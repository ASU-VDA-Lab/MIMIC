module fake_netlist_6_959_n_4544 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4544);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4544;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_2576;
wire n_1458;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_700;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3904;
wire n_3757;
wire n_4178;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_544;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_4417;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3655;
wire n_3452;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4255;
wire n_4071;
wire n_4403;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_451;
wire n_824;
wire n_686;
wire n_4297;
wire n_4102;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3910;
wire n_1699;
wire n_3812;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_433;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_4372;
wire n_982;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4161;
wire n_4130;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_612;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_2254;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_437;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_2178;
wire n_701;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_678;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_627;
wire n_595;
wire n_3253;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3337;
wire n_3450;
wire n_3431;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1627;
wire n_1295;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_673;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_872;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4540;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3426;
wire n_1788;
wire n_3158;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3353;
wire n_3018;
wire n_3150;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2650;
wire n_581;
wire n_2002;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2717;
wire n_1723;
wire n_2191;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3580;
wire n_705;
wire n_3418;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_446;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_4459;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1774;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_623;
wire n_3103;
wire n_3032;
wire n_3638;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3641;
wire n_767;
wire n_3591;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_4533;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_444;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_4362;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_4430;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_4428;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2502;
wire n_2131;
wire n_488;
wire n_2226;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3816;
wire n_3386;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2995;
wire n_2955;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_501;
wire n_956;
wire n_2276;
wire n_960;
wire n_3234;
wire n_4422;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_4126;
wire n_3870;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3250;
wire n_3276;
wire n_1934;
wire n_3194;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_4420;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3926;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1397;
wire n_1037;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4192;
wire n_4109;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4174;
wire n_1870;
wire n_2964;
wire n_4144;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_450;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_4258;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2699;
wire n_2272;
wire n_2200;
wire n_3029;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4135;
wire n_4209;
wire n_2871;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_2258;
wire n_1485;
wire n_1640;
wire n_4040;
wire n_804;
wire n_4461;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_431;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1794;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_706;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_4493;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2923;
wire n_2888;
wire n_2715;
wire n_2793;
wire n_1804;
wire n_2885;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2588;
wire n_2070;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_4203;
wire n_3515;
wire n_1150;
wire n_4505;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_875;
wire n_4462;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4543;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4173;
wire n_2752;
wire n_4157;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_691;
wire n_535;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_452;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_445;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2465;
wire n_1112;
wire n_2275;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1737;
wire n_1464;
wire n_653;
wire n_2430;
wire n_1414;
wire n_3584;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_576;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_839;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_3868;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_4115;
wire n_2999;
wire n_3796;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_570;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4353;
wire n_1789;
wire n_2531;
wire n_4104;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4351;
wire n_4346;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_436;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_756;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_635;
wire n_1194;
wire n_3374;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4538;
wire n_2640;
wire n_3695;
wire n_4254;
wire n_1051;
wire n_3976;
wire n_4051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4522;
wire n_4148;
wire n_2461;
wire n_2215;
wire n_571;
wire n_2001;
wire n_4341;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_679;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_665;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3896;
wire n_2774;
wire n_3815;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_827;
wire n_531;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_394),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_400),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_282),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_168),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_249),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_191),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_356),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_361),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_180),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_127),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_201),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_412),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_37),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_230),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_281),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_242),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_62),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_188),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_422),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_276),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_182),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_102),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_78),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_220),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_205),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_136),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_83),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_50),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_299),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_50),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_367),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_123),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_354),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_271),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_193),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_405),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_138),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_288),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_32),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_189),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_103),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_106),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_225),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_397),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_74),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_86),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_301),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_339),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_104),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_371),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_318),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_34),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_379),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_246),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_306),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_415),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_259),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_30),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_420),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_331),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_319),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_45),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_190),
.Y(n_497)
);

INVx4_ASAP7_75t_R g498 ( 
.A(n_107),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_364),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_258),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_188),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_386),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_43),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_290),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_201),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_298),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_184),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_269),
.Y(n_509)
);

BUFx8_ASAP7_75t_SL g510 ( 
.A(n_99),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_125),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_384),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_83),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_408),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_95),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_106),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_270),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_407),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_51),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_228),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_325),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_47),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_17),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_35),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_343),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_423),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_409),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_218),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_419),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_414),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_401),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_45),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_0),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_177),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_344),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_13),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_272),
.Y(n_537)
);

BUFx8_ASAP7_75t_SL g538 ( 
.A(n_279),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_64),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_121),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_26),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_126),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_383),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_145),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_322),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_257),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_86),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_224),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_6),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_425),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_350),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_342),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_78),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_359),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_351),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_163),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_358),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_402),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_129),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_341),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_57),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_42),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_413),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_382),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_94),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_378),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_118),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_233),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_173),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_295),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_428),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_126),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_391),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_247),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_363),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_374),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_232),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_138),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_284),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_330),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_192),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_155),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_151),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_196),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_4),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_114),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_190),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_166),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_74),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_147),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_161),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_122),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_268),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_392),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_309),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_264),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_8),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_113),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_135),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_357),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_173),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_196),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_326),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_110),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_240),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_197),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_7),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_137),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_102),
.Y(n_609)
);

BUFx2_ASAP7_75t_SL g610 ( 
.A(n_33),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_103),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_139),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_416),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_48),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_6),
.Y(n_615)
);

BUFx5_ASAP7_75t_L g616 ( 
.A(n_87),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_227),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_191),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_112),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_113),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_410),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_104),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_327),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_254),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_107),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_315),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_144),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_143),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_13),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_42),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_136),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_174),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_210),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_404),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_147),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_395),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_219),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_17),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_70),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_287),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_43),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_417),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_108),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_33),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_115),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_89),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_3),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_280),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_229),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_121),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_244),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_213),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_36),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_112),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_256),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_58),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_360),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_177),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_355),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_65),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_101),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_189),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_19),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_3),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_427),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_122),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_7),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_93),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_123),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_385),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_1),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_260),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_311),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_56),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_429),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_149),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_292),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_321),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_368),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_37),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_34),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_67),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_69),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_411),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_255),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_192),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_130),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_156),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_424),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_418),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_76),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_64),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_130),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_90),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_317),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_406),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_93),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_273),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_115),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_71),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_377),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_234),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_0),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_253),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_166),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_365),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_403),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_163),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_23),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_167),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_430),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_362),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_159),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_349),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_62),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_81),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_387),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_117),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_314),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_21),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_333),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_380),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_120),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_11),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_41),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_56),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_16),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_211),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_426),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_304),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_9),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_296),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_262),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_19),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_116),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_198),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_128),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_49),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_389),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_261),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_399),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_340),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_346),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_222),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_11),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_213),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_118),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_211),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_171),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_165),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_180),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_167),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_23),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_144),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_275),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_16),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_373),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_133),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_202),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_376),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_390),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_510),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_654),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_616),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_616),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_616),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_699),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_501),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_616),
.Y(n_769)
);

CKINVDCx16_ASAP7_75t_R g770 ( 
.A(n_560),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_616),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_536),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_616),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_515),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_616),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_448),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_503),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_616),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_720),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_720),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_508),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_671),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_720),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_511),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_720),
.Y(n_785)
);

BUFx5_ASAP7_75t_L g786 ( 
.A(n_435),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_720),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_720),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_720),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_681),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_443),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_720),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_565),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_565),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_516),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_513),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_519),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_565),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_513),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_533),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_520),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_533),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_581),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_581),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_629),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_522),
.Y(n_806)
);

CKINVDCx14_ASAP7_75t_R g807 ( 
.A(n_442),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_629),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_455),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_532),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_688),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_688),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_539),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_434),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_534),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_434),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_747),
.B(n_1),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_434),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_434),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_540),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_544),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_434),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_437),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_437),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_647),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_437),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_437),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_437),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_569),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_660),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_547),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_553),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_569),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_440),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_561),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_562),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_567),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_636),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_569),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_569),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_569),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_572),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_450),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_582),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_584),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_583),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_458),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_459),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_449),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_460),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_461),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_714),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_449),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_475),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_480),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_676),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_496),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_633),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_680),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_506),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_583),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_687),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_627),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_523),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_473),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_627),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_524),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_528),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_644),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_542),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_548),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_448),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_697),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_644),
.Y(n_874)
);

NOR2xp67_ASAP7_75t_L g875 ( 
.A(n_466),
.B(n_2),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_588),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_549),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_556),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_716),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_589),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_559),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_578),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_585),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_586),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_591),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_650),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_650),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_592),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_465),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_473),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_597),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_710),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_587),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_710),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_590),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_521),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_752),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_473),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_521),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_448),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_543),
.Y(n_901)
);

CKINVDCx16_ASAP7_75t_R g902 ( 
.A(n_711),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_607),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_614),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_618),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_619),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_620),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_440),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_622),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_630),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_637),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_598),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_441),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_441),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_723),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_445),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_645),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_599),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_646),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_612),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_652),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_653),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_667),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_445),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_669),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_683),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_723),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_601),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_726),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_602),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_604),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_726),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_606),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_608),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_686),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_691),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_612),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_692),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_609),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_452),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_700),
.Y(n_941)
);

INVxp33_ASAP7_75t_L g942 ( 
.A(n_703),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_724),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_611),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_725),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_452),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_728),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_734),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_617),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_448),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_745),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_543),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_625),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_545),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_448),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_628),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_545),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_447),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_451),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_690),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_631),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_488),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_612),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_632),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_690),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_456),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_635),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_638),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_656),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_639),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_489),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_526),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_535),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_537),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_546),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_641),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_643),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_649),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_656),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_478),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_551),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_554),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_658),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_456),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_690),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_656),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_555),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_478),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_661),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_564),
.Y(n_990)
);

BUFx8_ASAP7_75t_SL g991 ( 
.A(n_538),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_579),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_600),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_662),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_663),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_457),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_664),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_603),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_640),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_666),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_613),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_668),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_457),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_674),
.Y(n_1004)
);

INVxp33_ASAP7_75t_SL g1005 ( 
.A(n_462),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_621),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_642),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_659),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_655),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_684),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_682),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_696),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_702),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_518),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_719),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_729),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_610),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_466),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_690),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_739),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_690),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_693),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_694),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_755),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_760),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_462),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_761),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_468),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_468),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_760),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_464),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_505),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_464),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_505),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_469),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_527),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_527),
.Y(n_1037)
);

INVxp33_ASAP7_75t_L g1038 ( 
.A(n_557),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_469),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_471),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_557),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_717),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_471),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_474),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_717),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_478),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_465),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_474),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_472),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_760),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_472),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_476),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_568),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_568),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_476),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_541),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_594),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_477),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_594),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_757),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_757),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_760),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_615),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_760),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_477),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_479),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_615),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_705),
.B(n_2),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_759),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_479),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_705),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_708),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_708),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_431),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_483),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_431),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_483),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_432),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_432),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_433),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_481),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_433),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_436),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_486),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_436),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_481),
.Y(n_1086)
);

INVxp33_ASAP7_75t_L g1087 ( 
.A(n_486),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_438),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_438),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_577),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_439),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_492),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_481),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_759),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_439),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_444),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_444),
.Y(n_1097)
);

INVxp67_ASAP7_75t_SL g1098 ( 
.A(n_730),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_492),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_446),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_446),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_453),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_453),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_497),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_454),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_454),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_497),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_709),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_463),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_709),
.Y(n_1110)
);

INVxp67_ASAP7_75t_SL g1111 ( 
.A(n_634),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_463),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_713),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_704),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_713),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_715),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_715),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_718),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_718),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_467),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_467),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_563),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_732),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_727),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_727),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_1081),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_816),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_818),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_815),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_819),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_814),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_814),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_991),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_822),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_823),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_826),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_827),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1038),
.B(n_514),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_815),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_828),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_829),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_1081),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_833),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_825),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_762),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1056),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_825),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_856),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_840),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1074),
.B(n_502),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_763),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_793),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_762),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_856),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_794),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_798),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_824),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_824),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_1081),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_839),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_839),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_768),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_768),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_862),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_841),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_841),
.Y(n_1166)
);

INVxp67_ASAP7_75t_SL g1167 ( 
.A(n_1081),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_862),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_873),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_958),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_873),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_1014),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_959),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_777),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_1090),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_777),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_962),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_781),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_971),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_781),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_784),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_1123),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_972),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_973),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_784),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_908),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_974),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_1069),
.B(n_470),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_807),
.B(n_657),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1081),
.B(n_1120),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_908),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_795),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_795),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_975),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_797),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_981),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_982),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_987),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_990),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_992),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_797),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_1017),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_993),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_998),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_801),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_965),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_940),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1001),
.Y(n_1208)
);

INVxp33_ASAP7_75t_SL g1209 ( 
.A(n_763),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_940),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_946),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1006),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_767),
.Y(n_1213)
);

INVxp33_ASAP7_75t_L g1214 ( 
.A(n_913),
.Y(n_1214)
);

INVxp67_ASAP7_75t_SL g1215 ( 
.A(n_1076),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_801),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1007),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_946),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_806),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_806),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1008),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_996),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1010),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1012),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_965),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_L g1226 ( 
.A(n_1078),
.B(n_470),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1079),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1080),
.B(n_482),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1013),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_996),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1003),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1015),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1016),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_810),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1020),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1003),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1024),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1031),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1027),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1031),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_843),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_810),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_847),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_848),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1066),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1066),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_850),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_851),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_985),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1082),
.B(n_504),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_849),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_854),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_855),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1083),
.B(n_563),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_813),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_767),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1070),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1070),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_813),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_857),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_1085),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1075),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_820),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_860),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_820),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_L g1266 ( 
.A(n_1088),
.B(n_482),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_864),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_867),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_868),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1075),
.Y(n_1270)
);

INVxp33_ASAP7_75t_L g1271 ( 
.A(n_916),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_870),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_871),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1077),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1077),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1108),
.Y(n_1276)
);

INVxp67_ASAP7_75t_SL g1277 ( 
.A(n_1089),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_877),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_821),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_878),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1058),
.B(n_731),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_881),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_882),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_883),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_924),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_884),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1108),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_821),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_966),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_831),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_776),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_831),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1116),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_893),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1116),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_895),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_832),
.Y(n_1297)
);

NOR2xp67_ASAP7_75t_L g1298 ( 
.A(n_1091),
.B(n_484),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_985),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_832),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_969),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_791),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_835),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_903),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_904),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_905),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_835),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1019),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1019),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_906),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_836),
.Y(n_1311)
);

BUFx2_ASAP7_75t_SL g1312 ( 
.A(n_1111),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_809),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_836),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_907),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_830),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_837),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_909),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_859),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_910),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_879),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_911),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_837),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_917),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_897),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1021),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_919),
.Y(n_1327)
);

INVxp33_ASAP7_75t_L g1328 ( 
.A(n_1035),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_842),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_842),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1095),
.B(n_484),
.Y(n_1331)
);

INVxp33_ASAP7_75t_SL g1332 ( 
.A(n_844),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_849),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1096),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_921),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_922),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_923),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1097),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_844),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_770),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_845),
.Y(n_1341)
);

INVxp33_ASAP7_75t_SL g1342 ( 
.A(n_845),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_876),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_925),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_876),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_926),
.Y(n_1346)
);

INVxp67_ASAP7_75t_SL g1347 ( 
.A(n_1100),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_935),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_776),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_936),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_938),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_838),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_941),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_902),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_943),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_898),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_880),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_945),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_947),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_880),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1021),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_885),
.Y(n_1362)
);

XOR2xp5_ASAP7_75t_L g1363 ( 
.A(n_1114),
.B(n_740),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_885),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_888),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_948),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_888),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_891),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_891),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_912),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_912),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_918),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_918),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_928),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_951),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_1101),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_799),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_928),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1124),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_800),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_802),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_803),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1125),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1092),
.B(n_731),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_930),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_930),
.Y(n_1386)
);

CKINVDCx16_ASAP7_75t_R g1387 ( 
.A(n_980),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_980),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_931),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_931),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_933),
.Y(n_1391)
);

INVxp33_ASAP7_75t_SL g1392 ( 
.A(n_933),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_934),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_834),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_934),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_939),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1102),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_939),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1103),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_853),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1119),
.B(n_735),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_944),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_944),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_834),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1105),
.B(n_485),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_949),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_804),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_805),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_808),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_949),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_811),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_764),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_953),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_765),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_953),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1106),
.B(n_507),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1109),
.B(n_485),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_766),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1112),
.B(n_487),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1121),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_956),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_852),
.B(n_487),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_769),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_956),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_771),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_961),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_961),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_964),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_773),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_964),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_967),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1291),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1138),
.B(n_1068),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1251),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1377),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1126),
.B(n_899),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1380),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1146),
.A2(n_1005),
.B1(n_736),
.B2(n_737),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1215),
.A2(n_1009),
.B1(n_1098),
.B2(n_999),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1381),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1131),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1142),
.B(n_901),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1412),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1152),
.B(n_952),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1131),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1132),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1414),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1418),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1423),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1356),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1155),
.B(n_954),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1425),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1227),
.A2(n_1026),
.B1(n_1039),
.B2(n_1033),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1132),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1159),
.B(n_786),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1382),
.Y(n_1456)
);

INVx5_ASAP7_75t_L g1457 ( 
.A(n_1291),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1291),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1285),
.A2(n_968),
.B1(n_970),
.B2(n_967),
.Y(n_1459)
);

AOI22x1_ASAP7_75t_SL g1460 ( 
.A1(n_1186),
.A2(n_736),
.B1(n_737),
.B2(n_735),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1321),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1167),
.B(n_786),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1161),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1407),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1291),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1251),
.B(n_846),
.Y(n_1466)
);

INVx5_ASAP7_75t_L g1467 ( 
.A(n_1349),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1349),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1161),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1408),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1409),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1261),
.A2(n_1026),
.B1(n_1039),
.B2(n_1033),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1206),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1206),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1411),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1241),
.Y(n_1476)
);

AND2x6_ASAP7_75t_L g1477 ( 
.A(n_1190),
.B(n_775),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1225),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1225),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1429),
.A2(n_783),
.B(n_778),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1333),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1249),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1156),
.B(n_957),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1243),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1249),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1127),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1254),
.B(n_853),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1128),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1302),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1299),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1299),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1363),
.A2(n_1005),
.B1(n_744),
.B2(n_746),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1349),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1308),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1302),
.Y(n_1495)
);

AND2x2_ASAP7_75t_SL g1496 ( 
.A(n_1189),
.B(n_1068),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1130),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1349),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1134),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1313),
.A2(n_744),
.B1(n_746),
.B2(n_738),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1277),
.B(n_896),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1308),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1135),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1313),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1136),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1309),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1137),
.Y(n_1507)
);

AND2x6_ASAP7_75t_L g1508 ( 
.A(n_1331),
.B(n_787),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1140),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_R g1510 ( 
.A(n_1133),
.B(n_968),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1289),
.A2(n_976),
.B1(n_977),
.B2(n_970),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1309),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1326),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1333),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1326),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1334),
.B(n_896),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1361),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1361),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1141),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1400),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1400),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1143),
.Y(n_1522)
);

BUFx8_ASAP7_75t_L g1523 ( 
.A(n_1281),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1338),
.B(n_846),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1157),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1149),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1150),
.A2(n_780),
.B(n_779),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1158),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1316),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1209),
.B(n_920),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1160),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1244),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1347),
.B(n_861),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1316),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1165),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1247),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1376),
.B(n_1047),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1248),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1387),
.B(n_976),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1252),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1253),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1166),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1260),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1170),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1250),
.A2(n_1416),
.B(n_780),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1226),
.B(n_988),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1173),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1177),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1179),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1420),
.B(n_861),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1319),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1264),
.Y(n_1553)
);

AND2x2_ASAP7_75t_SL g1554 ( 
.A(n_1422),
.B(n_1086),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_R g1555 ( 
.A(n_1145),
.B(n_977),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1183),
.B(n_1049),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1267),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1184),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1405),
.B(n_978),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1187),
.B(n_1051),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1194),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1228),
.B(n_786),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1384),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1401),
.A2(n_1043),
.B1(n_1044),
.B2(n_1040),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1196),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1268),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1197),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1379),
.A2(n_983),
.B1(n_989),
.B2(n_978),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1269),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1198),
.A2(n_789),
.B(n_788),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1266),
.B(n_786),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1199),
.B(n_863),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1298),
.B(n_1417),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1200),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1203),
.B(n_863),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1419),
.B(n_786),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1204),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1272),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1208),
.B(n_1053),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1212),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1273),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1217),
.B(n_1054),
.Y(n_1582)
);

CKINVDCx16_ASAP7_75t_R g1583 ( 
.A(n_1319),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1202),
.B(n_786),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1278),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1221),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1223),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1332),
.B(n_983),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1224),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1229),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1232),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1233),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1235),
.B(n_1057),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1237),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1239),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1342),
.B(n_989),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1280),
.Y(n_1597)
);

INVx5_ASAP7_75t_L g1598 ( 
.A(n_1388),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1282),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_L g1600 ( 
.A(n_1188),
.B(n_988),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_SL g1601 ( 
.A1(n_1325),
.A2(n_748),
.B1(n_749),
.B2(n_738),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1283),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1284),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1286),
.B(n_866),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1325),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1294),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1296),
.A2(n_792),
.B(n_1025),
.Y(n_1607)
);

AOI22x1_ASAP7_75t_R g1608 ( 
.A1(n_1340),
.A2(n_1110),
.B1(n_1094),
.B2(n_1067),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1304),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1394),
.A2(n_1043),
.B1(n_1044),
.B2(n_1040),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1305),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1306),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1151),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1310),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1315),
.A2(n_785),
.B(n_779),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1318),
.B(n_1059),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1320),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1322),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1324),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1327),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1335),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1336),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1172),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1337),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1344),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1346),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1348),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1350),
.B(n_786),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1351),
.B(n_866),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1353),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1355),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1404),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1172),
.A2(n_749),
.B1(n_750),
.B2(n_748),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1358),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1359),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1366),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1375),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1383),
.B(n_1060),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1162),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1300),
.B(n_869),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1312),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1163),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1303),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1392),
.B(n_994),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1343),
.Y(n_1645)
);

INVx5_ASAP7_75t_L g1646 ( 
.A(n_1345),
.Y(n_1646)
);

AND2x6_ASAP7_75t_L g1647 ( 
.A(n_1174),
.B(n_1086),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1421),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1213),
.Y(n_1649)
);

AND2x6_ASAP7_75t_L g1650 ( 
.A(n_1176),
.B(n_1093),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1178),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1180),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1256),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1181),
.B(n_869),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1185),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1192),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1193),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1195),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1175),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1201),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_L g1661 ( 
.A(n_1340),
.B(n_1046),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1214),
.B(n_1061),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1205),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1216),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1219),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1220),
.B(n_874),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1234),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1271),
.B(n_874),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1242),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1255),
.B(n_786),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1328),
.A2(n_785),
.B(n_1025),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1259),
.B(n_994),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1263),
.B(n_886),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1265),
.A2(n_1064),
.B(n_1030),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1279),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1288),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1431),
.B(n_995),
.Y(n_1677)
);

BUFx8_ASAP7_75t_L g1678 ( 
.A(n_1352),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1290),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1292),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1297),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1307),
.B(n_995),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1311),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1314),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1317),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1323),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1329),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1330),
.B(n_886),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1339),
.A2(n_1000),
.B1(n_1002),
.B2(n_997),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1341),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1175),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1360),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1368),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1369),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1372),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1389),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1390),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1391),
.B(n_887),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1393),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1396),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1182),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1402),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1403),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1406),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1410),
.Y(n_1705)
);

BUFx3_ASAP7_75t_L g1706 ( 
.A(n_1413),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1415),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1426),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1427),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1428),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1153),
.B(n_997),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1357),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1357),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1362),
.B(n_1000),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1352),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1354),
.B(n_887),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1354),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1362),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1182),
.B(n_892),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1364),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1510),
.Y(n_1721)
);

NOR2xp67_ASAP7_75t_L g1722 ( 
.A(n_1450),
.B(n_1002),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1555),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1615),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_R g1725 ( 
.A(n_1489),
.B(n_1048),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1548),
.B(n_1004),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1641),
.B(n_1093),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1548),
.B(n_1436),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1461),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1668),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1623),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_1583),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1719),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1615),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1466),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1466),
.Y(n_1736)
);

AOI21x1_ASAP7_75t_L g1737 ( 
.A1(n_1562),
.A2(n_1064),
.B(n_1030),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1481),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1623),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1719),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1466),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1489),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_R g1743 ( 
.A(n_1659),
.B(n_1129),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1590),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1659),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_R g1746 ( 
.A(n_1605),
.B(n_1129),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1605),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1590),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_R g1749 ( 
.A(n_1663),
.B(n_1139),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1504),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1592),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1678),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1678),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1668),
.B(n_1087),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1678),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1598),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1654),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1481),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_R g1759 ( 
.A(n_1663),
.B(n_1139),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1651),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1651),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1592),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1607),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1607),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1706),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1706),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1504),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1639),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_1639),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1688),
.B(n_937),
.Y(n_1770)
);

CKINVDCx14_ASAP7_75t_R g1771 ( 
.A(n_1691),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1495),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1691),
.Y(n_1773)
);

BUFx10_ASAP7_75t_L g1774 ( 
.A(n_1711),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1639),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1607),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1639),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1595),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1639),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1642),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1642),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_R g1782 ( 
.A(n_1632),
.B(n_1048),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1719),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1595),
.Y(n_1784)
);

NOR2xp67_ASAP7_75t_L g1785 ( 
.A(n_1598),
.B(n_1652),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1642),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1716),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1642),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1599),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1642),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1599),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1656),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1433),
.A2(n_1011),
.B1(n_1022),
.B2(n_1004),
.Y(n_1793)
);

INVxp33_ASAP7_75t_SL g1794 ( 
.A(n_1530),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1603),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_R g1796 ( 
.A(n_1663),
.B(n_1144),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1559),
.B(n_1563),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1656),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1656),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1656),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1603),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1656),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1667),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1667),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1514),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1667),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1667),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1667),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1572),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1683),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1641),
.B(n_1011),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1701),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1683),
.Y(n_1813)
);

AND2x6_ASAP7_75t_L g1814 ( 
.A(n_1670),
.B(n_1122),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1570),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1683),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1572),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1683),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_R g1819 ( 
.A(n_1710),
.B(n_1144),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1572),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1575),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1575),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1575),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1442),
.B(n_1022),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1570),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_R g1826 ( 
.A(n_1710),
.B(n_1147),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1441),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1716),
.Y(n_1828)
);

CKINVDCx20_ASAP7_75t_R g1829 ( 
.A(n_1701),
.Y(n_1829)
);

CKINVDCx16_ASAP7_75t_R g1830 ( 
.A(n_1529),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_1534),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1604),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1683),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1685),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1688),
.B(n_986),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1573),
.B(n_1023),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1570),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1685),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_R g1839 ( 
.A(n_1632),
.B(n_1052),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1685),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1443),
.B(n_1023),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1716),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1685),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1574),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1552),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1685),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1687),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1687),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1443),
.B(n_1122),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1674),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1687),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1604),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1687),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1441),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1687),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1604),
.Y(n_1857)
);

CKINVDCx20_ASAP7_75t_R g1858 ( 
.A(n_1523),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1696),
.Y(n_1859)
);

CKINVDCx20_ASAP7_75t_R g1860 ( 
.A(n_1523),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1629),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_R g1862 ( 
.A(n_1710),
.B(n_1147),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1433),
.B(n_979),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1629),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1629),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_1523),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1544),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1598),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1598),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1696),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1715),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1445),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1696),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1574),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1696),
.Y(n_1875)
);

INVx3_ASAP7_75t_L g1876 ( 
.A(n_1674),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1445),
.Y(n_1877)
);

INVxp67_ASAP7_75t_R g1878 ( 
.A(n_1675),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_R g1879 ( 
.A(n_1598),
.B(n_1148),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1696),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1709),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1544),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1547),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1662),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1564),
.B(n_914),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1709),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1447),
.B(n_1052),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1446),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1446),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1654),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1709),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1547),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1709),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1610),
.B(n_914),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1448),
.B(n_1065),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1717),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1709),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1550),
.Y(n_1898)
);

CKINVDCx20_ASAP7_75t_R g1899 ( 
.A(n_1717),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1550),
.Y(n_1900)
);

AND3x2_ASAP7_75t_L g1901 ( 
.A(n_1679),
.B(n_774),
.C(n_984),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1652),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1652),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1700),
.Y(n_1904)
);

NOR2xp67_ASAP7_75t_L g1905 ( 
.A(n_1700),
.B(n_865),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1700),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1558),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1454),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1588),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1454),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1717),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1717),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1561),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1596),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1717),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1561),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1463),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1492),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1654),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1514),
.Y(n_1920)
);

NOR2xp67_ASAP7_75t_L g1921 ( 
.A(n_1689),
.B(n_890),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1565),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1463),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1520),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1520),
.Y(n_1925)
);

NOR2xp67_ASAP7_75t_L g1926 ( 
.A(n_1459),
.B(n_963),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1672),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1565),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1666),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1469),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1558),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1469),
.Y(n_1932)
);

NAND2xp33_ASAP7_75t_R g1933 ( 
.A(n_1714),
.B(n_1065),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1558),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1580),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1677),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1682),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1657),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1657),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1658),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1473),
.Y(n_1941)
);

BUFx3_ASAP7_75t_L g1942 ( 
.A(n_1434),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1658),
.Y(n_1943)
);

NOR2xp67_ASAP7_75t_L g1944 ( 
.A(n_1511),
.B(n_782),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1660),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1666),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1660),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_R g1948 ( 
.A(n_1655),
.B(n_1148),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1664),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1664),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1580),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1666),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1673),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1665),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1665),
.Y(n_1955)
);

CKINVDCx20_ASAP7_75t_R g1956 ( 
.A(n_1633),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1586),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1473),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1669),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1669),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1586),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1496),
.B(n_1084),
.Y(n_1962)
);

NAND2xp33_ASAP7_75t_R g1963 ( 
.A(n_1643),
.B(n_1084),
.Y(n_1963)
);

OAI22xp33_ASAP7_75t_R g1964 ( 
.A1(n_1718),
.A2(n_979),
.B1(n_772),
.B2(n_1094),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1474),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1539),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1681),
.Y(n_1967)
);

CKINVDCx20_ASAP7_75t_R g1968 ( 
.A(n_1500),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1681),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1684),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1673),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1449),
.B(n_1099),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_R g1973 ( 
.A(n_1655),
.B(n_1154),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1589),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1496),
.B(n_1099),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1434),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1589),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1453),
.B(n_1104),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1684),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1662),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1695),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_R g1982 ( 
.A(n_1676),
.B(n_1154),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1695),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1591),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1591),
.Y(n_1985)
);

BUFx3_ASAP7_75t_L g1986 ( 
.A(n_1521),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1474),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1699),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1699),
.Y(n_1989)
);

INVxp33_ASAP7_75t_SL g1990 ( 
.A(n_1438),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1478),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1702),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1702),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1704),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1704),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1478),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_R g1997 ( 
.A(n_1676),
.B(n_1164),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1479),
.Y(n_1998)
);

CKINVDCx20_ASAP7_75t_R g1999 ( 
.A(n_1601),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1521),
.Y(n_2000)
);

CKINVDCx20_ASAP7_75t_R g2001 ( 
.A(n_1460),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1460),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1707),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_R g2004 ( 
.A(n_1708),
.B(n_1164),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1707),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1594),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1673),
.Y(n_2007)
);

AND2x6_ASAP7_75t_L g2008 ( 
.A(n_1600),
.B(n_1110),
.Y(n_2008)
);

CKINVDCx20_ASAP7_75t_R g2009 ( 
.A(n_1568),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1674),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_R g2011 ( 
.A(n_1643),
.B(n_1104),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1608),
.Y(n_2012)
);

INVxp67_ASAP7_75t_SL g2013 ( 
.A(n_1506),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1594),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1647),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1770),
.B(n_1718),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1721),
.Y(n_2017)
);

AND2x6_ASAP7_75t_L g2018 ( 
.A(n_1763),
.B(n_1501),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1735),
.Y(n_2019)
);

BUFx10_ASAP7_75t_L g2020 ( 
.A(n_1978),
.Y(n_2020)
);

NOR2x1p5_ASAP7_75t_L g2021 ( 
.A(n_1768),
.B(n_1708),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1763),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_1896),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1728),
.B(n_1501),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1835),
.B(n_1516),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1738),
.B(n_1640),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1736),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1730),
.B(n_1516),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1741),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1730),
.B(n_1554),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1757),
.B(n_1646),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1764),
.Y(n_2032)
);

INVx6_ASAP7_75t_L g2033 ( 
.A(n_1844),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1907),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1797),
.B(n_1645),
.Y(n_2035)
);

OAI22xp33_ASAP7_75t_SL g2036 ( 
.A1(n_1962),
.A2(n_1648),
.B1(n_1645),
.B2(n_1649),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1907),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1764),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1809),
.Y(n_2039)
);

INVx5_ASAP7_75t_L g2040 ( 
.A(n_1907),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1817),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1844),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1757),
.B(n_1646),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1726),
.B(n_1894),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1723),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1836),
.B(n_1554),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1885),
.B(n_1845),
.Y(n_2047)
);

INVx4_ASAP7_75t_SL g2048 ( 
.A(n_1814),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1827),
.Y(n_2049)
);

INVx4_ASAP7_75t_SL g2050 ( 
.A(n_1814),
.Y(n_2050)
);

INVx5_ASAP7_75t_L g2051 ( 
.A(n_1907),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1820),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1884),
.B(n_1980),
.Y(n_2053)
);

INVxp33_ASAP7_75t_L g2054 ( 
.A(n_1746),
.Y(n_2054)
);

INVx4_ASAP7_75t_L g2055 ( 
.A(n_1844),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1821),
.Y(n_2056)
);

INVx1_ASAP7_75t_SL g2057 ( 
.A(n_1729),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1738),
.B(n_1640),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1822),
.Y(n_2059)
);

INVx1_ASAP7_75t_SL g2060 ( 
.A(n_1754),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1827),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1855),
.Y(n_2062)
);

INVx4_ASAP7_75t_L g2063 ( 
.A(n_1844),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1855),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1823),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1975),
.B(n_1863),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1874),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1890),
.B(n_1698),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1872),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1872),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1832),
.Y(n_2071)
);

AND2x2_ASAP7_75t_SL g2072 ( 
.A(n_1874),
.B(n_1576),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1733),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_L g2074 ( 
.A1(n_1815),
.A2(n_1837),
.B1(n_1825),
.B2(n_1814),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1852),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1744),
.B(n_1748),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1857),
.Y(n_2077)
);

BUFx3_ASAP7_75t_L g2078 ( 
.A(n_1896),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_1927),
.B(n_1648),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1877),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1877),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1971),
.B(n_1646),
.Y(n_2082)
);

BUFx3_ASAP7_75t_L g2083 ( 
.A(n_1899),
.Y(n_2083)
);

BUFx3_ASAP7_75t_L g2084 ( 
.A(n_1899),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1861),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1874),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1888),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1936),
.B(n_1472),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_1815),
.A2(n_1508),
.B1(n_1477),
.B2(n_1480),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_1937),
.B(n_1680),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1864),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1751),
.B(n_1524),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1909),
.B(n_1686),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1931),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1914),
.B(n_1690),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1794),
.B(n_1692),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1888),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1889),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1794),
.B(n_1693),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1772),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1889),
.Y(n_2101)
);

OR2x6_ASAP7_75t_L g2102 ( 
.A(n_1971),
.B(n_1720),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1824),
.B(n_1694),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1769),
.B(n_1646),
.Y(n_2104)
);

NAND2xp33_ASAP7_75t_L g2105 ( 
.A(n_2015),
.B(n_1647),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1758),
.B(n_1640),
.Y(n_2106)
);

INVx2_ASAP7_75t_SL g2107 ( 
.A(n_1915),
.Y(n_2107)
);

INVx1_ASAP7_75t_SL g2108 ( 
.A(n_1750),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1865),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1867),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1919),
.B(n_1697),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1908),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1882),
.Y(n_2113)
);

INVx2_ASAP7_75t_SL g2114 ( 
.A(n_1938),
.Y(n_2114)
);

INVx4_ASAP7_75t_SL g2115 ( 
.A(n_1814),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1883),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1775),
.B(n_1646),
.Y(n_2117)
);

NAND2xp33_ASAP7_75t_L g2118 ( 
.A(n_2015),
.B(n_1647),
.Y(n_2118)
);

INVx4_ASAP7_75t_L g2119 ( 
.A(n_1874),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1892),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1908),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1777),
.B(n_1584),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1898),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1762),
.B(n_1524),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1900),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_1830),
.B(n_1720),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1778),
.B(n_1524),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1879),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_1911),
.Y(n_2129)
);

INVx8_ASAP7_75t_L g2130 ( 
.A(n_1911),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1929),
.B(n_1698),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1784),
.B(n_1533),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_1750),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_1740),
.B(n_1649),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1910),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1779),
.B(n_1558),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1913),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1910),
.Y(n_2138)
);

NAND2xp33_ASAP7_75t_L g2139 ( 
.A(n_1780),
.B(n_1647),
.Y(n_2139)
);

INVx4_ASAP7_75t_SL g2140 ( 
.A(n_1814),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1917),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1789),
.B(n_1533),
.Y(n_2142)
);

NAND2xp33_ASAP7_75t_SL g2143 ( 
.A(n_1781),
.B(n_1703),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1946),
.B(n_1698),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1931),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1917),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1743),
.Y(n_2147)
);

BUFx3_ASAP7_75t_L g2148 ( 
.A(n_1912),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1923),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_1952),
.B(n_1705),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1916),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1931),
.Y(n_2152)
);

INVx6_ASAP7_75t_L g2153 ( 
.A(n_1942),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1922),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1791),
.B(n_1533),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1928),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1923),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1930),
.Y(n_2158)
);

BUFx10_ASAP7_75t_L g2159 ( 
.A(n_1901),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1930),
.Y(n_2160)
);

NAND3xp33_ASAP7_75t_L g2161 ( 
.A(n_1793),
.B(n_1613),
.C(n_1439),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_1912),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_1953),
.B(n_1653),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1786),
.B(n_1558),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1795),
.B(n_1551),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_1727),
.A2(n_1508),
.B1(n_1814),
.B2(n_2007),
.Y(n_2166)
);

INVx1_ASAP7_75t_SL g2167 ( 
.A(n_1767),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1801),
.B(n_1551),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1854),
.B(n_1551),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1942),
.B(n_1508),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1932),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_1931),
.Y(n_2172)
);

BUFx10_ASAP7_75t_L g2173 ( 
.A(n_1747),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_1727),
.A2(n_1508),
.B1(n_1650),
.B2(n_1647),
.Y(n_2174)
);

AND3x1_ASAP7_75t_L g2175 ( 
.A(n_1887),
.B(n_1713),
.C(n_1712),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1932),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1976),
.B(n_1508),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_1939),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1749),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1934),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_1815),
.A2(n_1508),
.B1(n_1477),
.B2(n_1480),
.Y(n_2181)
);

INVx6_ASAP7_75t_L g2182 ( 
.A(n_1976),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1825),
.A2(n_1477),
.B1(n_1480),
.B2(n_774),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_1940),
.B(n_1653),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1935),
.B(n_1449),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_1758),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1951),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1722),
.B(n_1487),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1759),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_1825),
.A2(n_1477),
.B1(n_875),
.B2(n_1647),
.Y(n_2190)
);

INVx5_ASAP7_75t_L g2191 ( 
.A(n_1934),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1957),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1961),
.B(n_1452),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1974),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1788),
.B(n_1577),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_1790),
.B(n_1487),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1783),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_1895),
.B(n_1644),
.C(n_1113),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1941),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1792),
.B(n_1638),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1798),
.B(n_1799),
.Y(n_2201)
);

NAND2xp33_ASAP7_75t_SL g2202 ( 
.A(n_1800),
.B(n_1364),
.Y(n_2202)
);

INVx5_ASAP7_75t_L g2203 ( 
.A(n_1934),
.Y(n_2203)
);

INVx2_ASAP7_75t_SL g2204 ( 
.A(n_1943),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1802),
.B(n_1638),
.Y(n_2205)
);

BUFx10_ASAP7_75t_L g2206 ( 
.A(n_1731),
.Y(n_2206)
);

INVx4_ASAP7_75t_L g2207 ( 
.A(n_1803),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1804),
.B(n_1577),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1806),
.B(n_1577),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_1787),
.B(n_1712),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1941),
.Y(n_2211)
);

CKINVDCx5p33_ASAP7_75t_R g2212 ( 
.A(n_1796),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_1807),
.B(n_1537),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1958),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_1837),
.A2(n_1477),
.B1(n_1650),
.B2(n_1671),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_1934),
.Y(n_2216)
);

BUFx2_ASAP7_75t_L g2217 ( 
.A(n_1767),
.Y(n_2217)
);

INVx3_ASAP7_75t_L g2218 ( 
.A(n_1958),
.Y(n_2218)
);

INVx11_ASAP7_75t_L g2219 ( 
.A(n_2008),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1977),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1984),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1965),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1985),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_1808),
.B(n_1577),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2006),
.Y(n_2225)
);

BUFx10_ASAP7_75t_L g2226 ( 
.A(n_1739),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1810),
.B(n_1577),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1965),
.Y(n_2228)
);

AND2x6_ASAP7_75t_L g2229 ( 
.A(n_1850),
.B(n_1537),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1987),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1805),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2014),
.B(n_1452),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_SL g2233 ( 
.A(n_1813),
.B(n_1606),
.Y(n_2233)
);

INVx2_ASAP7_75t_SL g2234 ( 
.A(n_1945),
.Y(n_2234)
);

NAND2xp33_ASAP7_75t_L g2235 ( 
.A(n_1816),
.B(n_1650),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1849),
.B(n_1549),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1987),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1991),
.Y(n_2238)
);

AND2x6_ASAP7_75t_L g2239 ( 
.A(n_1850),
.B(n_1546),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_1837),
.A2(n_1477),
.B1(n_1650),
.B2(n_1671),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_1828),
.B(n_984),
.Y(n_2241)
);

NAND2xp33_ASAP7_75t_L g2242 ( 
.A(n_1818),
.B(n_1650),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1991),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_1947),
.B(n_1587),
.Y(n_2244)
);

AO22x2_ASAP7_75t_L g2245 ( 
.A1(n_1850),
.A2(n_790),
.B1(n_858),
.B2(n_1018),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_1949),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1996),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_1833),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1996),
.Y(n_2249)
);

INVx2_ASAP7_75t_SL g2250 ( 
.A(n_1950),
.Y(n_2250)
);

BUFx3_ASAP7_75t_L g2251 ( 
.A(n_1805),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1998),
.Y(n_2252)
);

INVx4_ASAP7_75t_SL g2253 ( 
.A(n_2008),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_1876),
.A2(n_1650),
.B1(n_1549),
.B2(n_1609),
.Y(n_2254)
);

INVx4_ASAP7_75t_L g2255 ( 
.A(n_1834),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1954),
.B(n_1587),
.Y(n_2256)
);

BUFx3_ASAP7_75t_L g2257 ( 
.A(n_1838),
.Y(n_2257)
);

CKINVDCx16_ASAP7_75t_R g2258 ( 
.A(n_1819),
.Y(n_2258)
);

AND3x1_ASAP7_75t_L g2259 ( 
.A(n_1972),
.B(n_1661),
.C(n_1560),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_1840),
.B(n_1606),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1998),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1724),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1724),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_1734),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1734),
.Y(n_2265)
);

INVx3_ASAP7_75t_L g2266 ( 
.A(n_1776),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1776),
.Y(n_2267)
);

INVx1_ASAP7_75t_SL g2268 ( 
.A(n_1831),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1955),
.B(n_1587),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_1959),
.B(n_1626),
.Y(n_2270)
);

AND2x2_ASAP7_75t_SL g2271 ( 
.A(n_1876),
.B(n_1626),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1776),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1986),
.Y(n_2273)
);

INVx5_ASAP7_75t_L g2274 ( 
.A(n_1876),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_2010),
.A2(n_1549),
.B1(n_1609),
.B2(n_1567),
.Y(n_2275)
);

INVx2_ASAP7_75t_SL g2276 ( 
.A(n_1960),
.Y(n_2276)
);

INVx5_ASAP7_75t_L g2277 ( 
.A(n_2010),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2010),
.A2(n_1990),
.B1(n_1727),
.B2(n_1964),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1842),
.Y(n_2279)
);

NAND2x1p5_ASAP7_75t_L g2280 ( 
.A(n_1986),
.B(n_2000),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1727),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1737),
.Y(n_2282)
);

OR2x2_ASAP7_75t_L g2283 ( 
.A(n_1841),
.B(n_1055),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1843),
.B(n_1055),
.Y(n_2284)
);

NAND2xp33_ASAP7_75t_L g2285 ( 
.A(n_1846),
.B(n_1606),
.Y(n_2285)
);

INVx4_ASAP7_75t_SL g2286 ( 
.A(n_2008),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1727),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1727),
.B(n_1567),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_1785),
.B(n_1476),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_1967),
.Y(n_2290)
);

NAND2xp33_ASAP7_75t_L g2291 ( 
.A(n_1847),
.B(n_1848),
.Y(n_2291)
);

OR2x6_ASAP7_75t_L g2292 ( 
.A(n_1905),
.B(n_1556),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2008),
.B(n_1567),
.Y(n_2293)
);

INVx4_ASAP7_75t_L g2294 ( 
.A(n_1851),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2008),
.B(n_1609),
.Y(n_2295)
);

BUFx6f_ASAP7_75t_L g2296 ( 
.A(n_2000),
.Y(n_2296)
);

AND2x4_ASAP7_75t_L g2297 ( 
.A(n_1853),
.B(n_1484),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2013),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_1969),
.B(n_1626),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1970),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_1856),
.Y(n_2301)
);

INVx2_ASAP7_75t_SL g2302 ( 
.A(n_1979),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_L g2303 ( 
.A1(n_1990),
.A2(n_1612),
.B1(n_1622),
.B2(n_817),
.Y(n_2303)
);

BUFx3_ASAP7_75t_L g2304 ( 
.A(n_1859),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1981),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1983),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2008),
.B(n_1612),
.Y(n_2307)
);

HB1xp67_ASAP7_75t_L g2308 ( 
.A(n_1870),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_1745),
.B(n_1811),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1756),
.B(n_1612),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_1933),
.A2(n_1622),
.B1(n_1619),
.B2(n_1606),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2024),
.B(n_1873),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2035),
.B(n_1875),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2035),
.B(n_1880),
.Y(n_2314)
);

OR2x6_ASAP7_75t_L g2315 ( 
.A(n_2130),
.B(n_1926),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_2025),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2103),
.B(n_1881),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2218),
.Y(n_2318)
);

NAND2xp33_ASAP7_75t_L g2319 ( 
.A(n_2229),
.B(n_1886),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2103),
.B(n_1891),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2213),
.B(n_2200),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2218),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2216),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2090),
.B(n_1893),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2039),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2046),
.B(n_1897),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2271),
.B(n_1988),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_2216),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2028),
.B(n_1989),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2090),
.B(n_1992),
.Y(n_2330)
);

NAND2xp33_ASAP7_75t_L g2331 ( 
.A(n_2229),
.B(n_1756),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_2205),
.B(n_1993),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2169),
.B(n_1994),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2030),
.B(n_1995),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2228),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2244),
.B(n_2005),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2044),
.B(n_2060),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2053),
.B(n_2003),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2016),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_2283),
.B(n_1774),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2053),
.B(n_1622),
.Y(n_2341)
);

INVxp33_ASAP7_75t_L g2342 ( 
.A(n_2184),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2041),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_2244),
.B(n_1902),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2188),
.B(n_1903),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2284),
.B(n_1878),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2052),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2228),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2066),
.B(n_1774),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2068),
.B(n_1904),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2271),
.B(n_1868),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2256),
.B(n_1906),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2049),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_2017),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_2256),
.B(n_2299),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2269),
.B(n_2299),
.Y(n_2356)
);

BUFx3_ASAP7_75t_L g2357 ( 
.A(n_2023),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2269),
.B(n_1774),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_L g2359 ( 
.A(n_2229),
.B(n_1868),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2270),
.B(n_1869),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2270),
.B(n_1869),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2076),
.B(n_1920),
.Y(n_2362)
);

INVx4_ASAP7_75t_L g2363 ( 
.A(n_2042),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2092),
.B(n_1924),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2056),
.Y(n_2365)
);

NAND3xp33_ASAP7_75t_L g2366 ( 
.A(n_2079),
.B(n_2184),
.C(n_2161),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2049),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_2096),
.B(n_1760),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2059),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2079),
.B(n_1761),
.Y(n_2370)
);

OAI221xp5_ASAP7_75t_L g2371 ( 
.A1(n_2088),
.A2(n_1944),
.B1(n_1921),
.B2(n_2011),
.C(n_1963),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_2096),
.B(n_1765),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_2216),
.Y(n_2373)
);

INVx2_ASAP7_75t_SL g2374 ( 
.A(n_2100),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2196),
.B(n_1766),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2124),
.B(n_1925),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2127),
.B(n_1606),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2132),
.B(n_1619),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2131),
.B(n_1826),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2099),
.B(n_1862),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2061),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2142),
.B(n_1619),
.Y(n_2382)
);

NOR2x1p5_ASAP7_75t_L g2383 ( 
.A(n_2257),
.B(n_1752),
.Y(n_2383)
);

INVx2_ASAP7_75t_SL g2384 ( 
.A(n_2023),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2061),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2155),
.B(n_2165),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2099),
.B(n_1966),
.Y(n_2387)
);

NAND2xp33_ASAP7_75t_L g2388 ( 
.A(n_2229),
.B(n_1948),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2078),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2168),
.B(n_1619),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2144),
.B(n_2065),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2114),
.B(n_1973),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2071),
.B(n_1619),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_2216),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2178),
.B(n_1982),
.Y(n_2395)
);

NAND3xp33_ASAP7_75t_L g2396 ( 
.A(n_2088),
.B(n_1839),
.C(n_1782),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2273),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2093),
.B(n_1966),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2093),
.B(n_2009),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2075),
.B(n_1624),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2077),
.B(n_1624),
.Y(n_2401)
);

BUFx3_ASAP7_75t_L g2402 ( 
.A(n_2078),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2085),
.B(n_2091),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2062),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2109),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2303),
.B(n_1624),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2019),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2303),
.B(n_1624),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2027),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2029),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2083),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_2095),
.B(n_2009),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2204),
.B(n_1771),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2237),
.Y(n_2414)
);

AOI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2229),
.A2(n_1968),
.B1(n_1999),
.B2(n_1918),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2234),
.B(n_1997),
.Y(n_2416)
);

INVx8_ASAP7_75t_L g2417 ( 
.A(n_2130),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2246),
.B(n_2004),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2062),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2163),
.B(n_1624),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2163),
.B(n_1625),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2249),
.Y(n_2422)
);

AND2x2_ASAP7_75t_SL g2423 ( 
.A(n_2291),
.B(n_1597),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2261),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2111),
.B(n_1625),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2111),
.B(n_1625),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_2072),
.B(n_1625),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2150),
.B(n_1625),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_2083),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_SL g2430 ( 
.A(n_2250),
.B(n_1521),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2150),
.B(n_1532),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2018),
.B(n_1536),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2095),
.B(n_1365),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2069),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2018),
.B(n_2185),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2276),
.B(n_1521),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2018),
.B(n_1538),
.Y(n_2437)
);

NAND3xp33_ASAP7_75t_L g2438 ( 
.A(n_2300),
.B(n_2306),
.C(n_2305),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2018),
.B(n_2193),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2290),
.B(n_1556),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_2302),
.B(n_1521),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2018),
.B(n_1540),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2232),
.B(n_1541),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2084),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2069),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2072),
.B(n_1571),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2297),
.B(n_1543),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2110),
.B(n_1553),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2080),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2036),
.B(n_1526),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2113),
.B(n_1557),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2080),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2081),
.Y(n_2453)
);

AOI22xp33_ASAP7_75t_L g2454 ( 
.A1(n_2183),
.A2(n_1968),
.B1(n_1999),
.B2(n_1918),
.Y(n_2454)
);

INVxp67_ASAP7_75t_L g2455 ( 
.A(n_2073),
.Y(n_2455)
);

AOI22xp5_ASAP7_75t_L g2456 ( 
.A1(n_2259),
.A2(n_1367),
.B1(n_1370),
.B2(n_1365),
.Y(n_2456)
);

NAND2xp33_ASAP7_75t_L g2457 ( 
.A(n_2042),
.B(n_1752),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2308),
.B(n_1560),
.Y(n_2458)
);

INVx4_ASAP7_75t_L g2459 ( 
.A(n_2042),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_R g2460 ( 
.A(n_2045),
.B(n_1725),
.Y(n_2460)
);

INVxp67_ASAP7_75t_L g2461 ( 
.A(n_2073),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2297),
.B(n_1566),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2257),
.B(n_1526),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2081),
.Y(n_2464)
);

NAND3xp33_ASAP7_75t_SL g2465 ( 
.A(n_2057),
.B(n_1370),
.C(n_1367),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_2301),
.B(n_1526),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2116),
.B(n_1569),
.Y(n_2467)
);

NOR2x1p5_ASAP7_75t_L g2468 ( 
.A(n_2301),
.B(n_1753),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2087),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2087),
.Y(n_2470)
);

NOR2xp67_ASAP7_75t_SL g2471 ( 
.A(n_2304),
.B(n_1753),
.Y(n_2471)
);

NOR2xp67_ASAP7_75t_L g2472 ( 
.A(n_2207),
.B(n_1755),
.Y(n_2472)
);

OAI221xp5_ASAP7_75t_L g2473 ( 
.A1(n_2241),
.A2(n_1585),
.B1(n_1611),
.B2(n_1581),
.C(n_1578),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2097),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2304),
.B(n_1526),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2120),
.B(n_1614),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2097),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2123),
.B(n_1618),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2047),
.B(n_1371),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2125),
.B(n_1627),
.Y(n_2480)
);

INVx2_ASAP7_75t_SL g2481 ( 
.A(n_2084),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2040),
.B(n_2051),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_2026),
.B(n_1631),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2201),
.B(n_1371),
.Y(n_2484)
);

INVx8_ASAP7_75t_L g2485 ( 
.A(n_2130),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2026),
.B(n_1634),
.Y(n_2486)
);

AO221x1_ASAP7_75t_L g2487 ( 
.A1(n_2245),
.A2(n_796),
.B1(n_812),
.B2(n_2012),
.C(n_1636),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2137),
.B(n_1635),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2098),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2098),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2101),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2201),
.B(n_1373),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2101),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2112),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2151),
.B(n_1637),
.Y(n_2495)
);

OAI221xp5_ASAP7_75t_L g2496 ( 
.A1(n_2134),
.A2(n_1440),
.B1(n_1456),
.B2(n_1437),
.C(n_1435),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2154),
.B(n_1486),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2054),
.B(n_1373),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2112),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2156),
.B(n_1486),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_2054),
.B(n_2020),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2187),
.B(n_1488),
.Y(n_2502)
);

NOR3xp33_ASAP7_75t_L g2503 ( 
.A(n_2198),
.B(n_1113),
.C(n_1107),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2121),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2040),
.B(n_1526),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2121),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2020),
.B(n_1374),
.Y(n_2507)
);

NOR2xp33_ASAP7_75t_L g2508 ( 
.A(n_2308),
.B(n_1374),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2192),
.B(n_1488),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_2197),
.B(n_1378),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2058),
.B(n_1464),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_L g2512 ( 
.A(n_2278),
.B(n_1115),
.C(n_1107),
.Y(n_2512)
);

INVx1_ASAP7_75t_SL g2513 ( 
.A(n_2126),
.Y(n_2513)
);

OR2x6_ASAP7_75t_L g2514 ( 
.A(n_2129),
.B(n_1597),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2040),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2194),
.B(n_1497),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2058),
.B(n_2106),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_L g2518 ( 
.A(n_2042),
.B(n_1755),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2220),
.B(n_1497),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2135),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2135),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2138),
.Y(n_2522)
);

INVx2_ASAP7_75t_SL g2523 ( 
.A(n_2129),
.Y(n_2523)
);

AND2x4_ASAP7_75t_L g2524 ( 
.A(n_2106),
.B(n_1602),
.Y(n_2524)
);

INVx2_ASAP7_75t_SL g2525 ( 
.A(n_2148),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2197),
.B(n_1579),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2221),
.B(n_2223),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2138),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2141),
.Y(n_2529)
);

AOI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2143),
.A2(n_1385),
.B1(n_1386),
.B2(n_1378),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2141),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2146),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2186),
.B(n_2231),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2225),
.B(n_1499),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2146),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2210),
.B(n_1385),
.Y(n_2536)
);

AOI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2292),
.A2(n_1395),
.B1(n_1398),
.B2(n_1386),
.Y(n_2537)
);

INVx1_ASAP7_75t_SL g2538 ( 
.A(n_2108),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2153),
.B(n_1499),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2149),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2107),
.B(n_1579),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2149),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2157),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2040),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_SL g2545 ( 
.A(n_2173),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2207),
.B(n_1395),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_2248),
.B(n_1470),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_L g2548 ( 
.A(n_2067),
.B(n_1471),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2157),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2133),
.Y(n_2550)
);

OAI22xp33_ASAP7_75t_L g2551 ( 
.A1(n_2292),
.A2(n_1956),
.B1(n_1617),
.B2(n_1620),
.Y(n_2551)
);

NAND3xp33_ASAP7_75t_L g2552 ( 
.A(n_2278),
.B(n_1117),
.C(n_1115),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2248),
.B(n_1475),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2255),
.B(n_1602),
.Y(n_2554)
);

INVx2_ASAP7_75t_SL g2555 ( 
.A(n_2148),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_2354),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2325),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2343),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2347),
.Y(n_2559)
);

NOR2xp67_ASAP7_75t_L g2560 ( 
.A(n_2366),
.B(n_2255),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2365),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2369),
.Y(n_2562)
);

INVxp67_ASAP7_75t_L g2563 ( 
.A(n_2513),
.Y(n_2563)
);

BUFx3_ASAP7_75t_L g2564 ( 
.A(n_2357),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2405),
.Y(n_2565)
);

BUFx4f_ASAP7_75t_L g2566 ( 
.A(n_2417),
.Y(n_2566)
);

HB1xp67_ASAP7_75t_L g2567 ( 
.A(n_2455),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2407),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2402),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2409),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2353),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_2533),
.B(n_2186),
.Y(n_2572)
);

AO22x2_ASAP7_75t_L g2573 ( 
.A1(n_2396),
.A2(n_2512),
.B1(n_2552),
.B2(n_2327),
.Y(n_2573)
);

INVxp67_ASAP7_75t_L g2574 ( 
.A(n_2337),
.Y(n_2574)
);

INVxp67_ASAP7_75t_L g2575 ( 
.A(n_2337),
.Y(n_2575)
);

OAI221xp5_ASAP7_75t_L g2576 ( 
.A1(n_2371),
.A2(n_2175),
.B1(n_2309),
.B2(n_2202),
.C(n_2268),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2374),
.Y(n_2577)
);

INVx4_ASAP7_75t_L g2578 ( 
.A(n_2417),
.Y(n_2578)
);

NAND2x1p5_ASAP7_75t_L g2579 ( 
.A(n_2533),
.B(n_2055),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2410),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2403),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2317),
.B(n_2294),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2527),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2321),
.B(n_2162),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2429),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2414),
.Y(n_2586)
);

AO22x2_ASAP7_75t_L g2587 ( 
.A1(n_2327),
.A2(n_2117),
.B1(n_2104),
.B2(n_2253),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2342),
.B(n_2320),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2422),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2424),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2367),
.Y(n_2591)
);

CKINVDCx20_ASAP7_75t_R g2592 ( 
.A(n_2460),
.Y(n_2592)
);

INVxp67_ASAP7_75t_L g2593 ( 
.A(n_2510),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2381),
.Y(n_2594)
);

AOI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2399),
.A2(n_1424),
.B1(n_1430),
.B2(n_1398),
.Y(n_2595)
);

AOI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2399),
.A2(n_1430),
.B1(n_1424),
.B2(n_1831),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2412),
.A2(n_1871),
.B1(n_1812),
.B2(n_1829),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2385),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2404),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2419),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2445),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2449),
.Y(n_2602)
);

AO22x2_ASAP7_75t_L g2603 ( 
.A1(n_2355),
.A2(n_2117),
.B1(n_2104),
.B2(n_2253),
.Y(n_2603)
);

NAND2x1p5_ASAP7_75t_L g2604 ( 
.A(n_2515),
.B(n_2055),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2452),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2453),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2313),
.B(n_2294),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2474),
.Y(n_2608)
);

AO22x2_ASAP7_75t_L g2609 ( 
.A1(n_2355),
.A2(n_2286),
.B1(n_2253),
.B2(n_2164),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2489),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2491),
.Y(n_2611)
);

AOI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2412),
.A2(n_1871),
.B1(n_1812),
.B2(n_1829),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2494),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2506),
.Y(n_2614)
);

AO22x2_ASAP7_75t_L g2615 ( 
.A1(n_2356),
.A2(n_2286),
.B1(n_2164),
.B2(n_2195),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2444),
.Y(n_2616)
);

AND2x4_ASAP7_75t_L g2617 ( 
.A(n_2517),
.B(n_2231),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2521),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2524),
.B(n_2251),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2528),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2529),
.Y(n_2621)
);

OAI221xp5_ASAP7_75t_L g2622 ( 
.A1(n_2433),
.A2(n_2167),
.B1(n_2279),
.B2(n_2102),
.C(n_1118),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2535),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_L g2624 ( 
.A(n_2314),
.B(n_1186),
.Y(n_2624)
);

AO22x2_ASAP7_75t_L g2625 ( 
.A1(n_2356),
.A2(n_2286),
.B1(n_2195),
.B2(n_2208),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2540),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2549),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2433),
.A2(n_1773),
.B1(n_1207),
.B2(n_1210),
.Y(n_2628)
);

AO22x2_ASAP7_75t_L g2629 ( 
.A1(n_2351),
.A2(n_2208),
.B1(n_2209),
.B2(n_2136),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2333),
.B(n_2326),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2434),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2464),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2375),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2312),
.B(n_2153),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2469),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2524),
.B(n_2251),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2526),
.B(n_2102),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2470),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2384),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2477),
.Y(n_2640)
);

AOI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2398),
.A2(n_1773),
.B1(n_1207),
.B2(n_1210),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2490),
.Y(n_2642)
);

NAND2x1p5_ASAP7_75t_L g2643 ( 
.A(n_2515),
.B(n_2063),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2514),
.B(n_2021),
.Y(n_2644)
);

NAND2x1_ASAP7_75t_L g2645 ( 
.A(n_2515),
.B(n_2264),
.Y(n_2645)
);

INVxp67_ASAP7_75t_L g2646 ( 
.A(n_2510),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2493),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2499),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2338),
.B(n_2153),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2458),
.B(n_2102),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2504),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2520),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2334),
.B(n_2182),
.Y(n_2653)
);

NOR2xp67_ASAP7_75t_L g2654 ( 
.A(n_2438),
.B(n_2128),
.Y(n_2654)
);

AO22x2_ASAP7_75t_L g2655 ( 
.A1(n_2351),
.A2(n_2209),
.B1(n_2224),
.B2(n_2136),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2522),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2387),
.B(n_2258),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2514),
.B(n_2292),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2387),
.B(n_2379),
.Y(n_2659)
);

CKINVDCx20_ASAP7_75t_R g2660 ( 
.A(n_2460),
.Y(n_2660)
);

NOR2x1p5_ASAP7_75t_L g2661 ( 
.A(n_2465),
.B(n_2352),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2316),
.B(n_2182),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_2368),
.B(n_1191),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2316),
.B(n_2182),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2531),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2532),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2542),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2543),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2497),
.Y(n_2669)
);

NAND2x1p5_ASAP7_75t_L g2670 ( 
.A(n_2515),
.B(n_2063),
.Y(n_2670)
);

NAND2x1_ASAP7_75t_L g2671 ( 
.A(n_2544),
.B(n_2264),
.Y(n_2671)
);

AO22x2_ASAP7_75t_L g2672 ( 
.A1(n_2450),
.A2(n_2227),
.B1(n_2233),
.B2(n_2224),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2455),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2389),
.Y(n_2674)
);

BUFx8_ASAP7_75t_L g2675 ( 
.A(n_2545),
.Y(n_2675)
);

AO22x2_ASAP7_75t_L g2676 ( 
.A1(n_2450),
.A2(n_2233),
.B1(n_2260),
.B2(n_2227),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2500),
.Y(n_2677)
);

INVx6_ASAP7_75t_L g2678 ( 
.A(n_2383),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2502),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2368),
.B(n_1191),
.Y(n_2680)
);

AO22x2_ASAP7_75t_L g2681 ( 
.A1(n_2358),
.A2(n_2260),
.B1(n_2050),
.B2(n_2115),
.Y(n_2681)
);

BUFx8_ASAP7_75t_L g2682 ( 
.A(n_2545),
.Y(n_2682)
);

AO22x2_ASAP7_75t_L g2683 ( 
.A1(n_2330),
.A2(n_2050),
.B1(n_2115),
.B2(n_2048),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2514),
.B(n_2119),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2372),
.B(n_2179),
.Y(n_2685)
);

AO22x2_ASAP7_75t_L g2686 ( 
.A1(n_2324),
.A2(n_2050),
.B1(n_2115),
.B2(n_2048),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2411),
.B(n_2481),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2431),
.B(n_2122),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2509),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2318),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2516),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2519),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2322),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2372),
.B(n_1211),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2523),
.B(n_2119),
.Y(n_2695)
);

AO22x1_ASAP7_75t_L g2696 ( 
.A1(n_2398),
.A2(n_2536),
.B1(n_2479),
.B2(n_2507),
.Y(n_2696)
);

AOI22xp5_ASAP7_75t_L g2697 ( 
.A1(n_2479),
.A2(n_1218),
.B1(n_1222),
.B2(n_1211),
.Y(n_2697)
);

AO22x2_ASAP7_75t_L g2698 ( 
.A1(n_2380),
.A2(n_2140),
.B1(n_2048),
.B2(n_2031),
.Y(n_2698)
);

AND2x2_ASAP7_75t_SL g2699 ( 
.A(n_2454),
.B(n_2217),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2538),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2534),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2391),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2335),
.Y(n_2703)
);

OAI221xp5_ASAP7_75t_L g2704 ( 
.A1(n_2454),
.A2(n_2329),
.B1(n_2503),
.B2(n_2536),
.C(n_2362),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2448),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2451),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2484),
.A2(n_1222),
.B1(n_1230),
.B2(n_1218),
.Y(n_2707)
);

AO22x2_ASAP7_75t_L g2708 ( 
.A1(n_2427),
.A2(n_2140),
.B1(n_2031),
.B2(n_2082),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2467),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2476),
.Y(n_2710)
);

AOI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2484),
.A2(n_1231),
.B1(n_1236),
.B2(n_1230),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2478),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2480),
.Y(n_2713)
);

AO22x2_ASAP7_75t_L g2714 ( 
.A1(n_2427),
.A2(n_2140),
.B1(n_2082),
.B2(n_2043),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2345),
.B(n_2122),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2488),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2495),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2340),
.B(n_2189),
.Y(n_2718)
);

AO22x2_ASAP7_75t_L g2719 ( 
.A1(n_2487),
.A2(n_2043),
.B1(n_2245),
.B2(n_2281),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2348),
.Y(n_2720)
);

AO22x2_ASAP7_75t_L g2721 ( 
.A1(n_2336),
.A2(n_2245),
.B1(n_2287),
.B2(n_2293),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2539),
.Y(n_2722)
);

OAI221xp5_ASAP7_75t_L g2723 ( 
.A1(n_2503),
.A2(n_1118),
.B1(n_1117),
.B2(n_1046),
.C(n_2212),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2339),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2339),
.Y(n_2725)
);

NAND2x1p5_ASAP7_75t_L g2726 ( 
.A(n_2544),
.B(n_2067),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2541),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2461),
.Y(n_2728)
);

NAND2x1p5_ASAP7_75t_L g2729 ( 
.A(n_2544),
.B(n_2067),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2346),
.B(n_2173),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2461),
.Y(n_2731)
);

AO22x2_ASAP7_75t_L g2732 ( 
.A1(n_2360),
.A2(n_2370),
.B1(n_2408),
.B2(n_2406),
.Y(n_2732)
);

AO22x2_ASAP7_75t_L g2733 ( 
.A1(n_2360),
.A2(n_2307),
.B1(n_2295),
.B2(n_2263),
.Y(n_2733)
);

OR2x6_ASAP7_75t_SL g2734 ( 
.A(n_2350),
.B(n_2147),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2364),
.B(n_2236),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2397),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2496),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2440),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2443),
.Y(n_2739)
);

OAI22xp5_ASAP7_75t_L g2740 ( 
.A1(n_2361),
.A2(n_2190),
.B1(n_2181),
.B2(n_2089),
.Y(n_2740)
);

AO22x2_ASAP7_75t_L g2741 ( 
.A1(n_2344),
.A2(n_2265),
.B1(n_2298),
.B2(n_2262),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2393),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2550),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2400),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2401),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2397),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2483),
.Y(n_2747)
);

AND2x4_ASAP7_75t_L g2748 ( 
.A(n_2525),
.B(n_2067),
.Y(n_2748)
);

AO22x2_ASAP7_75t_L g2749 ( 
.A1(n_2332),
.A2(n_2265),
.B1(n_2282),
.B2(n_2310),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2486),
.Y(n_2750)
);

AO22x2_ASAP7_75t_L g2751 ( 
.A1(n_2425),
.A2(n_2282),
.B1(n_2177),
.B2(n_2170),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_SL g2752 ( 
.A(n_2556),
.B(n_1742),
.Y(n_2752)
);

AO32x1_ASAP7_75t_L g2753 ( 
.A1(n_2740),
.A2(n_1018),
.A3(n_2555),
.B1(n_2459),
.B2(n_2363),
.Y(n_2753)
);

OAI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2630),
.A2(n_2376),
.B(n_2386),
.Y(n_2754)
);

BUFx2_ASAP7_75t_SL g2755 ( 
.A(n_2564),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2735),
.A2(n_2285),
.B(n_2319),
.Y(n_2756)
);

AOI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2688),
.A2(n_2235),
.B(n_2139),
.Y(n_2757)
);

INVx5_ASAP7_75t_L g2758 ( 
.A(n_2585),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2624),
.B(n_2588),
.Y(n_2759)
);

OAI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2704),
.A2(n_2680),
.B1(n_2694),
.B2(n_2663),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2659),
.B(n_2492),
.Y(n_2761)
);

OAI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2574),
.A2(n_2415),
.B1(n_2340),
.B2(n_2530),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2739),
.A2(n_2242),
.B(n_2105),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2715),
.A2(n_2118),
.B(n_2331),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2705),
.B(n_2349),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2557),
.Y(n_2766)
);

O2A1O1Ixp33_ASAP7_75t_L g2767 ( 
.A1(n_2576),
.A2(n_2551),
.B(n_2392),
.C(n_2395),
.Y(n_2767)
);

OAI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2575),
.A2(n_2415),
.B1(n_2508),
.B2(n_2537),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2607),
.A2(n_2359),
.B(n_2181),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2706),
.B(n_2349),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2654),
.B(n_2551),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2709),
.B(n_2492),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2751),
.A2(n_2089),
.B(n_2426),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2700),
.B(n_1231),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2751),
.A2(n_2428),
.B(n_2446),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_2699),
.A2(n_2498),
.B1(n_2507),
.B2(n_2508),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2640),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_SL g2778 ( 
.A(n_2710),
.B(n_2456),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2743),
.B(n_1236),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_SL g2780 ( 
.A(n_2566),
.B(n_1742),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2712),
.B(n_2713),
.Y(n_2781)
);

O2A1O1Ixp33_ASAP7_75t_L g2782 ( 
.A1(n_2622),
.A2(n_2498),
.B(n_2447),
.C(n_2462),
.Y(n_2782)
);

AO21x1_ASAP7_75t_L g2783 ( 
.A1(n_2582),
.A2(n_2737),
.B(n_2421),
.Y(n_2783)
);

OA21x2_ASAP7_75t_L g2784 ( 
.A1(n_2742),
.A2(n_1545),
.B(n_1527),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2593),
.A2(n_2546),
.B1(n_2501),
.B2(n_2416),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2669),
.A2(n_2446),
.B(n_2378),
.Y(n_2786)
);

OAI22xp5_ASAP7_75t_L g2787 ( 
.A1(n_2646),
.A2(n_2546),
.B1(n_2501),
.B2(n_2418),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2573),
.A2(n_2315),
.B1(n_2423),
.B2(n_1240),
.Y(n_2788)
);

O2A1O1Ixp33_ASAP7_75t_L g2789 ( 
.A1(n_2723),
.A2(n_2547),
.B(n_2553),
.C(n_2388),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2716),
.B(n_2413),
.Y(n_2790)
);

OAI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2560),
.A2(n_2439),
.B(n_2435),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2571),
.Y(n_2792)
);

NOR2xp67_ASAP7_75t_L g2793 ( 
.A(n_2563),
.B(n_2472),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2572),
.B(n_2619),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_L g2795 ( 
.A(n_2595),
.B(n_1238),
.Y(n_2795)
);

AOI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2677),
.A2(n_2382),
.B(n_2377),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2606),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2623),
.Y(n_2798)
);

O2A1O1Ixp33_ASAP7_75t_L g2799 ( 
.A1(n_2685),
.A2(n_2511),
.B(n_2518),
.C(n_2457),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2558),
.Y(n_2800)
);

AOI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2657),
.A2(n_1169),
.B1(n_1171),
.B2(n_1168),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2717),
.B(n_2702),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2679),
.B(n_2341),
.Y(n_2803)
);

INVxp67_ASAP7_75t_L g2804 ( 
.A(n_2567),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2689),
.A2(n_2390),
.B(n_2190),
.Y(n_2805)
);

OAI22xp5_ASAP7_75t_L g2806 ( 
.A1(n_2596),
.A2(n_2315),
.B1(n_1956),
.B2(n_2311),
.Y(n_2806)
);

AOI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2691),
.A2(n_2548),
.B(n_2074),
.Y(n_2807)
);

OAI21xp5_ASAP7_75t_L g2808 ( 
.A1(n_2634),
.A2(n_2420),
.B(n_2432),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2692),
.A2(n_2074),
.B(n_2423),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2633),
.A2(n_2315),
.B1(n_1240),
.B2(n_1245),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2701),
.A2(n_2191),
.B(n_2051),
.Y(n_2811)
);

AOI21xp5_ASAP7_75t_L g2812 ( 
.A1(n_2732),
.A2(n_2191),
.B(n_2051),
.Y(n_2812)
);

BUFx2_ASAP7_75t_L g2813 ( 
.A(n_2572),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2581),
.B(n_2417),
.Y(n_2814)
);

NOR2x1p5_ASAP7_75t_SL g2815 ( 
.A(n_2744),
.B(n_2158),
.Y(n_2815)
);

OAI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2583),
.A2(n_1245),
.B1(n_1246),
.B2(n_1238),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2732),
.A2(n_2191),
.B(n_2051),
.Y(n_2817)
);

A2O1A1Ixp33_ASAP7_75t_L g2818 ( 
.A1(n_2653),
.A2(n_2466),
.B(n_2475),
.C(n_2463),
.Y(n_2818)
);

OAI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2597),
.A2(n_1257),
.B1(n_1258),
.B2(n_1246),
.Y(n_2819)
);

OAI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2649),
.A2(n_2442),
.B(n_2437),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2722),
.B(n_2485),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2559),
.Y(n_2822)
);

AOI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2609),
.A2(n_2203),
.B(n_2191),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2561),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_L g2825 ( 
.A(n_2696),
.B(n_1257),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2641),
.B(n_1258),
.Y(n_2826)
);

HB1xp67_ASAP7_75t_L g2827 ( 
.A(n_2673),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_2612),
.B(n_2628),
.Y(n_2828)
);

OAI321xp33_ASAP7_75t_L g2829 ( 
.A1(n_2697),
.A2(n_2473),
.A3(n_2475),
.B1(n_2466),
.B2(n_2463),
.C(n_1071),
.Y(n_2829)
);

NOR2xp67_ASAP7_75t_L g2830 ( 
.A(n_2578),
.B(n_2554),
.Y(n_2830)
);

O2A1O1Ixp33_ASAP7_75t_L g2831 ( 
.A1(n_2718),
.A2(n_1620),
.B(n_1621),
.C(n_1617),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2707),
.B(n_1262),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2609),
.A2(n_2203),
.B(n_2274),
.Y(n_2833)
);

INVx2_ASAP7_75t_SL g2834 ( 
.A(n_2569),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2711),
.B(n_1262),
.Y(n_2835)
);

O2A1O1Ixp33_ASAP7_75t_L g2836 ( 
.A1(n_2661),
.A2(n_1630),
.B(n_1621),
.C(n_2430),
.Y(n_2836)
);

OAI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2745),
.A2(n_2166),
.B(n_2289),
.Y(n_2837)
);

A2O1A1Ixp33_ASAP7_75t_L g2838 ( 
.A1(n_2747),
.A2(n_2174),
.B(n_2289),
.C(n_2436),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_2584),
.B(n_1270),
.Y(n_2839)
);

A2O1A1Ixp33_ASAP7_75t_L g2840 ( 
.A1(n_2750),
.A2(n_2658),
.B(n_2738),
.C(n_2727),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2637),
.B(n_2485),
.Y(n_2841)
);

OAI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2662),
.A2(n_1545),
.B(n_2288),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_2644),
.B(n_2206),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2619),
.B(n_2468),
.Y(n_2844)
);

OAI21xp33_ASAP7_75t_L g2845 ( 
.A1(n_2573),
.A2(n_1274),
.B(n_1270),
.Y(n_2845)
);

INVx2_ASAP7_75t_SL g2846 ( 
.A(n_2616),
.Y(n_2846)
);

OAI21xp33_ASAP7_75t_L g2847 ( 
.A1(n_2724),
.A2(n_1275),
.B(n_1274),
.Y(n_2847)
);

NOR3xp33_ASAP7_75t_L g2848 ( 
.A(n_2730),
.B(n_1593),
.C(n_1582),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_SL g2849 ( 
.A(n_2644),
.B(n_2206),
.Y(n_2849)
);

O2A1O1Ixp33_ASAP7_75t_L g2850 ( 
.A1(n_2664),
.A2(n_1630),
.B(n_2441),
.C(n_1276),
.Y(n_2850)
);

A2O1A1Ixp33_ASAP7_75t_L g2851 ( 
.A1(n_2658),
.A2(n_1505),
.B(n_1507),
.C(n_1503),
.Y(n_2851)
);

INVx5_ASAP7_75t_L g2852 ( 
.A(n_2678),
.Y(n_2852)
);

CKINVDCx8_ASAP7_75t_R g2853 ( 
.A(n_2636),
.Y(n_2853)
);

INVx2_ASAP7_75t_SL g2854 ( 
.A(n_2678),
.Y(n_2854)
);

OR2x2_ASAP7_75t_L g2855 ( 
.A(n_2725),
.B(n_2485),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2650),
.B(n_1444),
.Y(n_2856)
);

BUFx2_ASAP7_75t_L g2857 ( 
.A(n_2577),
.Y(n_2857)
);

BUFx4f_ASAP7_75t_L g2858 ( 
.A(n_2636),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2617),
.A2(n_1169),
.B1(n_1171),
.B2(n_1168),
.Y(n_2859)
);

A2O1A1Ixp33_ASAP7_75t_L g2860 ( 
.A1(n_2586),
.A2(n_1505),
.B(n_1507),
.C(n_1503),
.Y(n_2860)
);

INVx2_ASAP7_75t_SL g2861 ( 
.A(n_2674),
.Y(n_2861)
);

OAI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2734),
.A2(n_1276),
.B1(n_1287),
.B2(n_1275),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2617),
.B(n_1444),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2728),
.B(n_1451),
.Y(n_2864)
);

AOI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2681),
.A2(n_2203),
.B(n_2274),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2562),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2565),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2684),
.B(n_2226),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2731),
.B(n_1451),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2687),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2592),
.B(n_1287),
.Y(n_2871)
);

OAI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2639),
.A2(n_1295),
.B1(n_1293),
.B2(n_2254),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2681),
.A2(n_2203),
.B(n_2274),
.Y(n_2873)
);

NAND2xp33_ASAP7_75t_L g2874 ( 
.A(n_2579),
.B(n_2544),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2568),
.B(n_1483),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2684),
.B(n_2086),
.Y(n_2876)
);

AOI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2672),
.A2(n_2277),
.B(n_2274),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2660),
.A2(n_1295),
.B1(n_1293),
.B2(n_1732),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2672),
.A2(n_2277),
.B(n_2240),
.Y(n_2879)
);

NAND2xp33_ASAP7_75t_L g2880 ( 
.A(n_2604),
.B(n_2086),
.Y(n_2880)
);

BUFx3_ASAP7_75t_L g2881 ( 
.A(n_2687),
.Y(n_2881)
);

AOI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2676),
.A2(n_2277),
.B(n_2240),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_2695),
.B(n_2226),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2570),
.B(n_1483),
.Y(n_2884)
);

OAI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2720),
.A2(n_2183),
.B(n_2254),
.Y(n_2885)
);

INVx11_ASAP7_75t_L g2886 ( 
.A(n_2675),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2580),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2589),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2590),
.Y(n_2889)
);

OR2x2_ASAP7_75t_L g2890 ( 
.A(n_2591),
.B(n_796),
.Y(n_2890)
);

BUFx2_ASAP7_75t_L g2891 ( 
.A(n_2748),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2594),
.Y(n_2892)
);

INVx4_ASAP7_75t_L g2893 ( 
.A(n_2643),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2598),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2748),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2676),
.A2(n_2277),
.B(n_2215),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2690),
.B(n_2471),
.Y(n_2897)
);

INVx11_ASAP7_75t_L g2898 ( 
.A(n_2675),
.Y(n_2898)
);

INVx8_ASAP7_75t_L g2899 ( 
.A(n_2695),
.Y(n_2899)
);

OAI321xp33_ASAP7_75t_L g2900 ( 
.A1(n_2631),
.A2(n_1073),
.A3(n_1072),
.B1(n_1063),
.B2(n_812),
.C(n_1582),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2693),
.B(n_1593),
.Y(n_2901)
);

AOI21xp33_ASAP7_75t_L g2902 ( 
.A1(n_2719),
.A2(n_1301),
.B(n_2215),
.Y(n_2902)
);

A2O1A1Ixp33_ASAP7_75t_L g2903 ( 
.A1(n_2632),
.A2(n_1519),
.B(n_1522),
.C(n_1509),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2703),
.B(n_1616),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2736),
.B(n_1732),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2603),
.A2(n_2505),
.B(n_2482),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2746),
.B(n_1301),
.Y(n_2907)
);

AND2x4_ASAP7_75t_L g2908 ( 
.A(n_2599),
.B(n_2086),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2600),
.Y(n_2909)
);

AOI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2603),
.A2(n_2505),
.B(n_2482),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2629),
.A2(n_2275),
.B(n_2032),
.Y(n_2911)
);

BUFx6f_ASAP7_75t_L g2912 ( 
.A(n_2726),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2729),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2629),
.A2(n_2655),
.B(n_2733),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2601),
.B(n_1616),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2602),
.B(n_1858),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2605),
.B(n_1509),
.Y(n_2917)
);

AOI22xp33_ASAP7_75t_L g2918 ( 
.A1(n_2719),
.A2(n_2721),
.B1(n_2655),
.B2(n_2615),
.Y(n_2918)
);

AO32x1_ASAP7_75t_L g2919 ( 
.A1(n_2635),
.A2(n_2459),
.A3(n_2363),
.B1(n_2158),
.B2(n_2199),
.Y(n_2919)
);

INVx2_ASAP7_75t_SL g2920 ( 
.A(n_2682),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2670),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2733),
.A2(n_2275),
.B(n_2032),
.Y(n_2922)
);

AOI22xp33_ASAP7_75t_L g2923 ( 
.A1(n_2721),
.A2(n_1860),
.B1(n_1866),
.B2(n_1858),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2608),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_SL g2925 ( 
.A(n_2610),
.B(n_1860),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2611),
.B(n_1519),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2613),
.B(n_1522),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2587),
.A2(n_1866),
.B1(n_2033),
.B2(n_2086),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2614),
.B(n_2064),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2618),
.B(n_563),
.Y(n_2930)
);

O2A1O1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2638),
.A2(n_942),
.B(n_1029),
.C(n_1028),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2620),
.Y(n_2932)
);

BUFx8_ASAP7_75t_L g2933 ( 
.A(n_2682),
.Y(n_2933)
);

INVx3_ASAP7_75t_L g2934 ( 
.A(n_2645),
.Y(n_2934)
);

OR2x6_ASAP7_75t_L g2935 ( 
.A(n_2683),
.B(n_2033),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2621),
.B(n_2001),
.Y(n_2936)
);

AOI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2749),
.A2(n_1527),
.B(n_2171),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2626),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2587),
.A2(n_2033),
.B1(n_2219),
.B2(n_2002),
.Y(n_2939)
);

OAI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2627),
.A2(n_2239),
.B(n_2160),
.Y(n_2940)
);

AND2x6_ASAP7_75t_L g2941 ( 
.A(n_2642),
.B(n_2323),
.Y(n_2941)
);

AOI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2741),
.A2(n_2038),
.B(n_2022),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2647),
.B(n_2070),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2756),
.A2(n_2741),
.B(n_2686),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2766),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2754),
.A2(n_2686),
.B(n_2683),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2796),
.A2(n_2625),
.B(n_2615),
.Y(n_2947)
);

AOI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2760),
.A2(n_2625),
.B1(n_2749),
.B2(n_2002),
.Y(n_2948)
);

AO21x1_ASAP7_75t_L g2949 ( 
.A1(n_2771),
.A2(n_2651),
.B(n_2648),
.Y(n_2949)
);

O2A1O1Ixp33_ASAP7_75t_L g2950 ( 
.A1(n_2845),
.A2(n_2656),
.B(n_2665),
.C(n_2652),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_R g2951 ( 
.A(n_2780),
.B(n_2001),
.Y(n_2951)
);

INVxp67_ASAP7_75t_L g2952 ( 
.A(n_2827),
.Y(n_2952)
);

BUFx6f_ASAP7_75t_L g2953 ( 
.A(n_2852),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2800),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2776),
.A2(n_2698),
.B1(n_2714),
.B2(n_2708),
.Y(n_2955)
);

NAND2x1p5_ASAP7_75t_L g2956 ( 
.A(n_2758),
.B(n_2323),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2887),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2822),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2769),
.A2(n_2708),
.B(n_2714),
.Y(n_2959)
);

O2A1O1Ixp33_ASAP7_75t_L g2960 ( 
.A1(n_2828),
.A2(n_2667),
.B(n_2668),
.C(n_2666),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2761),
.B(n_595),
.Y(n_2961)
);

AOI22xp5_ASAP7_75t_L g2962 ( 
.A1(n_2825),
.A2(n_2159),
.B1(n_2698),
.B2(n_889),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2764),
.A2(n_2671),
.B(n_2645),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2759),
.B(n_2774),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2772),
.B(n_1542),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2781),
.B(n_1542),
.Y(n_2966)
);

INVx4_ASAP7_75t_L g2967 ( 
.A(n_2852),
.Y(n_2967)
);

INVx1_ASAP7_75t_SL g2968 ( 
.A(n_2857),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2879),
.A2(n_2671),
.B(n_2038),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2765),
.B(n_1032),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2832),
.A2(n_2835),
.B1(n_2795),
.B2(n_2848),
.Y(n_2971)
);

OAI22x1_ASAP7_75t_L g2972 ( 
.A1(n_2778),
.A2(n_751),
.B1(n_753),
.B2(n_750),
.Y(n_2972)
);

A2O1A1Ixp33_ASAP7_75t_L g2973 ( 
.A1(n_2767),
.A2(n_491),
.B(n_493),
.C(n_490),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2824),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2777),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_2779),
.B(n_2159),
.Y(n_2976)
);

BUFx3_ASAP7_75t_L g2977 ( 
.A(n_2852),
.Y(n_2977)
);

OAI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2850),
.A2(n_2239),
.B(n_1628),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2839),
.B(n_490),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2882),
.A2(n_2022),
.B(n_2266),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2770),
.B(n_1034),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2802),
.B(n_1036),
.Y(n_2982)
);

BUFx6f_ASAP7_75t_L g2983 ( 
.A(n_2858),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2866),
.Y(n_2984)
);

INVx2_ASAP7_75t_SL g2985 ( 
.A(n_2758),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2896),
.A2(n_2266),
.B(n_2267),
.Y(n_2986)
);

INVx3_ASAP7_75t_L g2987 ( 
.A(n_2895),
.Y(n_2987)
);

A2O1A1Ixp33_ASAP7_75t_L g2988 ( 
.A1(n_2782),
.A2(n_493),
.B(n_494),
.C(n_491),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2799),
.B(n_2785),
.Y(n_2989)
);

AND2x4_ASAP7_75t_L g2990 ( 
.A(n_2876),
.B(n_2323),
.Y(n_2990)
);

BUFx8_ASAP7_75t_L g2991 ( 
.A(n_2920),
.Y(n_2991)
);

INVxp67_ASAP7_75t_L g2992 ( 
.A(n_2870),
.Y(n_2992)
);

OAI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2788),
.A2(n_753),
.B1(n_754),
.B2(n_751),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2867),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2792),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_SL g2996 ( 
.A(n_2787),
.B(n_2323),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2803),
.B(n_1037),
.Y(n_2997)
);

NAND2x1p5_ASAP7_75t_L g2998 ( 
.A(n_2758),
.B(n_2328),
.Y(n_2998)
);

NOR2xp33_ASAP7_75t_SL g2999 ( 
.A(n_2752),
.B(n_2328),
.Y(n_2999)
);

AOI21x1_ASAP7_75t_L g3000 ( 
.A1(n_2812),
.A2(n_1042),
.B(n_1041),
.Y(n_3000)
);

OAI21xp33_ASAP7_75t_L g3001 ( 
.A1(n_2768),
.A2(n_756),
.B(n_754),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2797),
.Y(n_3002)
);

OAI22xp5_ASAP7_75t_L g3003 ( 
.A1(n_2923),
.A2(n_2801),
.B1(n_2762),
.B2(n_2806),
.Y(n_3003)
);

BUFx6f_ASAP7_75t_L g3004 ( 
.A(n_2858),
.Y(n_3004)
);

A2O1A1Ixp33_ASAP7_75t_L g3005 ( 
.A1(n_2789),
.A2(n_495),
.B(n_499),
.C(n_494),
.Y(n_3005)
);

BUFx12f_ASAP7_75t_L g3006 ( 
.A(n_2933),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2794),
.B(n_595),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2790),
.B(n_1045),
.Y(n_3008)
);

O2A1O1Ixp5_ASAP7_75t_L g3009 ( 
.A1(n_2783),
.A2(n_2037),
.B(n_2094),
.C(n_2034),
.Y(n_3009)
);

OAI22x1_ASAP7_75t_L g3010 ( 
.A1(n_2859),
.A2(n_758),
.B1(n_756),
.B2(n_499),
.Y(n_3010)
);

AOI22xp5_ASAP7_75t_L g3011 ( 
.A1(n_2826),
.A2(n_889),
.B1(n_758),
.B2(n_500),
.Y(n_3011)
);

BUFx2_ASAP7_75t_L g3012 ( 
.A(n_2813),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2804),
.B(n_2171),
.Y(n_3013)
);

INVxp67_ASAP7_75t_SL g3014 ( 
.A(n_2938),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2871),
.B(n_495),
.Y(n_3015)
);

AOI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2757),
.A2(n_2272),
.B(n_2267),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2888),
.Y(n_3017)
);

OAI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2878),
.A2(n_2280),
.B1(n_2230),
.B2(n_2238),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2889),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_SL g3020 ( 
.A(n_2853),
.B(n_2328),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2805),
.A2(n_2272),
.B(n_2328),
.Y(n_3021)
);

A2O1A1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2829),
.A2(n_500),
.B(n_712),
.C(n_707),
.Y(n_3022)
);

AOI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2862),
.A2(n_889),
.B1(n_707),
.B2(n_721),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2816),
.B(n_2819),
.Y(n_3024)
);

AOI21x1_ASAP7_75t_L g3025 ( 
.A1(n_2817),
.A2(n_2199),
.B(n_2176),
.Y(n_3025)
);

AOI221xp5_ASAP7_75t_L g3026 ( 
.A1(n_2902),
.A2(n_722),
.B1(n_741),
.B2(n_721),
.C(n_712),
.Y(n_3026)
);

CKINVDCx5p33_ASAP7_75t_R g3027 ( 
.A(n_2933),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2877),
.A2(n_2807),
.B(n_2763),
.Y(n_3028)
);

OR2x6_ASAP7_75t_L g3029 ( 
.A(n_2935),
.B(n_2914),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2814),
.B(n_2176),
.Y(n_3030)
);

INVx3_ASAP7_75t_L g3031 ( 
.A(n_2895),
.Y(n_3031)
);

AOI22xp5_ASAP7_75t_L g3032 ( 
.A1(n_2847),
.A2(n_733),
.B1(n_595),
.B2(n_722),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2794),
.B(n_733),
.Y(n_3033)
);

A2O1A1Ixp33_ASAP7_75t_L g3034 ( 
.A1(n_2840),
.A2(n_742),
.B(n_743),
.C(n_741),
.Y(n_3034)
);

XNOR2xp5_ASAP7_75t_L g3035 ( 
.A(n_2810),
.B(n_742),
.Y(n_3035)
);

HB1xp67_ASAP7_75t_L g3036 ( 
.A(n_2891),
.Y(n_3036)
);

A2O1A1Ixp33_ASAP7_75t_L g3037 ( 
.A1(n_2836),
.A2(n_743),
.B(n_509),
.C(n_517),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2798),
.B(n_2214),
.Y(n_3038)
);

AO32x2_ASAP7_75t_L g3039 ( 
.A1(n_2939),
.A2(n_498),
.A3(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2786),
.A2(n_2394),
.B(n_2373),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2881),
.Y(n_3041)
);

HB1xp67_ASAP7_75t_L g3042 ( 
.A(n_2892),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2809),
.A2(n_2394),
.B(n_2373),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2880),
.A2(n_2394),
.B(n_2373),
.Y(n_3044)
);

O2A1O1Ixp33_ASAP7_75t_L g3045 ( 
.A1(n_2925),
.A2(n_892),
.B(n_915),
.C(n_894),
.Y(n_3045)
);

INVxp67_ASAP7_75t_L g3046 ( 
.A(n_2905),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_SL g3047 ( 
.A(n_2821),
.B(n_2373),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2856),
.B(n_2214),
.Y(n_3048)
);

AOI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_2916),
.A2(n_733),
.B1(n_525),
.B2(n_529),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2894),
.Y(n_3050)
);

O2A1O1Ixp33_ASAP7_75t_L g3051 ( 
.A1(n_2851),
.A2(n_915),
.B(n_927),
.C(n_894),
.Y(n_3051)
);

BUFx6f_ASAP7_75t_L g3052 ( 
.A(n_2895),
.Y(n_3052)
);

AND2x2_ASAP7_75t_SL g3053 ( 
.A(n_2874),
.B(n_2394),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2909),
.B(n_2222),
.Y(n_3054)
);

OAI21x1_ASAP7_75t_L g3055 ( 
.A1(n_2937),
.A2(n_2243),
.B(n_2222),
.Y(n_3055)
);

O2A1O1Ixp33_ASAP7_75t_L g3056 ( 
.A1(n_2872),
.A2(n_929),
.B(n_932),
.C(n_927),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_2834),
.Y(n_3057)
);

AOI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2865),
.A2(n_2280),
.B(n_2037),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2924),
.Y(n_3059)
);

HB1xp67_ASAP7_75t_L g3060 ( 
.A(n_2932),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2863),
.B(n_2243),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2875),
.B(n_2247),
.Y(n_3062)
);

NOR2xp33_ASAP7_75t_L g3063 ( 
.A(n_2936),
.B(n_512),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2793),
.B(n_2273),
.Y(n_3064)
);

A2O1A1Ixp33_ASAP7_75t_L g3065 ( 
.A1(n_2900),
.A2(n_531),
.B(n_550),
.C(n_530),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2943),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2873),
.A2(n_2094),
.B(n_2034),
.Y(n_3067)
);

A2O1A1Ixp33_ASAP7_75t_SL g3068 ( 
.A1(n_2791),
.A2(n_1531),
.B(n_1525),
.C(n_2211),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2841),
.B(n_929),
.Y(n_3069)
);

OAI22xp5_ASAP7_75t_L g3070 ( 
.A1(n_2897),
.A2(n_2152),
.B1(n_2172),
.B2(n_2145),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2855),
.B(n_2808),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2833),
.A2(n_2152),
.B(n_2145),
.Y(n_3072)
);

AOI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2773),
.A2(n_2252),
.B(n_2247),
.Y(n_3073)
);

OAI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2838),
.A2(n_2239),
.B(n_2252),
.Y(n_3074)
);

BUFx6f_ASAP7_75t_L g3075 ( 
.A(n_2846),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_R g3076 ( 
.A(n_2854),
.B(n_2273),
.Y(n_3076)
);

AOI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2775),
.A2(n_2180),
.B(n_2172),
.Y(n_3077)
);

AOI31xp33_ASAP7_75t_L g3078 ( 
.A1(n_2843),
.A2(n_558),
.A3(n_566),
.B(n_552),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2908),
.Y(n_3079)
);

O2A1O1Ixp33_ASAP7_75t_L g3080 ( 
.A1(n_2818),
.A2(n_932),
.B(n_2180),
.C(n_1531),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2907),
.B(n_570),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2884),
.B(n_2239),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2885),
.A2(n_2296),
.B(n_2273),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2930),
.B(n_571),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2823),
.A2(n_2296),
.B(n_1462),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2864),
.B(n_2239),
.Y(n_3086)
);

O2A1O1Ixp33_ASAP7_75t_L g3087 ( 
.A1(n_2883),
.A2(n_1531),
.B(n_1525),
.C(n_1482),
.Y(n_3087)
);

BUFx2_ASAP7_75t_L g3088 ( 
.A(n_2899),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_2861),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2837),
.A2(n_2296),
.B(n_1455),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2940),
.A2(n_2296),
.B(n_1525),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2919),
.A2(n_1482),
.B(n_1479),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2830),
.B(n_1528),
.Y(n_3093)
);

CKINVDCx5p33_ASAP7_75t_R g3094 ( 
.A(n_2886),
.Y(n_3094)
);

O2A1O1Ixp33_ASAP7_75t_L g3095 ( 
.A1(n_2860),
.A2(n_1485),
.B(n_1491),
.C(n_1490),
.Y(n_3095)
);

CKINVDCx5p33_ASAP7_75t_R g3096 ( 
.A(n_2898),
.Y(n_3096)
);

A2O1A1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2831),
.A2(n_574),
.B(n_575),
.C(n_573),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2869),
.B(n_576),
.Y(n_3098)
);

OAI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2820),
.A2(n_593),
.B(n_580),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2919),
.A2(n_1490),
.B(n_1485),
.Y(n_3100)
);

CKINVDCx5p33_ASAP7_75t_R g3101 ( 
.A(n_2755),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2929),
.Y(n_3102)
);

INVx1_ASAP7_75t_SL g3103 ( 
.A(n_2890),
.Y(n_3103)
);

AND2x4_ASAP7_75t_L g3104 ( 
.A(n_2876),
.B(n_231),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2908),
.Y(n_3105)
);

CKINVDCx16_ASAP7_75t_R g3106 ( 
.A(n_2844),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2919),
.A2(n_1494),
.B(n_1491),
.Y(n_3107)
);

XNOR2xp5_ASAP7_75t_L g3108 ( 
.A(n_2844),
.B(n_596),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_2935),
.Y(n_3109)
);

AOI22xp5_ASAP7_75t_L g3110 ( 
.A1(n_2849),
.A2(n_623),
.B1(n_624),
.B2(n_605),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2915),
.B(n_626),
.Y(n_3111)
);

O2A1O1Ixp33_ASAP7_75t_L g3112 ( 
.A1(n_2928),
.A2(n_1512),
.B(n_1515),
.C(n_1494),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2868),
.B(n_1528),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2901),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2893),
.B(n_2921),
.Y(n_3115)
);

BUFx2_ASAP7_75t_L g3116 ( 
.A(n_2899),
.Y(n_3116)
);

AOI222xp33_ASAP7_75t_L g3117 ( 
.A1(n_2904),
.A2(n_706),
.B1(n_701),
.B2(n_698),
.C1(n_695),
.C2(n_689),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2811),
.A2(n_1515),
.B(n_1512),
.Y(n_3118)
);

NOR3xp33_ASAP7_75t_L g3119 ( 
.A(n_2931),
.B(n_651),
.C(n_648),
.Y(n_3119)
);

AND2x4_ASAP7_75t_L g3120 ( 
.A(n_2913),
.B(n_235),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2917),
.B(n_665),
.Y(n_3121)
);

NOR3xp33_ASAP7_75t_L g3122 ( 
.A(n_2903),
.B(n_672),
.C(n_670),
.Y(n_3122)
);

BUFx6f_ASAP7_75t_L g3123 ( 
.A(n_2912),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_2893),
.B(n_1528),
.Y(n_3124)
);

INVxp67_ASAP7_75t_SL g3125 ( 
.A(n_2942),
.Y(n_3125)
);

AND2x4_ASAP7_75t_L g3126 ( 
.A(n_2913),
.B(n_236),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2926),
.B(n_673),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2912),
.Y(n_3128)
);

BUFx2_ASAP7_75t_L g3129 ( 
.A(n_2912),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2927),
.B(n_675),
.Y(n_3130)
);

OAI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_2918),
.A2(n_2921),
.B1(n_2906),
.B2(n_2910),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2941),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2941),
.Y(n_3133)
);

OA21x2_ASAP7_75t_L g3134 ( 
.A1(n_2911),
.A2(n_1518),
.B(n_678),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2934),
.B(n_677),
.Y(n_3135)
);

BUFx2_ASAP7_75t_L g3136 ( 
.A(n_2941),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2941),
.A2(n_685),
.B1(n_679),
.B2(n_1535),
.Y(n_3137)
);

OAI22xp5_ASAP7_75t_L g3138 ( 
.A1(n_2934),
.A2(n_1493),
.B1(n_1498),
.B2(n_1432),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2842),
.B(n_1528),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2815),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_2922),
.B(n_237),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2784),
.B(n_238),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2784),
.Y(n_3143)
);

OAI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2753),
.A2(n_1518),
.B(n_1513),
.Y(n_3144)
);

NAND3xp33_ASAP7_75t_SL g3145 ( 
.A(n_2753),
.B(n_5),
.C(n_9),
.Y(n_3145)
);

HB1xp67_ASAP7_75t_L g3146 ( 
.A(n_2753),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2766),
.Y(n_3147)
);

BUFx6f_ASAP7_75t_L g3148 ( 
.A(n_2953),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2945),
.Y(n_3149)
);

AND2x4_ASAP7_75t_L g3150 ( 
.A(n_3109),
.B(n_239),
.Y(n_3150)
);

INVx3_ASAP7_75t_L g3151 ( 
.A(n_3123),
.Y(n_3151)
);

CKINVDCx5p33_ASAP7_75t_R g3152 ( 
.A(n_3006),
.Y(n_3152)
);

INVx1_ASAP7_75t_SL g3153 ( 
.A(n_3103),
.Y(n_3153)
);

OR2x2_ASAP7_75t_L g3154 ( 
.A(n_3042),
.B(n_776),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2953),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3147),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2954),
.Y(n_3157)
);

INVx3_ASAP7_75t_L g3158 ( 
.A(n_3123),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_3003),
.A2(n_1535),
.B1(n_1528),
.B2(n_1506),
.Y(n_3159)
);

BUFx10_ASAP7_75t_L g3160 ( 
.A(n_3027),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2958),
.Y(n_3161)
);

NAND2x1p5_ASAP7_75t_L g3162 ( 
.A(n_2967),
.B(n_1432),
.Y(n_3162)
);

INVxp67_ASAP7_75t_L g3163 ( 
.A(n_2968),
.Y(n_3163)
);

INVx4_ASAP7_75t_L g3164 ( 
.A(n_2953),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_3060),
.Y(n_3165)
);

BUFx2_ASAP7_75t_L g3166 ( 
.A(n_3036),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2974),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2984),
.Y(n_3168)
);

INVx1_ASAP7_75t_SL g3169 ( 
.A(n_3089),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_3029),
.B(n_241),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2994),
.Y(n_3171)
);

INVx1_ASAP7_75t_SL g3172 ( 
.A(n_3057),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_3014),
.B(n_10),
.Y(n_3173)
);

INVx2_ASAP7_75t_SL g3174 ( 
.A(n_3075),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3017),
.Y(n_3175)
);

INVx1_ASAP7_75t_SL g3176 ( 
.A(n_3101),
.Y(n_3176)
);

INVx3_ASAP7_75t_L g3177 ( 
.A(n_3123),
.Y(n_3177)
);

NOR2x1_ASAP7_75t_L g3178 ( 
.A(n_2989),
.B(n_776),
.Y(n_3178)
);

CKINVDCx11_ASAP7_75t_R g3179 ( 
.A(n_3075),
.Y(n_3179)
);

OR2x2_ASAP7_75t_L g3180 ( 
.A(n_2952),
.B(n_776),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3019),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3050),
.Y(n_3182)
);

OAI22xp5_ASAP7_75t_L g3183 ( 
.A1(n_2971),
.A2(n_1535),
.B1(n_1493),
.B2(n_1498),
.Y(n_3183)
);

HB1xp67_ASAP7_75t_L g3184 ( 
.A(n_3059),
.Y(n_3184)
);

HB1xp67_ASAP7_75t_L g3185 ( 
.A(n_2957),
.Y(n_3185)
);

AOI222xp33_ASAP7_75t_L g3186 ( 
.A1(n_3001),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_18),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3066),
.B(n_12),
.Y(n_3187)
);

BUFx4f_ASAP7_75t_L g3188 ( 
.A(n_2983),
.Y(n_3188)
);

INVx5_ASAP7_75t_L g3189 ( 
.A(n_2967),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2975),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3143),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3125),
.Y(n_3192)
);

OR2x6_ASAP7_75t_L g3193 ( 
.A(n_3029),
.B(n_872),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3114),
.B(n_14),
.Y(n_3194)
);

OAI22x1_ASAP7_75t_L g3195 ( 
.A1(n_2948),
.A2(n_20),
.B1(n_15),
.B2(n_18),
.Y(n_3195)
);

AND2x4_ASAP7_75t_L g3196 ( 
.A(n_3029),
.B(n_243),
.Y(n_3196)
);

BUFx4f_ASAP7_75t_L g3197 ( 
.A(n_2983),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2995),
.Y(n_3198)
);

OR2x6_ASAP7_75t_L g3199 ( 
.A(n_2946),
.B(n_872),
.Y(n_3199)
);

AND3x1_ASAP7_75t_SL g3200 ( 
.A(n_3026),
.B(n_20),
.C(n_21),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2964),
.B(n_22),
.Y(n_3201)
);

AOI221x1_ASAP7_75t_L g3202 ( 
.A1(n_2972),
.A2(n_950),
.B1(n_955),
.B2(n_900),
.C(n_872),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_3046),
.B(n_22),
.Y(n_3203)
);

BUFx12f_ASAP7_75t_L g3204 ( 
.A(n_3094),
.Y(n_3204)
);

AND2x4_ASAP7_75t_L g3205 ( 
.A(n_3136),
.B(n_245),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3032),
.A2(n_1535),
.B1(n_1493),
.B2(n_1498),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3002),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3140),
.Y(n_3208)
);

INVx3_ASAP7_75t_L g3209 ( 
.A(n_3128),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_3102),
.Y(n_3210)
);

BUFx3_ASAP7_75t_L g3211 ( 
.A(n_3075),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_3128),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_2977),
.Y(n_3213)
);

INVx1_ASAP7_75t_SL g3214 ( 
.A(n_3012),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_3079),
.Y(n_3215)
);

INVx1_ASAP7_75t_SL g3216 ( 
.A(n_3041),
.Y(n_3216)
);

INVx5_ASAP7_75t_L g3217 ( 
.A(n_3141),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3105),
.B(n_24),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_3139),
.A2(n_1535),
.B(n_1517),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2949),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_3052),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_3015),
.B(n_24),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_3129),
.B(n_25),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_3013),
.Y(n_3224)
);

BUFx6f_ASAP7_75t_L g3225 ( 
.A(n_3052),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_3052),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2999),
.B(n_1506),
.Y(n_3227)
);

INVx2_ASAP7_75t_SL g3228 ( 
.A(n_2991),
.Y(n_3228)
);

CKINVDCx20_ASAP7_75t_R g3229 ( 
.A(n_3096),
.Y(n_3229)
);

HB1xp67_ASAP7_75t_L g3230 ( 
.A(n_3071),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3024),
.B(n_25),
.Y(n_3231)
);

OAI22xp33_ASAP7_75t_L g3232 ( 
.A1(n_3032),
.A2(n_900),
.B1(n_950),
.B2(n_872),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_2983),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3035),
.A2(n_1432),
.B1(n_900),
.B2(n_950),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_3076),
.Y(n_3235)
);

BUFx2_ASAP7_75t_L g3236 ( 
.A(n_2992),
.Y(n_3236)
);

INVx2_ASAP7_75t_SL g3237 ( 
.A(n_2991),
.Y(n_3237)
);

OAI22x1_ASAP7_75t_L g3238 ( 
.A1(n_2948),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3069),
.B(n_27),
.Y(n_3239)
);

CKINVDCx11_ASAP7_75t_R g3240 ( 
.A(n_3106),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_2988),
.A2(n_1517),
.B(n_1506),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3048),
.B(n_28),
.Y(n_3242)
);

BUFx8_ASAP7_75t_L g3243 ( 
.A(n_3007),
.Y(n_3243)
);

AOI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3063),
.A2(n_1513),
.B1(n_1502),
.B2(n_1506),
.Y(n_3244)
);

NOR2xp67_ASAP7_75t_L g3245 ( 
.A(n_2985),
.B(n_3008),
.Y(n_3245)
);

BUFx3_ASAP7_75t_L g3246 ( 
.A(n_3088),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2987),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3055),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3073),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3131),
.Y(n_3250)
);

HB1xp67_ASAP7_75t_L g3251 ( 
.A(n_2996),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2961),
.B(n_29),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_3116),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2987),
.Y(n_3254)
);

BUFx6f_ASAP7_75t_L g3255 ( 
.A(n_3004),
.Y(n_3255)
);

BUFx2_ASAP7_75t_L g3256 ( 
.A(n_3132),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3054),
.Y(n_3257)
);

BUFx3_ASAP7_75t_L g3258 ( 
.A(n_3031),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2947),
.Y(n_3259)
);

AND2x4_ASAP7_75t_L g3260 ( 
.A(n_3133),
.B(n_248),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_3133),
.Y(n_3261)
);

INVxp67_ASAP7_75t_SL g3262 ( 
.A(n_2960),
.Y(n_3262)
);

BUFx6f_ASAP7_75t_L g3263 ( 
.A(n_3004),
.Y(n_3263)
);

OR2x6_ASAP7_75t_L g3264 ( 
.A(n_2959),
.B(n_872),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2950),
.Y(n_3265)
);

AOI221xp5_ASAP7_75t_L g3266 ( 
.A1(n_2993),
.A2(n_1062),
.B1(n_1050),
.B2(n_960),
.C(n_955),
.Y(n_3266)
);

A2O1A1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_2973),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3039),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_3031),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3047),
.Y(n_3270)
);

BUFx6f_ASAP7_75t_L g3271 ( 
.A(n_3004),
.Y(n_3271)
);

INVx2_ASAP7_75t_SL g3272 ( 
.A(n_2990),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_3038),
.Y(n_3273)
);

BUFx12f_ASAP7_75t_L g3274 ( 
.A(n_3033),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_2951),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_2955),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_2990),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3028),
.A2(n_1517),
.B(n_1513),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_3108),
.Y(n_3279)
);

OR2x6_ASAP7_75t_L g3280 ( 
.A(n_2944),
.B(n_900),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3146),
.Y(n_3281)
);

OAI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_3049),
.A2(n_3023),
.B1(n_3011),
.B2(n_2962),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3030),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_SL g3284 ( 
.A(n_3053),
.B(n_1517),
.Y(n_3284)
);

AOI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3119),
.A2(n_1502),
.B1(n_1517),
.B2(n_950),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3025),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3086),
.B(n_31),
.Y(n_3287)
);

AND2x4_ASAP7_75t_L g3288 ( 
.A(n_3115),
.B(n_250),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_3122),
.A2(n_1502),
.B1(n_950),
.B2(n_955),
.Y(n_3289)
);

INVx5_ASAP7_75t_L g3290 ( 
.A(n_3141),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3009),
.Y(n_3291)
);

AND2x4_ASAP7_75t_L g3292 ( 
.A(n_3043),
.B(n_251),
.Y(n_3292)
);

BUFx2_ASAP7_75t_L g3293 ( 
.A(n_2956),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3142),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2966),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_2979),
.A2(n_955),
.B1(n_960),
.B2(n_900),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3061),
.B(n_32),
.Y(n_3297)
);

BUFx12f_ASAP7_75t_L g3298 ( 
.A(n_3104),
.Y(n_3298)
);

A2O1A1Ixp33_ASAP7_75t_L g3299 ( 
.A1(n_3005),
.A2(n_3034),
.B(n_3081),
.C(n_3078),
.Y(n_3299)
);

O2A1O1Ixp33_ASAP7_75t_L g3300 ( 
.A1(n_3022),
.A2(n_38),
.B(n_35),
.C(n_36),
.Y(n_3300)
);

HB1xp67_ASAP7_75t_L g3301 ( 
.A(n_3082),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3134),
.Y(n_3302)
);

INVx1_ASAP7_75t_SL g3303 ( 
.A(n_3084),
.Y(n_3303)
);

INVx5_ASAP7_75t_L g3304 ( 
.A(n_3135),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_3104),
.B(n_252),
.Y(n_3305)
);

INVx3_ASAP7_75t_L g3306 ( 
.A(n_2998),
.Y(n_3306)
);

INVx4_ASAP7_75t_L g3307 ( 
.A(n_3120),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_3010),
.A2(n_960),
.B1(n_1050),
.B2(n_955),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_2976),
.B(n_38),
.Y(n_3309)
);

OR2x6_ASAP7_75t_L g3310 ( 
.A(n_3040),
.B(n_3083),
.Y(n_3310)
);

OAI22xp33_ASAP7_75t_SL g3311 ( 
.A1(n_3113),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3134),
.Y(n_3312)
);

BUFx6f_ASAP7_75t_L g3313 ( 
.A(n_3120),
.Y(n_3313)
);

A2O1A1Ixp33_ASAP7_75t_L g3314 ( 
.A1(n_3137),
.A2(n_44),
.B(n_39),
.C(n_40),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_3126),
.Y(n_3315)
);

BUFx2_ASAP7_75t_L g3316 ( 
.A(n_3126),
.Y(n_3316)
);

AOI21xp33_ASAP7_75t_L g3317 ( 
.A1(n_3099),
.A2(n_44),
.B(n_46),
.Y(n_3317)
);

AOI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_3117),
.A2(n_1050),
.B1(n_1062),
.B2(n_960),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_3062),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_2965),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2980),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2986),
.Y(n_3322)
);

INVxp67_ASAP7_75t_SL g3323 ( 
.A(n_2969),
.Y(n_3323)
);

AOI22xp33_ASAP7_75t_L g3324 ( 
.A1(n_2978),
.A2(n_1050),
.B1(n_1062),
.B2(n_960),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2970),
.B(n_46),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3000),
.Y(n_3326)
);

NAND2x1_ASAP7_75t_L g3327 ( 
.A(n_2963),
.B(n_1050),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3064),
.B(n_47),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2982),
.Y(n_3329)
);

INVxp67_ASAP7_75t_L g3330 ( 
.A(n_2981),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3039),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_3080),
.A2(n_1465),
.B(n_1458),
.Y(n_3332)
);

OAI22xp5_ASAP7_75t_L g3333 ( 
.A1(n_3137),
.A2(n_1062),
.B1(n_51),
.B2(n_48),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3039),
.Y(n_3334)
);

HB1xp67_ASAP7_75t_L g3335 ( 
.A(n_3074),
.Y(n_3335)
);

BUFx3_ASAP7_75t_L g3336 ( 
.A(n_3098),
.Y(n_3336)
);

BUFx2_ASAP7_75t_L g3337 ( 
.A(n_3070),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_2997),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3145),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3124),
.Y(n_3340)
);

INVxp67_ASAP7_75t_L g3341 ( 
.A(n_3111),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3093),
.Y(n_3342)
);

OAI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_3110),
.A2(n_1062),
.B1(n_53),
.B2(n_49),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3021),
.Y(n_3344)
);

BUFx6f_ASAP7_75t_L g3345 ( 
.A(n_3121),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3077),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3020),
.B(n_52),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3110),
.B(n_3018),
.Y(n_3348)
);

INVx3_ASAP7_75t_L g3349 ( 
.A(n_3127),
.Y(n_3349)
);

BUFx12f_ASAP7_75t_L g3350 ( 
.A(n_3045),
.Y(n_3350)
);

INVx4_ASAP7_75t_L g3351 ( 
.A(n_3044),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3130),
.B(n_52),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3090),
.B(n_53),
.Y(n_3353)
);

O2A1O1Ixp33_ASAP7_75t_L g3354 ( 
.A1(n_3065),
.A2(n_57),
.B(n_54),
.C(n_55),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3144),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3068),
.A2(n_1465),
.B(n_1458),
.Y(n_3356)
);

BUFx2_ASAP7_75t_L g3357 ( 
.A(n_3138),
.Y(n_3357)
);

BUFx6f_ASAP7_75t_L g3358 ( 
.A(n_3058),
.Y(n_3358)
);

BUFx6f_ASAP7_75t_L g3359 ( 
.A(n_3072),
.Y(n_3359)
);

INVx2_ASAP7_75t_SL g3360 ( 
.A(n_3067),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3056),
.B(n_54),
.Y(n_3361)
);

INVx3_ASAP7_75t_L g3362 ( 
.A(n_3261),
.Y(n_3362)
);

BUFx2_ASAP7_75t_L g3363 ( 
.A(n_3166),
.Y(n_3363)
);

BUFx2_ASAP7_75t_L g3364 ( 
.A(n_3165),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3294),
.B(n_3016),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3262),
.A2(n_3037),
.B(n_3097),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3175),
.Y(n_3367)
);

CKINVDCx20_ASAP7_75t_R g3368 ( 
.A(n_3229),
.Y(n_3368)
);

HB1xp67_ASAP7_75t_L g3369 ( 
.A(n_3230),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3149),
.Y(n_3370)
);

INVx5_ASAP7_75t_L g3371 ( 
.A(n_3193),
.Y(n_3371)
);

AND2x4_ASAP7_75t_L g3372 ( 
.A(n_3208),
.B(n_3085),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3214),
.B(n_3091),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3149),
.Y(n_3374)
);

CKINVDCx5p33_ASAP7_75t_R g3375 ( 
.A(n_3204),
.Y(n_3375)
);

OAI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_3299),
.A2(n_3051),
.B(n_3087),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_3181),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_SL g3378 ( 
.A(n_3152),
.B(n_3112),
.Y(n_3378)
);

BUFx2_ASAP7_75t_SL g3379 ( 
.A(n_3228),
.Y(n_3379)
);

INVx5_ASAP7_75t_L g3380 ( 
.A(n_3193),
.Y(n_3380)
);

BUFx12f_ASAP7_75t_L g3381 ( 
.A(n_3160),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3236),
.B(n_55),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3294),
.B(n_58),
.Y(n_3383)
);

INVx4_ASAP7_75t_L g3384 ( 
.A(n_3304),
.Y(n_3384)
);

BUFx6f_ASAP7_75t_L g3385 ( 
.A(n_3179),
.Y(n_3385)
);

AO32x1_ASAP7_75t_L g3386 ( 
.A1(n_3282),
.A2(n_3107),
.A3(n_3100),
.B1(n_3092),
.B2(n_63),
.Y(n_3386)
);

CKINVDCx5p33_ASAP7_75t_R g3387 ( 
.A(n_3240),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3182),
.Y(n_3388)
);

HB1xp67_ASAP7_75t_L g3389 ( 
.A(n_3185),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_3323),
.A2(n_3118),
.B(n_3095),
.Y(n_3390)
);

INVx4_ASAP7_75t_SL g3391 ( 
.A(n_3274),
.Y(n_3391)
);

OAI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_3318),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_3392)
);

OR2x6_ASAP7_75t_L g3393 ( 
.A(n_3307),
.B(n_1458),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_SL g3394 ( 
.A(n_3304),
.B(n_1458),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3156),
.Y(n_3395)
);

AOI21xp5_ASAP7_75t_L g3396 ( 
.A1(n_3317),
.A2(n_3227),
.B(n_3232),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3301),
.B(n_59),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3210),
.B(n_3338),
.Y(n_3398)
);

INVx2_ASAP7_75t_SL g3399 ( 
.A(n_3211),
.Y(n_3399)
);

OAI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3314),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3156),
.Y(n_3401)
);

OAI21x1_ASAP7_75t_SL g3402 ( 
.A1(n_3265),
.A2(n_65),
.B(n_66),
.Y(n_3402)
);

INVx2_ASAP7_75t_SL g3403 ( 
.A(n_3213),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3163),
.B(n_66),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_SL g3405 ( 
.A1(n_3222),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_3405)
);

INVxp67_ASAP7_75t_L g3406 ( 
.A(n_3336),
.Y(n_3406)
);

HB1xp67_ASAP7_75t_L g3407 ( 
.A(n_3184),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3191),
.Y(n_3408)
);

BUFx12f_ASAP7_75t_L g3409 ( 
.A(n_3160),
.Y(n_3409)
);

INVx3_ASAP7_75t_L g3410 ( 
.A(n_3261),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_3304),
.Y(n_3411)
);

AND2x4_ASAP7_75t_L g3412 ( 
.A(n_3208),
.B(n_68),
.Y(n_3412)
);

BUFx4_ASAP7_75t_SL g3413 ( 
.A(n_3275),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_3213),
.Y(n_3414)
);

CKINVDCx11_ASAP7_75t_R g3415 ( 
.A(n_3176),
.Y(n_3415)
);

OAI22xp33_ASAP7_75t_SL g3416 ( 
.A1(n_3199),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3338),
.B(n_72),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3224),
.B(n_73),
.Y(n_3418)
);

INVx4_ASAP7_75t_L g3419 ( 
.A(n_3213),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3241),
.A2(n_3278),
.B(n_3327),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3192),
.A2(n_1465),
.B(n_1458),
.Y(n_3421)
);

AND2x4_ASAP7_75t_L g3422 ( 
.A(n_3157),
.B(n_73),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3191),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3157),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3348),
.A2(n_3186),
.B1(n_3201),
.B2(n_3250),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3161),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3153),
.B(n_75),
.Y(n_3427)
);

AND2x4_ASAP7_75t_L g3428 ( 
.A(n_3161),
.B(n_75),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3246),
.B(n_3253),
.Y(n_3429)
);

BUFx2_ASAP7_75t_SL g3430 ( 
.A(n_3237),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3167),
.Y(n_3431)
);

BUFx3_ASAP7_75t_L g3432 ( 
.A(n_3174),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_3243),
.Y(n_3433)
);

AOI22xp33_ASAP7_75t_L g3434 ( 
.A1(n_3276),
.A2(n_79),
.B1(n_76),
.B2(n_77),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3303),
.B(n_77),
.Y(n_3435)
);

INVx1_ASAP7_75t_SL g3436 ( 
.A(n_3169),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3319),
.B(n_79),
.Y(n_3437)
);

CKINVDCx5p33_ASAP7_75t_R g3438 ( 
.A(n_3243),
.Y(n_3438)
);

OR2x6_ASAP7_75t_L g3439 ( 
.A(n_3307),
.B(n_1465),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3167),
.Y(n_3440)
);

AND2x4_ASAP7_75t_L g3441 ( 
.A(n_3168),
.B(n_3171),
.Y(n_3441)
);

INVx1_ASAP7_75t_SL g3442 ( 
.A(n_3172),
.Y(n_3442)
);

OAI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_3231),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3216),
.B(n_80),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3283),
.B(n_82),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3168),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3192),
.A2(n_1468),
.B(n_1465),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3267),
.A2(n_87),
.B1(n_84),
.B2(n_85),
.Y(n_3448)
);

BUFx2_ASAP7_75t_L g3449 ( 
.A(n_3256),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3171),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_3245),
.A2(n_88),
.B1(n_84),
.B2(n_85),
.Y(n_3451)
);

INVx2_ASAP7_75t_SL g3452 ( 
.A(n_3221),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3148),
.Y(n_3453)
);

INVx1_ASAP7_75t_SL g3454 ( 
.A(n_3235),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_3221),
.Y(n_3455)
);

INVx2_ASAP7_75t_SL g3456 ( 
.A(n_3221),
.Y(n_3456)
);

NAND2x1p5_ASAP7_75t_L g3457 ( 
.A(n_3217),
.B(n_1468),
.Y(n_3457)
);

OAI22xp5_ASAP7_75t_L g3458 ( 
.A1(n_3330),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3207),
.Y(n_3459)
);

AND2x6_ASAP7_75t_L g3460 ( 
.A(n_3170),
.B(n_91),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3349),
.B(n_91),
.Y(n_3461)
);

BUFx2_ASAP7_75t_L g3462 ( 
.A(n_3258),
.Y(n_3462)
);

AOI21xp33_ASAP7_75t_L g3463 ( 
.A1(n_3339),
.A2(n_92),
.B(n_94),
.Y(n_3463)
);

OAI22xp5_ASAP7_75t_L g3464 ( 
.A1(n_3341),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_3464)
);

INVx2_ASAP7_75t_SL g3465 ( 
.A(n_3225),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3190),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3316),
.B(n_96),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3198),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3349),
.B(n_97),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3251),
.B(n_97),
.Y(n_3470)
);

BUFx6f_ASAP7_75t_L g3471 ( 
.A(n_3148),
.Y(n_3471)
);

AND2x4_ASAP7_75t_L g3472 ( 
.A(n_3259),
.B(n_98),
.Y(n_3472)
);

BUFx6f_ASAP7_75t_L g3473 ( 
.A(n_3148),
.Y(n_3473)
);

OR2x6_ASAP7_75t_L g3474 ( 
.A(n_3199),
.B(n_3351),
.Y(n_3474)
);

BUFx6f_ASAP7_75t_L g3475 ( 
.A(n_3155),
.Y(n_3475)
);

BUFx2_ASAP7_75t_L g3476 ( 
.A(n_3164),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3259),
.B(n_98),
.Y(n_3477)
);

O2A1O1Ixp33_ASAP7_75t_L g3478 ( 
.A1(n_3354),
.A2(n_99),
.B(n_100),
.C(n_101),
.Y(n_3478)
);

OAI21x1_ASAP7_75t_L g3479 ( 
.A1(n_3312),
.A2(n_265),
.B(n_263),
.Y(n_3479)
);

OAI21x1_ASAP7_75t_L g3480 ( 
.A1(n_3302),
.A2(n_267),
.B(n_266),
.Y(n_3480)
);

INVx3_ASAP7_75t_L g3481 ( 
.A(n_3247),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3220),
.Y(n_3482)
);

OAI21x1_ASAP7_75t_L g3483 ( 
.A1(n_3302),
.A2(n_277),
.B(n_274),
.Y(n_3483)
);

AND2x2_ASAP7_75t_L g3484 ( 
.A(n_3315),
.B(n_100),
.Y(n_3484)
);

O2A1O1Ixp5_ASAP7_75t_L g3485 ( 
.A1(n_3339),
.A2(n_105),
.B(n_108),
.C(n_109),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3345),
.B(n_1468),
.Y(n_3486)
);

BUFx6f_ASAP7_75t_L g3487 ( 
.A(n_3155),
.Y(n_3487)
);

OR2x6_ASAP7_75t_L g3488 ( 
.A(n_3351),
.B(n_1468),
.Y(n_3488)
);

AND2x4_ASAP7_75t_L g3489 ( 
.A(n_3215),
.B(n_105),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3315),
.B(n_3345),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3295),
.B(n_109),
.Y(n_3491)
);

CKINVDCx16_ASAP7_75t_R g3492 ( 
.A(n_3298),
.Y(n_3492)
);

AND2x4_ASAP7_75t_L g3493 ( 
.A(n_3270),
.B(n_110),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3295),
.B(n_111),
.Y(n_3494)
);

BUFx6f_ASAP7_75t_L g3495 ( 
.A(n_3155),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3220),
.Y(n_3496)
);

BUFx2_ASAP7_75t_L g3497 ( 
.A(n_3164),
.Y(n_3497)
);

BUFx12f_ASAP7_75t_L g3498 ( 
.A(n_3345),
.Y(n_3498)
);

AND2x4_ASAP7_75t_L g3499 ( 
.A(n_3217),
.B(n_111),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_3217),
.B(n_1468),
.Y(n_3500)
);

OR2x6_ASAP7_75t_L g3501 ( 
.A(n_3170),
.B(n_278),
.Y(n_3501)
);

BUFx2_ASAP7_75t_L g3502 ( 
.A(n_3209),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3332),
.A2(n_1467),
.B(n_1457),
.Y(n_3503)
);

NOR2xp67_ASAP7_75t_L g3504 ( 
.A(n_3189),
.B(n_114),
.Y(n_3504)
);

CKINVDCx5p33_ASAP7_75t_R g3505 ( 
.A(n_3279),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3320),
.B(n_116),
.Y(n_3506)
);

CKINVDCx20_ASAP7_75t_R g3507 ( 
.A(n_3188),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3254),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3159),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_3509)
);

BUFx3_ASAP7_75t_L g3510 ( 
.A(n_3225),
.Y(n_3510)
);

INVx4_ASAP7_75t_L g3511 ( 
.A(n_3189),
.Y(n_3511)
);

O2A1O1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3300),
.A2(n_119),
.B(n_124),
.C(n_125),
.Y(n_3512)
);

AND2x4_ASAP7_75t_L g3513 ( 
.A(n_3290),
.B(n_124),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3257),
.Y(n_3514)
);

INVx2_ASAP7_75t_SL g3515 ( 
.A(n_3225),
.Y(n_3515)
);

AOI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_3350),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3324),
.A2(n_1467),
.B(n_1457),
.Y(n_3517)
);

INVx3_ASAP7_75t_L g3518 ( 
.A(n_3209),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3252),
.B(n_131),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3329),
.B(n_131),
.Y(n_3520)
);

INVx2_ASAP7_75t_SL g3521 ( 
.A(n_3151),
.Y(n_3521)
);

AOI21xp5_ASAP7_75t_L g3522 ( 
.A1(n_3310),
.A2(n_1467),
.B(n_1457),
.Y(n_3522)
);

AND2x4_ASAP7_75t_L g3523 ( 
.A(n_3290),
.B(n_132),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3281),
.Y(n_3524)
);

BUFx2_ASAP7_75t_L g3525 ( 
.A(n_3212),
.Y(n_3525)
);

CKINVDCx11_ASAP7_75t_R g3526 ( 
.A(n_3233),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3273),
.B(n_3335),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3281),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3277),
.B(n_3226),
.Y(n_3529)
);

INVx3_ASAP7_75t_L g3530 ( 
.A(n_3212),
.Y(n_3530)
);

INVx5_ASAP7_75t_L g3531 ( 
.A(n_3358),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3173),
.B(n_132),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_3385),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3527),
.B(n_3268),
.Y(n_3534)
);

CKINVDCx20_ASAP7_75t_R g3535 ( 
.A(n_3368),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3424),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3425),
.A2(n_3195),
.B1(n_3238),
.B2(n_3333),
.Y(n_3537)
);

BUFx2_ASAP7_75t_L g3538 ( 
.A(n_3498),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3424),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3369),
.B(n_3331),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3426),
.Y(n_3541)
);

AOI22xp33_ASAP7_75t_SL g3542 ( 
.A1(n_3460),
.A2(n_3353),
.B1(n_3290),
.B2(n_3311),
.Y(n_3542)
);

INVx6_ASAP7_75t_L g3543 ( 
.A(n_3385),
.Y(n_3543)
);

AOI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3366),
.A2(n_3361),
.B(n_3310),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_L g3545 ( 
.A1(n_3400),
.A2(n_3343),
.B1(n_3264),
.B2(n_3234),
.Y(n_3545)
);

BUFx3_ASAP7_75t_L g3546 ( 
.A(n_3385),
.Y(n_3546)
);

CKINVDCx14_ASAP7_75t_R g3547 ( 
.A(n_3387),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3441),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3441),
.Y(n_3549)
);

INVx6_ASAP7_75t_L g3550 ( 
.A(n_3381),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3481),
.Y(n_3551)
);

INVxp67_ASAP7_75t_SL g3552 ( 
.A(n_3407),
.Y(n_3552)
);

BUFx6f_ASAP7_75t_SL g3553 ( 
.A(n_3499),
.Y(n_3553)
);

AOI22xp5_ASAP7_75t_L g3554 ( 
.A1(n_3448),
.A2(n_3200),
.B1(n_3264),
.B2(n_3196),
.Y(n_3554)
);

BUFx10_ASAP7_75t_L g3555 ( 
.A(n_3433),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3426),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_SL g3557 ( 
.A1(n_3460),
.A2(n_3196),
.B1(n_3334),
.B2(n_3280),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3408),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_SL g3559 ( 
.A1(n_3460),
.A2(n_3280),
.B1(n_3292),
.B2(n_3313),
.Y(n_3559)
);

INVx5_ASAP7_75t_L g3560 ( 
.A(n_3409),
.Y(n_3560)
);

OAI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_3501),
.A2(n_3308),
.B1(n_3337),
.B2(n_3178),
.Y(n_3561)
);

AND2x4_ASAP7_75t_L g3562 ( 
.A(n_3384),
.B(n_3269),
.Y(n_3562)
);

INVx6_ASAP7_75t_L g3563 ( 
.A(n_3391),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3408),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_SL g3565 ( 
.A1(n_3460),
.A2(n_3292),
.B1(n_3313),
.B2(n_3305),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3389),
.B(n_3344),
.Y(n_3566)
);

BUFx12f_ASAP7_75t_L g3567 ( 
.A(n_3438),
.Y(n_3567)
);

INVx5_ASAP7_75t_L g3568 ( 
.A(n_3511),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3423),
.Y(n_3569)
);

AOI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3463),
.A2(n_3352),
.B1(n_3309),
.B2(n_3305),
.Y(n_3570)
);

BUFx2_ASAP7_75t_L g3571 ( 
.A(n_3384),
.Y(n_3571)
);

BUFx8_ASAP7_75t_SL g3572 ( 
.A(n_3505),
.Y(n_3572)
);

BUFx3_ASAP7_75t_L g3573 ( 
.A(n_3415),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3392),
.A2(n_3288),
.B1(n_3357),
.B2(n_3150),
.Y(n_3574)
);

BUFx4f_ASAP7_75t_L g3575 ( 
.A(n_3499),
.Y(n_3575)
);

INVx6_ASAP7_75t_L g3576 ( 
.A(n_3391),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3423),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_L g3578 ( 
.A1(n_3376),
.A2(n_3288),
.B1(n_3150),
.B2(n_3287),
.Y(n_3578)
);

CKINVDCx11_ASAP7_75t_R g3579 ( 
.A(n_3507),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3370),
.Y(n_3580)
);

CKINVDCx11_ASAP7_75t_R g3581 ( 
.A(n_3526),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_L g3582 ( 
.A1(n_3443),
.A2(n_3358),
.B1(n_3359),
.B2(n_3355),
.Y(n_3582)
);

AOI22xp33_ASAP7_75t_SL g3583 ( 
.A1(n_3416),
.A2(n_3313),
.B1(n_3205),
.B2(n_3358),
.Y(n_3583)
);

OAI21xp5_ASAP7_75t_SL g3584 ( 
.A1(n_3516),
.A2(n_3203),
.B(n_3325),
.Y(n_3584)
);

AOI22xp5_ASAP7_75t_L g3585 ( 
.A1(n_3451),
.A2(n_3347),
.B1(n_3206),
.B2(n_3205),
.Y(n_3585)
);

HB1xp67_ASAP7_75t_L g3586 ( 
.A(n_3364),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3374),
.Y(n_3587)
);

AOI22xp33_ASAP7_75t_SL g3588 ( 
.A1(n_3378),
.A2(n_3328),
.B1(n_3359),
.B2(n_3260),
.Y(n_3588)
);

CKINVDCx6p67_ASAP7_75t_R g3589 ( 
.A(n_3379),
.Y(n_3589)
);

BUFx6f_ASAP7_75t_L g3590 ( 
.A(n_3453),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_SL g3591 ( 
.A(n_3513),
.Y(n_3591)
);

INVx2_ASAP7_75t_SL g3592 ( 
.A(n_3429),
.Y(n_3592)
);

BUFx3_ASAP7_75t_L g3593 ( 
.A(n_3375),
.Y(n_3593)
);

OAI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3501),
.A2(n_3188),
.B1(n_3197),
.B2(n_3342),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_SL g3595 ( 
.A1(n_3500),
.A2(n_3202),
.B(n_3260),
.Y(n_3595)
);

BUFx2_ASAP7_75t_L g3596 ( 
.A(n_3411),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3398),
.B(n_3344),
.Y(n_3597)
);

AOI22xp33_ASAP7_75t_SL g3598 ( 
.A1(n_3513),
.A2(n_3359),
.B1(n_3189),
.B2(n_3360),
.Y(n_3598)
);

OAI22xp5_ASAP7_75t_SL g3599 ( 
.A1(n_3492),
.A2(n_3187),
.B1(n_3194),
.B2(n_3239),
.Y(n_3599)
);

INVx6_ASAP7_75t_L g3600 ( 
.A(n_3419),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3481),
.Y(n_3601)
);

CKINVDCx20_ASAP7_75t_R g3602 ( 
.A(n_3436),
.Y(n_3602)
);

BUFx2_ASAP7_75t_SL g3603 ( 
.A(n_3454),
.Y(n_3603)
);

INVx4_ASAP7_75t_L g3604 ( 
.A(n_3523),
.Y(n_3604)
);

AOI22xp5_ASAP7_75t_L g3605 ( 
.A1(n_3434),
.A2(n_3183),
.B1(n_3242),
.B2(n_3297),
.Y(n_3605)
);

AOI22xp5_ASAP7_75t_L g3606 ( 
.A1(n_3509),
.A2(n_3464),
.B1(n_3458),
.B2(n_3519),
.Y(n_3606)
);

INVx8_ASAP7_75t_L g3607 ( 
.A(n_3523),
.Y(n_3607)
);

BUFx2_ASAP7_75t_L g3608 ( 
.A(n_3411),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3363),
.B(n_3293),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3395),
.Y(n_3610)
);

BUFx3_ASAP7_75t_L g3611 ( 
.A(n_3462),
.Y(n_3611)
);

NAND2x1p5_ASAP7_75t_L g3612 ( 
.A(n_3531),
.B(n_3197),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3478),
.A2(n_3284),
.B1(n_3291),
.B2(n_3296),
.Y(n_3613)
);

INVx2_ASAP7_75t_SL g3614 ( 
.A(n_3490),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3450),
.Y(n_3615)
);

OAI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3474),
.A2(n_3285),
.B1(n_3255),
.B2(n_3233),
.Y(n_3616)
);

OAI22xp5_ASAP7_75t_L g3617 ( 
.A1(n_3512),
.A2(n_3474),
.B1(n_3371),
.B2(n_3380),
.Y(n_3617)
);

CKINVDCx6p67_ASAP7_75t_R g3618 ( 
.A(n_3430),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3401),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3396),
.A2(n_3326),
.B1(n_3277),
.B2(n_3289),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3472),
.A2(n_3277),
.B1(n_3346),
.B2(n_3322),
.Y(n_3621)
);

OAI22xp5_ASAP7_75t_L g3622 ( 
.A1(n_3371),
.A2(n_3244),
.B1(n_3272),
.B2(n_3340),
.Y(n_3622)
);

BUFx2_ASAP7_75t_SL g3623 ( 
.A(n_3403),
.Y(n_3623)
);

OAI22xp5_ASAP7_75t_L g3624 ( 
.A1(n_3371),
.A2(n_3306),
.B1(n_3233),
.B2(n_3255),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3431),
.Y(n_3625)
);

INVx4_ASAP7_75t_L g3626 ( 
.A(n_3453),
.Y(n_3626)
);

CKINVDCx11_ASAP7_75t_R g3627 ( 
.A(n_3442),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3440),
.Y(n_3628)
);

OAI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3383),
.A2(n_3180),
.B1(n_3223),
.B2(n_3346),
.Y(n_3629)
);

CKINVDCx20_ASAP7_75t_R g3630 ( 
.A(n_3406),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3446),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3367),
.Y(n_3632)
);

CKINVDCx11_ASAP7_75t_R g3633 ( 
.A(n_3453),
.Y(n_3633)
);

BUFx8_ASAP7_75t_L g3634 ( 
.A(n_3444),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3482),
.Y(n_3635)
);

AOI22xp33_ASAP7_75t_L g3636 ( 
.A1(n_3472),
.A2(n_3322),
.B1(n_3321),
.B2(n_3271),
.Y(n_3636)
);

AOI22xp5_ASAP7_75t_L g3637 ( 
.A1(n_3493),
.A2(n_3218),
.B1(n_3266),
.B2(n_3321),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3496),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3524),
.Y(n_3639)
);

BUFx10_ASAP7_75t_L g3640 ( 
.A(n_3493),
.Y(n_3640)
);

BUFx2_ASAP7_75t_L g3641 ( 
.A(n_3476),
.Y(n_3641)
);

OAI22xp5_ASAP7_75t_L g3642 ( 
.A1(n_3461),
.A2(n_3306),
.B1(n_3154),
.B2(n_3255),
.Y(n_3642)
);

BUFx8_ASAP7_75t_SL g3643 ( 
.A(n_3471),
.Y(n_3643)
);

BUFx2_ASAP7_75t_L g3644 ( 
.A(n_3497),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3377),
.Y(n_3645)
);

BUFx10_ASAP7_75t_L g3646 ( 
.A(n_3422),
.Y(n_3646)
);

BUFx2_ASAP7_75t_L g3647 ( 
.A(n_3449),
.Y(n_3647)
);

BUFx3_ASAP7_75t_L g3648 ( 
.A(n_3414),
.Y(n_3648)
);

INVx2_ASAP7_75t_SL g3649 ( 
.A(n_3414),
.Y(n_3649)
);

AOI22xp33_ASAP7_75t_SL g3650 ( 
.A1(n_3402),
.A2(n_3263),
.B1(n_3271),
.B2(n_3177),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3373),
.A2(n_3271),
.B1(n_3263),
.B2(n_3151),
.Y(n_3651)
);

BUFx3_ASAP7_75t_L g3652 ( 
.A(n_3432),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3399),
.Y(n_3653)
);

CKINVDCx11_ASAP7_75t_R g3654 ( 
.A(n_3471),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3529),
.Y(n_3655)
);

CKINVDCx6p67_ASAP7_75t_R g3656 ( 
.A(n_3510),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3524),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3528),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3388),
.Y(n_3659)
);

AOI22xp33_ASAP7_75t_SL g3660 ( 
.A1(n_3531),
.A2(n_3263),
.B1(n_3158),
.B2(n_3177),
.Y(n_3660)
);

BUFx2_ASAP7_75t_L g3661 ( 
.A(n_3502),
.Y(n_3661)
);

OAI22xp33_ASAP7_75t_L g3662 ( 
.A1(n_3380),
.A2(n_3158),
.B1(n_3249),
.B2(n_3286),
.Y(n_3662)
);

HB1xp67_ASAP7_75t_L g3663 ( 
.A(n_3528),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3459),
.Y(n_3664)
);

BUFx12f_ASAP7_75t_L g3665 ( 
.A(n_3427),
.Y(n_3665)
);

AOI22xp33_ASAP7_75t_L g3666 ( 
.A1(n_3365),
.A2(n_3249),
.B1(n_3286),
.B2(n_3219),
.Y(n_3666)
);

NAND2xp33_ASAP7_75t_SL g3667 ( 
.A(n_3422),
.B(n_3248),
.Y(n_3667)
);

INVx6_ASAP7_75t_L g3668 ( 
.A(n_3419),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3663),
.Y(n_3669)
);

BUFx2_ASAP7_75t_SL g3670 ( 
.A(n_3560),
.Y(n_3670)
);

AOI22xp33_ASAP7_75t_L g3671 ( 
.A1(n_3544),
.A2(n_3372),
.B1(n_3380),
.B2(n_3504),
.Y(n_3671)
);

CKINVDCx11_ASAP7_75t_R g3672 ( 
.A(n_3555),
.Y(n_3672)
);

OA21x2_ASAP7_75t_L g3673 ( 
.A1(n_3635),
.A2(n_3447),
.B(n_3421),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3638),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3536),
.Y(n_3675)
);

AO21x2_ASAP7_75t_L g3676 ( 
.A1(n_3662),
.A2(n_3522),
.B(n_3420),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3539),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3541),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3556),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3558),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3564),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3569),
.Y(n_3682)
);

OAI22xp5_ASAP7_75t_L g3683 ( 
.A1(n_3537),
.A2(n_3531),
.B1(n_3394),
.B2(n_3428),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3661),
.B(n_3525),
.Y(n_3684)
);

INVx1_ASAP7_75t_SL g3685 ( 
.A(n_3627),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3577),
.Y(n_3686)
);

INVx4_ASAP7_75t_L g3687 ( 
.A(n_3560),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3639),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3657),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3658),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3580),
.Y(n_3691)
);

AOI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3571),
.A2(n_3469),
.B(n_3397),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3587),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3610),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3615),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3664),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3619),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3584),
.A2(n_3485),
.B(n_3532),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3628),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3625),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3641),
.B(n_3518),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3597),
.A2(n_3530),
.B(n_3518),
.Y(n_3702)
);

OAI21x1_ASAP7_75t_L g3703 ( 
.A1(n_3566),
.A2(n_3530),
.B(n_3410),
.Y(n_3703)
);

OAI21xp5_ASAP7_75t_L g3704 ( 
.A1(n_3584),
.A2(n_3417),
.B(n_3520),
.Y(n_3704)
);

OAI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3666),
.A2(n_3410),
.B(n_3362),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3631),
.Y(n_3706)
);

HB1xp67_ASAP7_75t_L g3707 ( 
.A(n_3586),
.Y(n_3707)
);

BUFx2_ASAP7_75t_L g3708 ( 
.A(n_3596),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3632),
.Y(n_3709)
);

OAI21x1_ASAP7_75t_L g3710 ( 
.A1(n_3624),
.A2(n_3362),
.B(n_3248),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3645),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3659),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3540),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3644),
.B(n_3508),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3552),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3647),
.B(n_3548),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3549),
.Y(n_3717)
);

HB1xp67_ASAP7_75t_L g3718 ( 
.A(n_3608),
.Y(n_3718)
);

OAI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3636),
.A2(n_3390),
.B(n_3514),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3551),
.Y(n_3720)
);

OAI22xp33_ASAP7_75t_L g3721 ( 
.A1(n_3554),
.A2(n_3488),
.B1(n_3511),
.B2(n_3439),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3601),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3534),
.Y(n_3723)
);

AND2x4_ASAP7_75t_L g3724 ( 
.A(n_3568),
.B(n_3372),
.Y(n_3724)
);

INVx3_ASAP7_75t_L g3725 ( 
.A(n_3568),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3568),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3609),
.B(n_3521),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3649),
.B(n_3468),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3611),
.B(n_3466),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3646),
.Y(n_3730)
);

OAI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3554),
.A2(n_3542),
.B1(n_3545),
.B2(n_3559),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3646),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3640),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3562),
.Y(n_3734)
);

INVx1_ASAP7_75t_SL g3735 ( 
.A(n_3579),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3629),
.B(n_3470),
.Y(n_3736)
);

INVx8_ASAP7_75t_L g3737 ( 
.A(n_3533),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3562),
.Y(n_3738)
);

INVx3_ASAP7_75t_L g3739 ( 
.A(n_3589),
.Y(n_3739)
);

AOI22xp33_ASAP7_75t_L g3740 ( 
.A1(n_3599),
.A2(n_3477),
.B1(n_3412),
.B2(n_3428),
.Y(n_3740)
);

INVx2_ASAP7_75t_SL g3741 ( 
.A(n_3600),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3640),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3667),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3629),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3623),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3603),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3642),
.Y(n_3747)
);

INVxp67_ASAP7_75t_L g3748 ( 
.A(n_3599),
.Y(n_3748)
);

OA21x2_ASAP7_75t_L g3749 ( 
.A1(n_3621),
.A2(n_3494),
.B(n_3491),
.Y(n_3749)
);

AO31x2_ASAP7_75t_L g3750 ( 
.A1(n_3617),
.A2(n_3503),
.A3(n_3418),
.B(n_3437),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3626),
.Y(n_3751)
);

INVx1_ASAP7_75t_SL g3752 ( 
.A(n_3581),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3618),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3642),
.A2(n_3457),
.B(n_3486),
.Y(n_3754)
);

INVx3_ASAP7_75t_L g3755 ( 
.A(n_3600),
.Y(n_3755)
);

AOI21x1_ASAP7_75t_L g3756 ( 
.A1(n_3538),
.A2(n_3445),
.B(n_3506),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3648),
.Y(n_3757)
);

BUFx2_ASAP7_75t_L g3758 ( 
.A(n_3604),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_3655),
.B(n_3452),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3626),
.Y(n_3760)
);

INVx4_ASAP7_75t_L g3761 ( 
.A(n_3560),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_3614),
.B(n_3455),
.Y(n_3762)
);

BUFx8_ASAP7_75t_L g3763 ( 
.A(n_3533),
.Y(n_3763)
);

AO21x2_ASAP7_75t_L g3764 ( 
.A1(n_3616),
.A2(n_3405),
.B(n_3412),
.Y(n_3764)
);

HB1xp67_ASAP7_75t_L g3765 ( 
.A(n_3653),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3592),
.B(n_3652),
.Y(n_3766)
);

HB1xp67_ASAP7_75t_L g3767 ( 
.A(n_3590),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3668),
.Y(n_3768)
);

BUFx6f_ASAP7_75t_L g3769 ( 
.A(n_3533),
.Y(n_3769)
);

INVx3_ASAP7_75t_L g3770 ( 
.A(n_3668),
.Y(n_3770)
);

OAI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3622),
.A2(n_3483),
.B(n_3480),
.Y(n_3771)
);

NAND2x1p5_ASAP7_75t_L g3772 ( 
.A(n_3575),
.B(n_3471),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3604),
.B(n_3456),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3590),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3656),
.B(n_3465),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3590),
.Y(n_3776)
);

BUFx3_ASAP7_75t_L g3777 ( 
.A(n_3573),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3651),
.B(n_3382),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3553),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3612),
.A2(n_3594),
.B(n_3582),
.Y(n_3780)
);

BUFx3_ASAP7_75t_L g3781 ( 
.A(n_3563),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3553),
.Y(n_3782)
);

HB1xp67_ASAP7_75t_L g3783 ( 
.A(n_3602),
.Y(n_3783)
);

BUFx3_ASAP7_75t_L g3784 ( 
.A(n_3563),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3598),
.B(n_3467),
.Y(n_3785)
);

BUFx2_ASAP7_75t_R g3786 ( 
.A(n_3572),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3591),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3591),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3607),
.Y(n_3789)
);

BUFx3_ASAP7_75t_L g3790 ( 
.A(n_3576),
.Y(n_3790)
);

AOI21x1_ASAP7_75t_L g3791 ( 
.A1(n_3613),
.A2(n_3484),
.B(n_3489),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3607),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3650),
.B(n_3404),
.Y(n_3793)
);

AND2x2_ASAP7_75t_L g3794 ( 
.A(n_3660),
.B(n_3515),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_3675),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3675),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3677),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3677),
.Y(n_3798)
);

BUFx2_ASAP7_75t_L g3799 ( 
.A(n_3687),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3758),
.B(n_3546),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3691),
.Y(n_3801)
);

OAI21x1_ASAP7_75t_L g3802 ( 
.A1(n_3705),
.A2(n_3620),
.B(n_3595),
.Y(n_3802)
);

HB1xp67_ASAP7_75t_L g3803 ( 
.A(n_3707),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3679),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3694),
.Y(n_3805)
);

OA21x2_ASAP7_75t_L g3806 ( 
.A1(n_3710),
.A2(n_3570),
.B(n_3606),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3695),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3678),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3679),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3680),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3758),
.B(n_3557),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3681),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3708),
.B(n_3576),
.Y(n_3813)
);

INVxp67_ASAP7_75t_L g3814 ( 
.A(n_3670),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3682),
.Y(n_3815)
);

BUFx2_ASAP7_75t_L g3816 ( 
.A(n_3687),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3686),
.Y(n_3817)
);

INVx2_ASAP7_75t_SL g3818 ( 
.A(n_3737),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3688),
.Y(n_3819)
);

OR2x2_ASAP7_75t_L g3820 ( 
.A(n_3744),
.B(n_3607),
.Y(n_3820)
);

BUFx6f_ASAP7_75t_L g3821 ( 
.A(n_3672),
.Y(n_3821)
);

AND2x2_ASAP7_75t_L g3822 ( 
.A(n_3708),
.B(n_3575),
.Y(n_3822)
);

OR2x2_ASAP7_75t_L g3823 ( 
.A(n_3713),
.B(n_3613),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3689),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3681),
.Y(n_3825)
);

AOI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3726),
.A2(n_3435),
.B(n_3561),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3674),
.Y(n_3827)
);

HB1xp67_ASAP7_75t_L g3828 ( 
.A(n_3718),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3747),
.B(n_3583),
.Y(n_3829)
);

AND2x4_ASAP7_75t_L g3830 ( 
.A(n_3725),
.B(n_3593),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3755),
.B(n_3543),
.Y(n_3831)
);

INVx3_ASAP7_75t_L g3832 ( 
.A(n_3687),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3674),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3693),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3693),
.Y(n_3835)
);

HB1xp67_ASAP7_75t_L g3836 ( 
.A(n_3669),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3749),
.B(n_3489),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3720),
.Y(n_3838)
);

OR2x2_ASAP7_75t_L g3839 ( 
.A(n_3713),
.B(n_3637),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3720),
.Y(n_3840)
);

HB1xp67_ASAP7_75t_L g3841 ( 
.A(n_3699),
.Y(n_3841)
);

INVx1_ASAP7_75t_SL g3842 ( 
.A(n_3672),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3690),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3722),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3696),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3706),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3722),
.Y(n_3847)
);

HB1xp67_ASAP7_75t_L g3848 ( 
.A(n_3715),
.Y(n_3848)
);

INVx2_ASAP7_75t_SL g3849 ( 
.A(n_3737),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3697),
.Y(n_3850)
);

OAI21x1_ASAP7_75t_L g3851 ( 
.A1(n_3705),
.A2(n_3578),
.B(n_3479),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3755),
.B(n_3543),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3709),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3709),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3749),
.B(n_3637),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3749),
.B(n_3588),
.Y(n_3856)
);

BUFx6f_ASAP7_75t_L g3857 ( 
.A(n_3769),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3711),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3711),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3697),
.Y(n_3860)
);

CKINVDCx20_ASAP7_75t_R g3861 ( 
.A(n_3783),
.Y(n_3861)
);

OAI21x1_ASAP7_75t_L g3862 ( 
.A1(n_3710),
.A2(n_3574),
.B(n_3585),
.Y(n_3862)
);

OA21x2_ASAP7_75t_L g3863 ( 
.A1(n_3702),
.A2(n_3703),
.B(n_3780),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3712),
.Y(n_3864)
);

OR2x2_ASAP7_75t_L g3865 ( 
.A(n_3723),
.B(n_3488),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3712),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3755),
.B(n_3633),
.Y(n_3867)
);

CKINVDCx14_ASAP7_75t_R g3868 ( 
.A(n_3739),
.Y(n_3868)
);

AO21x2_ASAP7_75t_L g3869 ( 
.A1(n_3726),
.A2(n_3606),
.B(n_3605),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3700),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3770),
.B(n_3654),
.Y(n_3871)
);

BUFx2_ASAP7_75t_L g3872 ( 
.A(n_3761),
.Y(n_3872)
);

AND2x2_ASAP7_75t_L g3873 ( 
.A(n_3770),
.B(n_3550),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3770),
.B(n_3550),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3700),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3728),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3728),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3767),
.Y(n_3878)
);

BUFx2_ASAP7_75t_SL g3879 ( 
.A(n_3739),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3791),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3717),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3791),
.Y(n_3882)
);

BUFx4f_ASAP7_75t_SL g3883 ( 
.A(n_3752),
.Y(n_3883)
);

OR2x6_ASAP7_75t_L g3884 ( 
.A(n_3670),
.B(n_3761),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3774),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3733),
.B(n_3555),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3733),
.B(n_3630),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3774),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3776),
.Y(n_3889)
);

AO21x2_ASAP7_75t_L g3890 ( 
.A1(n_3698),
.A2(n_3676),
.B(n_3721),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3776),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3751),
.Y(n_3892)
);

OR2x2_ASAP7_75t_L g3893 ( 
.A(n_3750),
.B(n_3473),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3742),
.B(n_3565),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3751),
.Y(n_3895)
);

HB1xp67_ASAP7_75t_L g3896 ( 
.A(n_3692),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3702),
.Y(n_3897)
);

INVx3_ASAP7_75t_L g3898 ( 
.A(n_3761),
.Y(n_3898)
);

OR2x2_ASAP7_75t_L g3899 ( 
.A(n_3750),
.B(n_3473),
.Y(n_3899)
);

AND2x4_ASAP7_75t_L g3900 ( 
.A(n_3725),
.B(n_3473),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3760),
.Y(n_3901)
);

OR2x2_ASAP7_75t_L g3902 ( 
.A(n_3750),
.B(n_3475),
.Y(n_3902)
);

OR2x6_ASAP7_75t_L g3903 ( 
.A(n_3725),
.B(n_3393),
.Y(n_3903)
);

OAI21x1_ASAP7_75t_L g3904 ( 
.A1(n_3703),
.A2(n_3719),
.B(n_3780),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3742),
.B(n_3547),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3760),
.Y(n_3906)
);

AND2x2_ASAP7_75t_L g3907 ( 
.A(n_3724),
.B(n_3794),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3692),
.Y(n_3908)
);

OAI21x1_ASAP7_75t_L g3909 ( 
.A1(n_3719),
.A2(n_3585),
.B(n_3356),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3729),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3714),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3724),
.B(n_3665),
.Y(n_3912)
);

HB1xp67_ASAP7_75t_L g3913 ( 
.A(n_3764),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3729),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3734),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3738),
.Y(n_3916)
);

HB1xp67_ASAP7_75t_L g3917 ( 
.A(n_3764),
.Y(n_3917)
);

CKINVDCx20_ASAP7_75t_R g3918 ( 
.A(n_3883),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3867),
.B(n_3739),
.Y(n_3919)
);

NAND2x1_ASAP7_75t_L g3920 ( 
.A(n_3884),
.B(n_3743),
.Y(n_3920)
);

O2A1O1Ixp33_ASAP7_75t_SL g3921 ( 
.A1(n_3913),
.A2(n_3748),
.B(n_3731),
.C(n_3685),
.Y(n_3921)
);

CKINVDCx11_ASAP7_75t_R g3922 ( 
.A(n_3821),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3867),
.B(n_3753),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3871),
.B(n_3753),
.Y(n_3924)
);

AOI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3855),
.A2(n_3683),
.B(n_3704),
.Y(n_3925)
);

OAI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3917),
.A2(n_3671),
.B(n_3754),
.Y(n_3926)
);

BUFx2_ASAP7_75t_L g3927 ( 
.A(n_3821),
.Y(n_3927)
);

AO32x2_ASAP7_75t_L g3928 ( 
.A1(n_3818),
.A2(n_3741),
.A3(n_3756),
.B1(n_3736),
.B2(n_3793),
.Y(n_3928)
);

AND2x4_ASAP7_75t_L g3929 ( 
.A(n_3813),
.B(n_3781),
.Y(n_3929)
);

AO32x2_ASAP7_75t_L g3930 ( 
.A1(n_3818),
.A2(n_3741),
.A3(n_3756),
.B1(n_3765),
.B2(n_3732),
.Y(n_3930)
);

INVxp67_ASAP7_75t_L g3931 ( 
.A(n_3879),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3871),
.B(n_3800),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3800),
.B(n_3753),
.Y(n_3933)
);

OAI211xp5_ASAP7_75t_L g3934 ( 
.A1(n_3856),
.A2(n_3740),
.B(n_3785),
.C(n_3605),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3868),
.B(n_3781),
.Y(n_3935)
);

AND2x4_ASAP7_75t_L g3936 ( 
.A(n_3813),
.B(n_3784),
.Y(n_3936)
);

AO21x2_ASAP7_75t_L g3937 ( 
.A1(n_3896),
.A2(n_3782),
.B(n_3779),
.Y(n_3937)
);

OR2x2_ASAP7_75t_L g3938 ( 
.A(n_3839),
.B(n_3750),
.Y(n_3938)
);

NOR2xp33_ASAP7_75t_L g3939 ( 
.A(n_3821),
.B(n_3786),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3868),
.B(n_3784),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3843),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3821),
.B(n_3724),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_3890),
.A2(n_3735),
.B(n_3764),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3907),
.B(n_3790),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_3821),
.B(n_3787),
.Y(n_3945)
);

OR2x2_ASAP7_75t_L g3946 ( 
.A(n_3839),
.B(n_3823),
.Y(n_3946)
);

INVx5_ASAP7_75t_SL g3947 ( 
.A(n_3884),
.Y(n_3947)
);

OR2x2_ASAP7_75t_L g3948 ( 
.A(n_3823),
.B(n_3869),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3843),
.Y(n_3949)
);

OR2x2_ASAP7_75t_L g3950 ( 
.A(n_3869),
.B(n_3750),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3869),
.B(n_3788),
.Y(n_3951)
);

AND2x2_ASAP7_75t_L g3952 ( 
.A(n_3907),
.B(n_3790),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3873),
.B(n_3794),
.Y(n_3953)
);

OAI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3862),
.A2(n_3754),
.B(n_3771),
.Y(n_3954)
);

AND2x2_ASAP7_75t_L g3955 ( 
.A(n_3873),
.B(n_3773),
.Y(n_3955)
);

AND2x4_ASAP7_75t_L g3956 ( 
.A(n_3830),
.B(n_3730),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3803),
.B(n_3746),
.Y(n_3957)
);

CKINVDCx5p33_ASAP7_75t_R g3958 ( 
.A(n_3861),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3884),
.Y(n_3959)
);

OAI21x1_ASAP7_75t_L g3960 ( 
.A1(n_3904),
.A2(n_3745),
.B(n_3768),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3890),
.A2(n_3676),
.B1(n_3789),
.B2(n_3792),
.Y(n_3961)
);

OR2x2_ASAP7_75t_L g3962 ( 
.A(n_3837),
.B(n_3778),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3884),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3874),
.B(n_3773),
.Y(n_3964)
);

INVx5_ASAP7_75t_SL g3965 ( 
.A(n_3830),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3874),
.B(n_3716),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3845),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3830),
.B(n_3769),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3845),
.Y(n_3969)
);

A2O1A1Ixp33_ASAP7_75t_L g3970 ( 
.A1(n_3802),
.A2(n_3771),
.B(n_3777),
.C(n_3737),
.Y(n_3970)
);

BUFx2_ASAP7_75t_L g3971 ( 
.A(n_3822),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3831),
.B(n_3716),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3831),
.B(n_3684),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3852),
.B(n_3684),
.Y(n_3974)
);

AND2x2_ASAP7_75t_L g3975 ( 
.A(n_3852),
.B(n_3775),
.Y(n_3975)
);

INVxp67_ASAP7_75t_L g3976 ( 
.A(n_3879),
.Y(n_3976)
);

NOR2x1_ASAP7_75t_SL g3977 ( 
.A(n_3890),
.B(n_3676),
.Y(n_3977)
);

INVx5_ASAP7_75t_SL g3978 ( 
.A(n_3857),
.Y(n_3978)
);

OAI21x1_ASAP7_75t_L g3979 ( 
.A1(n_3904),
.A2(n_3772),
.B(n_3701),
.Y(n_3979)
);

AOI22xp5_ASAP7_75t_L g3980 ( 
.A1(n_3806),
.A2(n_3763),
.B1(n_3769),
.B2(n_3777),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3887),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3842),
.B(n_3769),
.Y(n_3982)
);

AOI22xp5_ASAP7_75t_L g3983 ( 
.A1(n_3886),
.A2(n_3757),
.B1(n_3766),
.B2(n_3775),
.Y(n_3983)
);

NAND2xp33_ASAP7_75t_L g3984 ( 
.A(n_3822),
.B(n_3772),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3912),
.B(n_3701),
.Y(n_3985)
);

OAI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3862),
.A2(n_3772),
.B(n_3766),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3905),
.B(n_3567),
.Y(n_3987)
);

CKINVDCx14_ASAP7_75t_R g3988 ( 
.A(n_3861),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_3886),
.B(n_3769),
.Y(n_3989)
);

OR2x6_ASAP7_75t_L g3990 ( 
.A(n_3814),
.B(n_3737),
.Y(n_3990)
);

OR2x6_ASAP7_75t_L g3991 ( 
.A(n_3912),
.B(n_3763),
.Y(n_3991)
);

OA21x2_ASAP7_75t_L g3992 ( 
.A1(n_3882),
.A2(n_3816),
.B(n_3799),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3853),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3878),
.B(n_3714),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3887),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3905),
.B(n_3727),
.Y(n_3996)
);

OR2x6_ASAP7_75t_L g3997 ( 
.A(n_3799),
.B(n_3763),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3811),
.B(n_3727),
.Y(n_3998)
);

INVxp67_ASAP7_75t_L g3999 ( 
.A(n_3816),
.Y(n_3999)
);

OAI211xp5_ASAP7_75t_L g4000 ( 
.A1(n_3880),
.A2(n_3673),
.B(n_3762),
.C(n_3759),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_L g4001 ( 
.A(n_3829),
.B(n_3535),
.Y(n_4001)
);

INVx2_ASAP7_75t_SL g4002 ( 
.A(n_3857),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3854),
.Y(n_4003)
);

OAI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_3802),
.A2(n_3673),
.B(n_3759),
.Y(n_4004)
);

AO32x2_ASAP7_75t_L g4005 ( 
.A1(n_3849),
.A2(n_3762),
.A3(n_3634),
.B1(n_3643),
.B2(n_3673),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3878),
.B(n_3634),
.Y(n_4006)
);

NAND2xp33_ASAP7_75t_R g4007 ( 
.A(n_3806),
.B(n_3413),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_SL g4008 ( 
.A(n_3828),
.B(n_3475),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3806),
.A2(n_3386),
.B(n_3393),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3857),
.Y(n_4010)
);

OAI21xp5_ASAP7_75t_L g4011 ( 
.A1(n_3909),
.A2(n_3517),
.B(n_3439),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3811),
.B(n_3475),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3894),
.B(n_3495),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3894),
.B(n_3495),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3858),
.Y(n_4015)
);

AND2x2_ASAP7_75t_L g4016 ( 
.A(n_3911),
.B(n_3495),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3911),
.B(n_3487),
.Y(n_4017)
);

OA21x2_ASAP7_75t_L g4018 ( 
.A1(n_3882),
.A2(n_3386),
.B(n_3487),
.Y(n_4018)
);

AO21x2_ASAP7_75t_L g4019 ( 
.A1(n_3908),
.A2(n_3386),
.B(n_133),
.Y(n_4019)
);

INVx3_ASAP7_75t_L g4020 ( 
.A(n_3832),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3910),
.B(n_3487),
.Y(n_4021)
);

INVx3_ASAP7_75t_L g4022 ( 
.A(n_3832),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3849),
.B(n_3162),
.Y(n_4023)
);

AOI221xp5_ASAP7_75t_L g4024 ( 
.A1(n_3872),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.C(n_139),
.Y(n_4024)
);

OAI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3909),
.A2(n_134),
.B(n_140),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3914),
.B(n_140),
.Y(n_4026)
);

A2O1A1Ixp33_ASAP7_75t_L g4027 ( 
.A1(n_3851),
.A2(n_141),
.B(n_142),
.C(n_143),
.Y(n_4027)
);

BUFx4f_ASAP7_75t_L g4028 ( 
.A(n_3872),
.Y(n_4028)
);

NOR2xp33_ASAP7_75t_L g4029 ( 
.A(n_3820),
.B(n_141),
.Y(n_4029)
);

O2A1O1Ixp33_ASAP7_75t_L g4030 ( 
.A1(n_3848),
.A2(n_142),
.B(n_145),
.C(n_146),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3900),
.B(n_3820),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3857),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3892),
.B(n_146),
.Y(n_4033)
);

AND2x6_ASAP7_75t_L g4034 ( 
.A(n_3832),
.B(n_148),
.Y(n_4034)
);

OAI22xp5_ASAP7_75t_L g4035 ( 
.A1(n_3826),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3900),
.B(n_150),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3941),
.Y(n_4037)
);

HB1xp67_ASAP7_75t_L g4038 ( 
.A(n_3992),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3932),
.B(n_3898),
.Y(n_4039)
);

AO31x2_ASAP7_75t_L g4040 ( 
.A1(n_3977),
.A2(n_3906),
.A3(n_3891),
.B(n_3901),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3941),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3919),
.B(n_3898),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3949),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_3923),
.B(n_3898),
.Y(n_4044)
);

INVx1_ASAP7_75t_SL g4045 ( 
.A(n_3922),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3949),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3992),
.Y(n_4047)
);

OAI33xp33_ASAP7_75t_L g4048 ( 
.A1(n_3999),
.A2(n_3895),
.A3(n_3901),
.B1(n_3885),
.B2(n_3888),
.B3(n_3889),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3924),
.B(n_3876),
.Y(n_4049)
);

HB1xp67_ASAP7_75t_L g4050 ( 
.A(n_3988),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3967),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3977),
.Y(n_4052)
);

INVx5_ASAP7_75t_L g4053 ( 
.A(n_4034),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3933),
.B(n_3876),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3967),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3971),
.B(n_3906),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3981),
.B(n_3915),
.Y(n_4057)
);

NOR2x1_ASAP7_75t_L g4058 ( 
.A(n_3943),
.B(n_3857),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3969),
.Y(n_4059)
);

OR2x2_ASAP7_75t_L g4060 ( 
.A(n_3946),
.B(n_3877),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3927),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_4020),
.Y(n_4062)
);

BUFx3_ASAP7_75t_L g4063 ( 
.A(n_3918),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3995),
.B(n_3916),
.Y(n_4064)
);

HB1xp67_ASAP7_75t_L g4065 ( 
.A(n_3937),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_4020),
.Y(n_4066)
);

HB1xp67_ASAP7_75t_L g4067 ( 
.A(n_3937),
.Y(n_4067)
);

AND2x2_ASAP7_75t_L g4068 ( 
.A(n_3944),
.B(n_3877),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3952),
.B(n_3891),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_4022),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3969),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_4022),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3935),
.B(n_3900),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_4029),
.B(n_3895),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3940),
.B(n_3885),
.Y(n_4075)
);

AND2x2_ASAP7_75t_L g4076 ( 
.A(n_3975),
.B(n_3836),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_3948),
.B(n_3850),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3993),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3930),
.Y(n_4079)
);

AO21x2_ASAP7_75t_L g4080 ( 
.A1(n_3980),
.A2(n_3897),
.B(n_3826),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3930),
.Y(n_4081)
);

INVx2_ASAP7_75t_R g4082 ( 
.A(n_3930),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3965),
.B(n_3903),
.Y(n_4083)
);

OR2x2_ASAP7_75t_L g4084 ( 
.A(n_3957),
.B(n_3850),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3993),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_4003),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3965),
.B(n_3903),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_3953),
.B(n_3903),
.Y(n_4088)
);

CKINVDCx8_ASAP7_75t_R g4089 ( 
.A(n_4034),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3973),
.B(n_3903),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4003),
.Y(n_4091)
);

OA21x2_ASAP7_75t_L g4092 ( 
.A1(n_3961),
.A2(n_3897),
.B(n_3893),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_3994),
.B(n_3860),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4015),
.Y(n_4094)
);

HB1xp67_ASAP7_75t_L g4095 ( 
.A(n_3998),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4015),
.Y(n_4096)
);

NOR2x1_ASAP7_75t_L g4097 ( 
.A(n_3997),
.B(n_3893),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3974),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3978),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_4033),
.Y(n_4100)
);

BUFx2_ASAP7_75t_L g4101 ( 
.A(n_3991),
.Y(n_4101)
);

OR2x2_ASAP7_75t_L g4102 ( 
.A(n_3962),
.B(n_3860),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_4010),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_3929),
.B(n_3863),
.Y(n_4104)
);

INVxp67_ASAP7_75t_L g4105 ( 
.A(n_4034),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3978),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4032),
.Y(n_4107)
);

OR2x2_ASAP7_75t_L g4108 ( 
.A(n_3938),
.B(n_3875),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3929),
.B(n_3863),
.Y(n_4109)
);

BUFx3_ASAP7_75t_L g4110 ( 
.A(n_3958),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4034),
.B(n_3801),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4026),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_3936),
.B(n_3863),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_4002),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3921),
.A2(n_4007),
.B1(n_3945),
.B2(n_3934),
.Y(n_4115)
);

AOI221xp5_ASAP7_75t_L g4116 ( 
.A1(n_3925),
.A2(n_3807),
.B1(n_3805),
.B2(n_3846),
.C(n_3817),
.Y(n_4116)
);

INVx3_ASAP7_75t_L g4117 ( 
.A(n_3920),
.Y(n_4117)
);

NAND3xp33_ASAP7_75t_SL g4118 ( 
.A(n_3980),
.B(n_3902),
.C(n_3899),
.Y(n_4118)
);

AOI322xp5_ASAP7_75t_L g4119 ( 
.A1(n_4024),
.A2(n_3841),
.A3(n_3808),
.B1(n_3810),
.B2(n_3824),
.C1(n_3819),
.C2(n_3815),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_4036),
.B(n_3881),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_4012),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_4028),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3936),
.B(n_3955),
.Y(n_4123)
);

HB1xp67_ASAP7_75t_L g4124 ( 
.A(n_3931),
.Y(n_4124)
);

HB1xp67_ASAP7_75t_L g4125 ( 
.A(n_3976),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3959),
.Y(n_4126)
);

BUFx6f_ASAP7_75t_L g4127 ( 
.A(n_4028),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_3964),
.B(n_3899),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_3966),
.B(n_3902),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_4061),
.B(n_3982),
.Y(n_4130)
);

NAND3xp33_ASAP7_75t_L g4131 ( 
.A(n_4115),
.B(n_4027),
.C(n_4025),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_R g4132 ( 
.A(n_4089),
.B(n_3939),
.Y(n_4132)
);

AOI221xp5_ASAP7_75t_L g4133 ( 
.A1(n_4116),
.A2(n_4035),
.B1(n_3926),
.B2(n_3970),
.C(n_4030),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_4050),
.B(n_3996),
.Y(n_4134)
);

AOI221xp5_ASAP7_75t_L g4135 ( 
.A1(n_4118),
.A2(n_4125),
.B1(n_4124),
.B2(n_4048),
.C(n_4067),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_4045),
.B(n_3991),
.Y(n_4136)
);

HB1xp67_ASAP7_75t_L g4137 ( 
.A(n_4065),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_4110),
.B(n_3985),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_4061),
.B(n_4031),
.Y(n_4139)
);

OAI221xp5_ASAP7_75t_SL g4140 ( 
.A1(n_4119),
.A2(n_3950),
.B1(n_4000),
.B2(n_3951),
.C(n_4009),
.Y(n_4140)
);

NOR3xp33_ASAP7_75t_L g4141 ( 
.A(n_4122),
.B(n_4105),
.C(n_4101),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_4110),
.B(n_4013),
.Y(n_4142)
);

HB1xp67_ASAP7_75t_L g4143 ( 
.A(n_4038),
.Y(n_4143)
);

AOI221xp5_ASAP7_75t_L g4144 ( 
.A1(n_4126),
.A2(n_3954),
.B1(n_3986),
.B2(n_4004),
.C(n_3963),
.Y(n_4144)
);

OAI21xp33_ASAP7_75t_L g4145 ( 
.A1(n_4076),
.A2(n_3942),
.B(n_3983),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_4073),
.B(n_4014),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4121),
.B(n_4006),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4121),
.B(n_3989),
.Y(n_4148)
);

AND2x2_ASAP7_75t_SL g4149 ( 
.A(n_4101),
.B(n_3987),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_4095),
.B(n_3989),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4073),
.B(n_3997),
.Y(n_4151)
);

AND2x2_ASAP7_75t_SL g4152 ( 
.A(n_4127),
.B(n_3984),
.Y(n_4152)
);

NAND4xp25_ASAP7_75t_L g4153 ( 
.A(n_4122),
.B(n_4001),
.C(n_3968),
.D(n_4008),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4112),
.B(n_3956),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_4063),
.B(n_3972),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_4112),
.B(n_4076),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4114),
.B(n_3956),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_4114),
.B(n_4016),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_4063),
.B(n_3990),
.Y(n_4159)
);

OAI221xp5_ASAP7_75t_SL g4160 ( 
.A1(n_4079),
.A2(n_3928),
.B1(n_3990),
.B2(n_4005),
.C(n_3947),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_SL g4161 ( 
.A(n_4053),
.B(n_3947),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_4068),
.B(n_4017),
.Y(n_4162)
);

NAND3xp33_ASAP7_75t_L g4163 ( 
.A(n_4053),
.B(n_4011),
.C(n_4021),
.Y(n_4163)
);

OAI221xp5_ASAP7_75t_SL g4164 ( 
.A1(n_4079),
.A2(n_3928),
.B1(n_4005),
.B2(n_3865),
.C(n_3833),
.Y(n_4164)
);

OAI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_4058),
.A2(n_3865),
.B1(n_4023),
.B2(n_3881),
.Y(n_4165)
);

OAI21xp33_ASAP7_75t_L g4166 ( 
.A1(n_4039),
.A2(n_3960),
.B(n_3864),
.Y(n_4166)
);

OAI21xp33_ASAP7_75t_L g4167 ( 
.A1(n_4039),
.A2(n_3866),
.B(n_3859),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_SL g4168 ( 
.A1(n_4089),
.A2(n_3928),
.B1(n_4005),
.B2(n_4018),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_SL g4169 ( 
.A(n_4053),
.B(n_3979),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_4123),
.B(n_3875),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_4068),
.B(n_3870),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4098),
.B(n_3838),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_4098),
.B(n_3838),
.Y(n_4173)
);

OAI21xp5_ASAP7_75t_SL g4174 ( 
.A1(n_4127),
.A2(n_3834),
.B(n_3827),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4060),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_4049),
.B(n_3840),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4123),
.B(n_3840),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_4049),
.B(n_3844),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4053),
.B(n_4103),
.Y(n_4179)
);

AOI221xp5_ASAP7_75t_L g4180 ( 
.A1(n_4081),
.A2(n_4127),
.B1(n_4107),
.B2(n_4056),
.C(n_4074),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_4042),
.B(n_3844),
.Y(n_4181)
);

OA21x2_ASAP7_75t_L g4182 ( 
.A1(n_4081),
.A2(n_3847),
.B(n_3834),
.Y(n_4182)
);

NAND3xp33_ASAP7_75t_L g4183 ( 
.A(n_4053),
.B(n_4018),
.C(n_3835),
.Y(n_4183)
);

NOR2xp33_ASAP7_75t_L g4184 ( 
.A(n_4149),
.B(n_4127),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4134),
.B(n_4100),
.Y(n_4185)
);

OR2x2_ASAP7_75t_L g4186 ( 
.A(n_4143),
.B(n_4082),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4143),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4135),
.B(n_4082),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_4182),
.Y(n_4189)
);

INVx2_ASAP7_75t_SL g4190 ( 
.A(n_4161),
.Y(n_4190)
);

BUFx3_ASAP7_75t_L g4191 ( 
.A(n_4136),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_4130),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_4132),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_4146),
.B(n_4042),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_4182),
.Y(n_4195)
);

NAND5xp2_ASAP7_75t_L g4196 ( 
.A(n_4140),
.B(n_4087),
.C(n_4083),
.D(n_4088),
.E(n_4044),
.Y(n_4196)
);

NAND3xp33_ASAP7_75t_L g4197 ( 
.A(n_4140),
.B(n_4127),
.C(n_4047),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4137),
.Y(n_4198)
);

BUFx3_ASAP7_75t_L g4199 ( 
.A(n_4137),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4141),
.B(n_4099),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4155),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4175),
.Y(n_4202)
);

INVx5_ASAP7_75t_SL g4203 ( 
.A(n_4149),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4142),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4138),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4151),
.B(n_4044),
.Y(n_4206)
);

AOI22xp33_ASAP7_75t_L g4207 ( 
.A1(n_4131),
.A2(n_4088),
.B1(n_4090),
.B2(n_4083),
.Y(n_4207)
);

INVxp67_ASAP7_75t_SL g4208 ( 
.A(n_4161),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4168),
.Y(n_4209)
);

AO22x1_ASAP7_75t_L g4210 ( 
.A1(n_4141),
.A2(n_4047),
.B1(n_4097),
.B2(n_4117),
.Y(n_4210)
);

AOI221xp5_ASAP7_75t_L g4211 ( 
.A1(n_4133),
.A2(n_4111),
.B1(n_4096),
.B2(n_4094),
.C(n_4078),
.Y(n_4211)
);

OR2x2_ASAP7_75t_L g4212 ( 
.A(n_4156),
.B(n_4060),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_4159),
.B(n_4087),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4172),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_4181),
.Y(n_4215)
);

INVxp67_ASAP7_75t_SL g4216 ( 
.A(n_4150),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4152),
.B(n_4117),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4152),
.B(n_4117),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4173),
.Y(n_4219)
);

INVx2_ASAP7_75t_L g4220 ( 
.A(n_4183),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4170),
.B(n_4090),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_4177),
.B(n_4062),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4169),
.Y(n_4223)
);

AND2x4_ASAP7_75t_L g4224 ( 
.A(n_4157),
.B(n_4062),
.Y(n_4224)
);

OR2x2_ASAP7_75t_L g4225 ( 
.A(n_4176),
.B(n_4084),
.Y(n_4225)
);

OA21x2_ASAP7_75t_L g4226 ( 
.A1(n_4180),
.A2(n_4052),
.B(n_4099),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4132),
.B(n_4054),
.Y(n_4227)
);

OAI22xp33_ASAP7_75t_L g4228 ( 
.A1(n_4153),
.A2(n_4092),
.B1(n_4052),
.B2(n_4106),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4171),
.Y(n_4229)
);

AO21x2_ASAP7_75t_L g4230 ( 
.A1(n_4179),
.A2(n_4041),
.B(n_4037),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4139),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4148),
.Y(n_4232)
);

A2O1A1Ixp33_ASAP7_75t_SL g4233 ( 
.A1(n_4160),
.A2(n_4164),
.B(n_4106),
.C(n_4147),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4145),
.B(n_4054),
.Y(n_4234)
);

HB1xp67_ASAP7_75t_L g4235 ( 
.A(n_4162),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4186),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4191),
.B(n_4075),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4199),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4199),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4227),
.B(n_4154),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4199),
.Y(n_4241)
);

AND2x4_ASAP7_75t_L g4242 ( 
.A(n_4191),
.B(n_4066),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4227),
.B(n_4158),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4198),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4203),
.B(n_4120),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4198),
.Y(n_4246)
);

OR2x2_ASAP7_75t_L g4247 ( 
.A(n_4186),
.B(n_4178),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4189),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4198),
.Y(n_4249)
);

AND2x2_ASAP7_75t_L g4250 ( 
.A(n_4191),
.B(n_4075),
.Y(n_4250)
);

HB1xp67_ASAP7_75t_L g4251 ( 
.A(n_4192),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4220),
.B(n_4084),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4187),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4203),
.B(n_4194),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4194),
.B(n_4206),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4187),
.Y(n_4256)
);

NAND2x1_ASAP7_75t_L g4257 ( 
.A(n_4217),
.B(n_4092),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4206),
.B(n_4069),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_4203),
.B(n_4069),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4203),
.B(n_4234),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4189),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4213),
.B(n_4066),
.Y(n_4262)
);

AND2x2_ASAP7_75t_L g4263 ( 
.A(n_4213),
.B(n_4070),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4189),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4195),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4195),
.Y(n_4266)
);

NOR2xp67_ASAP7_75t_L g4267 ( 
.A(n_4190),
.B(n_4165),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4203),
.B(n_4070),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4234),
.B(n_4174),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4217),
.B(n_4072),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4195),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4218),
.B(n_4072),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4201),
.B(n_4167),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4230),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4257),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4255),
.B(n_4221),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4257),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4274),
.Y(n_4278)
);

OR2x2_ASAP7_75t_L g4279 ( 
.A(n_4251),
.B(n_4201),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_4255),
.B(n_4221),
.Y(n_4280)
);

OR2x2_ASAP7_75t_L g4281 ( 
.A(n_4240),
.B(n_4201),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4237),
.B(n_4204),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4236),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4237),
.B(n_4204),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_4242),
.B(n_4218),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4236),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4258),
.B(n_4204),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_4243),
.B(n_4205),
.Y(n_4288)
);

INVxp67_ASAP7_75t_L g4289 ( 
.A(n_4250),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4249),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4249),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4248),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4250),
.B(n_4205),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4248),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4258),
.B(n_4208),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4262),
.B(n_4263),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4262),
.B(n_4205),
.Y(n_4297)
);

NOR2xp33_ASAP7_75t_L g4298 ( 
.A(n_4238),
.B(n_4193),
.Y(n_4298)
);

NAND2x1_ASAP7_75t_L g4299 ( 
.A(n_4242),
.B(n_4222),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4265),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4299),
.Y(n_4301)
);

OR2x2_ASAP7_75t_L g4302 ( 
.A(n_4296),
.B(n_4209),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4275),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4275),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4277),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4276),
.B(n_4263),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4277),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4295),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_SL g4309 ( 
.A(n_4295),
.B(n_4184),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4280),
.Y(n_4310)
);

AOI211xp5_ASAP7_75t_L g4311 ( 
.A1(n_4283),
.A2(n_4196),
.B(n_4233),
.C(n_4197),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4287),
.B(n_4207),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4294),
.Y(n_4313)
);

HB1xp67_ASAP7_75t_L g4314 ( 
.A(n_4285),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4285),
.B(n_4242),
.Y(n_4315)
);

INVxp33_ASAP7_75t_L g4316 ( 
.A(n_4298),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4285),
.B(n_4270),
.Y(n_4317)
);

OAI322xp33_ASAP7_75t_L g4318 ( 
.A1(n_4286),
.A2(n_4188),
.A3(n_4209),
.B1(n_4220),
.B2(n_4197),
.C1(n_4252),
.C2(n_4247),
.Y(n_4318)
);

AOI32xp33_ASAP7_75t_L g4319 ( 
.A1(n_4298),
.A2(n_4188),
.A3(n_4220),
.B1(n_4209),
.B2(n_4228),
.Y(n_4319)
);

NAND2x1p5_ASAP7_75t_L g4320 ( 
.A(n_4279),
.B(n_4239),
.Y(n_4320)
);

AOI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_4311),
.A2(n_4267),
.B1(n_4216),
.B2(n_4190),
.Y(n_4321)
);

INVx2_ASAP7_75t_SL g4322 ( 
.A(n_4314),
.Y(n_4322)
);

XNOR2x1_ASAP7_75t_L g4323 ( 
.A(n_4312),
.B(n_4281),
.Y(n_4323)
);

NOR2xp33_ASAP7_75t_L g4324 ( 
.A(n_4309),
.B(n_4200),
.Y(n_4324)
);

XNOR2xp5_ASAP7_75t_L g4325 ( 
.A(n_4311),
.B(n_4235),
.Y(n_4325)
);

AOI22xp5_ASAP7_75t_L g4326 ( 
.A1(n_4310),
.A2(n_4306),
.B1(n_4211),
.B2(n_4226),
.Y(n_4326)
);

INVxp67_ASAP7_75t_L g4327 ( 
.A(n_4315),
.Y(n_4327)
);

XOR2x2_ASAP7_75t_L g4328 ( 
.A(n_4320),
.B(n_4269),
.Y(n_4328)
);

XNOR2xp5_ASAP7_75t_L g4329 ( 
.A(n_4316),
.B(n_4270),
.Y(n_4329)
);

INVxp67_ASAP7_75t_L g4330 ( 
.A(n_4317),
.Y(n_4330)
);

XOR2x2_ASAP7_75t_L g4331 ( 
.A(n_4320),
.B(n_4260),
.Y(n_4331)
);

INVx2_ASAP7_75t_SL g4332 ( 
.A(n_4301),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4308),
.B(n_4272),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4303),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4302),
.B(n_4272),
.Y(n_4335)
);

XNOR2xp5_ASAP7_75t_L g4336 ( 
.A(n_4304),
.B(n_4254),
.Y(n_4336)
);

XOR2x2_ASAP7_75t_L g4337 ( 
.A(n_4305),
.B(n_4259),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4322),
.B(n_4268),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4333),
.B(n_4297),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4329),
.Y(n_4340)
);

AND2x4_ASAP7_75t_L g4341 ( 
.A(n_4335),
.B(n_4241),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4324),
.B(n_4268),
.Y(n_4342)
);

INVx1_ASAP7_75t_SL g4343 ( 
.A(n_4331),
.Y(n_4343)
);

INVx1_ASAP7_75t_SL g4344 ( 
.A(n_4328),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4332),
.B(n_4232),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_4326),
.B(n_4289),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4336),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4321),
.B(n_4289),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_4327),
.B(n_4232),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4338),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4341),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4341),
.B(n_4319),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4345),
.Y(n_4353)
);

AOI21xp33_ASAP7_75t_L g4354 ( 
.A1(n_4343),
.A2(n_4245),
.B(n_4323),
.Y(n_4354)
);

NOR3xp33_ASAP7_75t_L g4355 ( 
.A(n_4344),
.B(n_4330),
.C(n_4318),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4349),
.B(n_4232),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4342),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4351),
.Y(n_4358)
);

HB1xp67_ASAP7_75t_L g4359 ( 
.A(n_4356),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4352),
.Y(n_4360)
);

OAI21xp33_ASAP7_75t_L g4361 ( 
.A1(n_4354),
.A2(n_4196),
.B(n_4185),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_SL g4362 ( 
.A(n_4355),
.B(n_4223),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4353),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4350),
.B(n_4244),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4357),
.Y(n_4365)
);

OAI221xp5_ASAP7_75t_L g4366 ( 
.A1(n_4355),
.A2(n_4226),
.B1(n_4273),
.B2(n_4282),
.C(n_4284),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4351),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4351),
.Y(n_4368)
);

INVxp67_ASAP7_75t_L g4369 ( 
.A(n_4351),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4351),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4361),
.B(n_4246),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4367),
.B(n_4231),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4358),
.B(n_4202),
.Y(n_4373)
);

OAI221xp5_ASAP7_75t_L g4374 ( 
.A1(n_4366),
.A2(n_4226),
.B1(n_4325),
.B2(n_4293),
.C(n_4346),
.Y(n_4374)
);

INVx3_ASAP7_75t_SL g4375 ( 
.A(n_4365),
.Y(n_4375)
);

NOR2xp33_ASAP7_75t_L g4376 ( 
.A(n_4369),
.B(n_4318),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4368),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4370),
.B(n_4202),
.Y(n_4378)
);

AND2x2_ASAP7_75t_L g4379 ( 
.A(n_4363),
.B(n_4231),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4360),
.B(n_4288),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4364),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4364),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_4362),
.B(n_4253),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4359),
.B(n_4256),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_L g4385 ( 
.A(n_4366),
.B(n_4339),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4367),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4367),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4367),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4367),
.Y(n_4389)
);

OAI22xp5_ASAP7_75t_L g4390 ( 
.A1(n_4366),
.A2(n_4226),
.B1(n_4252),
.B2(n_4223),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_4361),
.B(n_4294),
.Y(n_4391)
);

AOI22xp33_ASAP7_75t_L g4392 ( 
.A1(n_4361),
.A2(n_4223),
.B1(n_4224),
.B2(n_4215),
.Y(n_4392)
);

INVx2_ASAP7_75t_SL g4393 ( 
.A(n_4372),
.Y(n_4393)
);

AOI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4376),
.A2(n_4340),
.B1(n_4347),
.B2(n_4337),
.Y(n_4394)
);

OAI322xp33_ASAP7_75t_L g4395 ( 
.A1(n_4390),
.A2(n_4271),
.A3(n_4261),
.B1(n_4264),
.B2(n_4307),
.C1(n_4348),
.C2(n_4334),
.Y(n_4395)
);

AND4x1_ASAP7_75t_L g4396 ( 
.A(n_4380),
.B(n_4313),
.C(n_4300),
.D(n_4292),
.Y(n_4396)
);

OAI322xp33_ASAP7_75t_L g4397 ( 
.A1(n_4390),
.A2(n_4266),
.A3(n_4265),
.B1(n_4291),
.B2(n_4290),
.C1(n_4278),
.C2(n_4247),
.Y(n_4397)
);

OAI22xp5_ASAP7_75t_L g4398 ( 
.A1(n_4392),
.A2(n_4215),
.B1(n_4224),
.B2(n_4229),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4373),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4378),
.Y(n_4400)
);

INVx2_ASAP7_75t_SL g4401 ( 
.A(n_4379),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4383),
.Y(n_4402)
);

CKINVDCx5p33_ASAP7_75t_R g4403 ( 
.A(n_4375),
.Y(n_4403)
);

AOI22xp5_ASAP7_75t_L g4404 ( 
.A1(n_4386),
.A2(n_4224),
.B1(n_4215),
.B2(n_4266),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4377),
.Y(n_4405)
);

AOI22xp5_ASAP7_75t_L g4406 ( 
.A1(n_4387),
.A2(n_4224),
.B1(n_4222),
.B2(n_4229),
.Y(n_4406)
);

O2A1O1Ixp33_ASAP7_75t_L g4407 ( 
.A1(n_4374),
.A2(n_4278),
.B(n_4160),
.C(n_4164),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4384),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4391),
.Y(n_4409)
);

AOI22x1_ASAP7_75t_L g4410 ( 
.A1(n_4388),
.A2(n_4212),
.B1(n_4219),
.B2(n_4214),
.Y(n_4410)
);

AOI22xp5_ASAP7_75t_L g4411 ( 
.A1(n_4389),
.A2(n_4222),
.B1(n_4219),
.B2(n_4214),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4391),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4371),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4381),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4385),
.A2(n_4222),
.B1(n_4210),
.B2(n_4230),
.Y(n_4415)
);

OA22x2_ASAP7_75t_L g4416 ( 
.A1(n_4382),
.A2(n_4085),
.B1(n_4037),
.B2(n_4041),
.Y(n_4416)
);

AOI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4376),
.A2(n_4210),
.B1(n_4230),
.B2(n_4212),
.Y(n_4417)
);

AOI22xp5_ASAP7_75t_L g4418 ( 
.A1(n_4376),
.A2(n_4230),
.B1(n_4144),
.B2(n_4163),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_4406),
.B(n_4225),
.Y(n_4419)
);

NOR3xp33_ASAP7_75t_L g4420 ( 
.A(n_4414),
.B(n_4225),
.C(n_4166),
.Y(n_4420)
);

NOR2x1_ASAP7_75t_L g4421 ( 
.A(n_4395),
.B(n_4397),
.Y(n_4421)
);

OAI211xp5_ASAP7_75t_SL g4422 ( 
.A1(n_4394),
.A2(n_4091),
.B(n_4086),
.C(n_4085),
.Y(n_4422)
);

INVxp67_ASAP7_75t_L g4423 ( 
.A(n_4404),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_4407),
.A2(n_4092),
.B(n_4046),
.Y(n_4424)
);

NOR4xp25_ASAP7_75t_L g4425 ( 
.A(n_4409),
.B(n_4043),
.C(n_4071),
.D(n_4046),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4405),
.B(n_4129),
.Y(n_4426)
);

NOR2x1_ASAP7_75t_L g4427 ( 
.A(n_4412),
.B(n_4043),
.Y(n_4427)
);

AOI211x1_ASAP7_75t_L g4428 ( 
.A1(n_4396),
.A2(n_4071),
.B(n_4059),
.C(n_4055),
.Y(n_4428)
);

AOI211xp5_ASAP7_75t_L g4429 ( 
.A1(n_4398),
.A2(n_4051),
.B(n_4077),
.C(n_4113),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_4416),
.Y(n_4430)
);

AOI22xp5_ASAP7_75t_L g4431 ( 
.A1(n_4403),
.A2(n_4080),
.B1(n_4113),
.B2(n_4109),
.Y(n_4431)
);

AOI211x1_ASAP7_75t_L g4432 ( 
.A1(n_4413),
.A2(n_4109),
.B(n_4104),
.C(n_4057),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4411),
.B(n_4080),
.Y(n_4433)
);

NOR2x1_ASAP7_75t_L g4434 ( 
.A(n_4408),
.B(n_4080),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_4415),
.B(n_4064),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4410),
.Y(n_4436)
);

OAI21xp5_ASAP7_75t_L g4437 ( 
.A1(n_4417),
.A2(n_4104),
.B(n_4077),
.Y(n_4437)
);

BUFx4_ASAP7_75t_R g4438 ( 
.A(n_4393),
.Y(n_4438)
);

AOI22xp5_ASAP7_75t_L g4439 ( 
.A1(n_4418),
.A2(n_4128),
.B1(n_4129),
.B2(n_4102),
.Y(n_4439)
);

AOI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_4401),
.A2(n_4128),
.B1(n_4102),
.B2(n_4093),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_4402),
.B(n_4093),
.Y(n_4441)
);

NOR3xp33_ASAP7_75t_L g4442 ( 
.A(n_4399),
.B(n_4400),
.C(n_4108),
.Y(n_4442)
);

NOR2x1_ASAP7_75t_L g4443 ( 
.A(n_4427),
.B(n_4108),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4426),
.Y(n_4444)
);

NAND5xp2_ASAP7_75t_L g4445 ( 
.A(n_4420),
.B(n_151),
.C(n_152),
.D(n_153),
.E(n_154),
.Y(n_4445)
);

INVxp33_ASAP7_75t_L g4446 ( 
.A(n_4441),
.Y(n_4446)
);

NOR3x1_ASAP7_75t_L g4447 ( 
.A(n_4436),
.B(n_3851),
.C(n_152),
.Y(n_4447)
);

NOR2x1_ASAP7_75t_L g4448 ( 
.A(n_4421),
.B(n_153),
.Y(n_4448)
);

AOI21xp5_ASAP7_75t_L g4449 ( 
.A1(n_4433),
.A2(n_4040),
.B(n_3833),
.Y(n_4449)
);

NOR4xp75_ASAP7_75t_L g4450 ( 
.A(n_4435),
.B(n_4040),
.C(n_155),
.D(n_156),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4432),
.B(n_4424),
.Y(n_4451)
);

OAI211xp5_ASAP7_75t_L g4452 ( 
.A1(n_4423),
.A2(n_154),
.B(n_157),
.C(n_158),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4440),
.B(n_4419),
.Y(n_4453)
);

OAI222xp33_ASAP7_75t_R g4454 ( 
.A1(n_4430),
.A2(n_4040),
.B1(n_158),
.B2(n_159),
.C1(n_160),
.C2(n_161),
.Y(n_4454)
);

AOI211xp5_ASAP7_75t_L g4455 ( 
.A1(n_4422),
.A2(n_157),
.B(n_160),
.C(n_162),
.Y(n_4455)
);

NOR3x1_ASAP7_75t_L g4456 ( 
.A(n_4437),
.B(n_162),
.C(n_164),
.Y(n_4456)
);

NOR4xp25_ASAP7_75t_L g4457 ( 
.A(n_4438),
.B(n_4442),
.C(n_4428),
.D(n_4425),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_4434),
.Y(n_4458)
);

NAND4xp75_ASAP7_75t_L g4459 ( 
.A(n_4439),
.B(n_164),
.C(n_165),
.D(n_168),
.Y(n_4459)
);

NOR2x1_ASAP7_75t_L g4460 ( 
.A(n_4459),
.B(n_4429),
.Y(n_4460)
);

NOR3xp33_ASAP7_75t_L g4461 ( 
.A(n_4453),
.B(n_4431),
.C(n_169),
.Y(n_4461)
);

NAND3xp33_ASAP7_75t_L g4462 ( 
.A(n_4448),
.B(n_169),
.C(n_170),
.Y(n_4462)
);

NOR2x1_ASAP7_75t_L g4463 ( 
.A(n_4452),
.B(n_170),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4443),
.Y(n_4464)
);

NOR3xp33_ASAP7_75t_L g4465 ( 
.A(n_4444),
.B(n_171),
.C(n_172),
.Y(n_4465)
);

AND4x1_ASAP7_75t_L g4466 ( 
.A(n_4457),
.B(n_172),
.C(n_174),
.D(n_175),
.Y(n_4466)
);

NAND5xp2_ASAP7_75t_L g4467 ( 
.A(n_4446),
.B(n_175),
.C(n_176),
.D(n_178),
.E(n_179),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_4455),
.B(n_4040),
.Y(n_4468)
);

NAND4xp25_ASAP7_75t_L g4469 ( 
.A(n_4456),
.B(n_176),
.C(n_178),
.D(n_179),
.Y(n_4469)
);

NOR3x1_ASAP7_75t_L g4470 ( 
.A(n_4451),
.B(n_181),
.C(n_182),
.Y(n_4470)
);

NOR2x1_ASAP7_75t_L g4471 ( 
.A(n_4445),
.B(n_181),
.Y(n_4471)
);

OR2x6_ASAP7_75t_L g4472 ( 
.A(n_4458),
.B(n_3847),
.Y(n_4472)
);

OR2x2_ASAP7_75t_L g4473 ( 
.A(n_4449),
.B(n_4040),
.Y(n_4473)
);

NOR3xp33_ASAP7_75t_L g4474 ( 
.A(n_4454),
.B(n_4450),
.C(n_4447),
.Y(n_4474)
);

AOI222xp33_ASAP7_75t_L g4475 ( 
.A1(n_4464),
.A2(n_4468),
.B1(n_4462),
.B2(n_4460),
.C1(n_4463),
.C2(n_4471),
.Y(n_4475)
);

AOI221xp5_ASAP7_75t_L g4476 ( 
.A1(n_4461),
.A2(n_3835),
.B1(n_3827),
.B2(n_3797),
.C(n_3798),
.Y(n_4476)
);

BUFx2_ASAP7_75t_L g4477 ( 
.A(n_4469),
.Y(n_4477)
);

AOI221xp5_ASAP7_75t_L g4478 ( 
.A1(n_4474),
.A2(n_3795),
.B1(n_3796),
.B2(n_3797),
.C(n_3798),
.Y(n_4478)
);

AOI221xp5_ASAP7_75t_L g4479 ( 
.A1(n_4465),
.A2(n_3795),
.B1(n_3796),
.B2(n_3804),
.C(n_3809),
.Y(n_4479)
);

AOI211x1_ASAP7_75t_L g4480 ( 
.A1(n_4466),
.A2(n_183),
.B(n_184),
.C(n_185),
.Y(n_4480)
);

NAND3xp33_ASAP7_75t_L g4481 ( 
.A(n_4472),
.B(n_183),
.C(n_185),
.Y(n_4481)
);

OAI221xp5_ASAP7_75t_L g4482 ( 
.A1(n_4472),
.A2(n_3804),
.B1(n_3809),
.B2(n_3812),
.C(n_3825),
.Y(n_4482)
);

AOI321xp33_ASAP7_75t_L g4483 ( 
.A1(n_4473),
.A2(n_186),
.A3(n_187),
.B1(n_193),
.B2(n_194),
.C(n_195),
.Y(n_4483)
);

NAND3xp33_ASAP7_75t_L g4484 ( 
.A(n_4470),
.B(n_186),
.C(n_187),
.Y(n_4484)
);

AOI221xp5_ASAP7_75t_L g4485 ( 
.A1(n_4467),
.A2(n_3812),
.B1(n_3825),
.B2(n_197),
.C(n_198),
.Y(n_4485)
);

A2O1A1Ixp33_ASAP7_75t_L g4486 ( 
.A1(n_4464),
.A2(n_194),
.B(n_195),
.C(n_199),
.Y(n_4486)
);

BUFx8_ASAP7_75t_L g4487 ( 
.A(n_4464),
.Y(n_4487)
);

OAI21xp5_ASAP7_75t_L g4488 ( 
.A1(n_4471),
.A2(n_199),
.B(n_200),
.Y(n_4488)
);

NOR2x1_ASAP7_75t_L g4489 ( 
.A(n_4464),
.B(n_200),
.Y(n_4489)
);

AOI22xp5_ASAP7_75t_L g4490 ( 
.A1(n_4474),
.A2(n_4019),
.B1(n_203),
.B2(n_204),
.Y(n_4490)
);

AOI221xp5_ASAP7_75t_SL g4491 ( 
.A1(n_4464),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.C(n_205),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4471),
.Y(n_4492)
);

AOI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_4492),
.A2(n_4019),
.B1(n_207),
.B2(n_208),
.Y(n_4493)
);

NOR2xp67_ASAP7_75t_L g4494 ( 
.A(n_4481),
.B(n_206),
.Y(n_4494)
);

NOR2xp67_ASAP7_75t_L g4495 ( 
.A(n_4484),
.B(n_206),
.Y(n_4495)
);

AOI22xp5_ASAP7_75t_L g4496 ( 
.A1(n_4487),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_4496)
);

NOR2xp67_ASAP7_75t_L g4497 ( 
.A(n_4488),
.B(n_209),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4489),
.Y(n_4498)
);

NOR2xp67_ASAP7_75t_L g4499 ( 
.A(n_4480),
.B(n_210),
.Y(n_4499)
);

XNOR2xp5_ASAP7_75t_L g4500 ( 
.A(n_4485),
.B(n_212),
.Y(n_4500)
);

NAND3xp33_ASAP7_75t_L g4501 ( 
.A(n_4487),
.B(n_212),
.C(n_214),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4483),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4477),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4486),
.Y(n_4504)
);

HB1xp67_ASAP7_75t_L g4505 ( 
.A(n_4491),
.Y(n_4505)
);

NOR2x2_ASAP7_75t_L g4506 ( 
.A(n_4475),
.B(n_214),
.Y(n_4506)
);

AOI22xp5_ASAP7_75t_L g4507 ( 
.A1(n_4478),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_4507)
);

AOI22xp33_ASAP7_75t_SL g4508 ( 
.A1(n_4482),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_4508)
);

AOI22xp5_ASAP7_75t_L g4509 ( 
.A1(n_4476),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_4509)
);

AOI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4503),
.A2(n_4479),
.B1(n_4490),
.B2(n_223),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4508),
.B(n_221),
.Y(n_4511)
);

NOR2xp33_ASAP7_75t_L g4512 ( 
.A(n_4502),
.B(n_221),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_4499),
.B(n_222),
.Y(n_4513)
);

NAND4xp75_ASAP7_75t_L g4514 ( 
.A(n_4495),
.B(n_223),
.C(n_224),
.D(n_225),
.Y(n_4514)
);

OAI322xp33_ASAP7_75t_L g4515 ( 
.A1(n_4498),
.A2(n_226),
.A3(n_227),
.B1(n_228),
.B2(n_229),
.C1(n_283),
.C2(n_285),
.Y(n_4515)
);

NOR2xp33_ASAP7_75t_L g4516 ( 
.A(n_4505),
.B(n_4504),
.Y(n_4516)
);

NAND4xp25_ASAP7_75t_L g4517 ( 
.A(n_4507),
.B(n_226),
.C(n_286),
.D(n_289),
.Y(n_4517)
);

HB1xp67_ASAP7_75t_L g4518 ( 
.A(n_4501),
.Y(n_4518)
);

AND2x4_ASAP7_75t_L g4519 ( 
.A(n_4497),
.B(n_291),
.Y(n_4519)
);

HB1xp67_ASAP7_75t_L g4520 ( 
.A(n_4494),
.Y(n_4520)
);

NOR3xp33_ASAP7_75t_L g4521 ( 
.A(n_4512),
.B(n_4506),
.C(n_4509),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4519),
.B(n_4500),
.Y(n_4522)
);

OAI22x1_ASAP7_75t_L g4523 ( 
.A1(n_4510),
.A2(n_4496),
.B1(n_4493),
.B2(n_297),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_SL g4524 ( 
.A(n_4513),
.B(n_293),
.Y(n_4524)
);

NAND3xp33_ASAP7_75t_L g4525 ( 
.A(n_4516),
.B(n_294),
.C(n_300),
.Y(n_4525)
);

NAND3xp33_ASAP7_75t_L g4526 ( 
.A(n_4518),
.B(n_302),
.C(n_303),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4524),
.Y(n_4527)
);

NOR3xp33_ASAP7_75t_L g4528 ( 
.A(n_4522),
.B(n_4520),
.C(n_4511),
.Y(n_4528)
);

INVx2_ASAP7_75t_SL g4529 ( 
.A(n_4523),
.Y(n_4529)
);

AOI22xp5_ASAP7_75t_L g4530 ( 
.A1(n_4528),
.A2(n_4521),
.B1(n_4514),
.B2(n_4517),
.Y(n_4530)
);

AO21x2_ASAP7_75t_L g4531 ( 
.A1(n_4527),
.A2(n_4519),
.B(n_4525),
.Y(n_4531)
);

NAND4xp75_ASAP7_75t_L g4532 ( 
.A(n_4530),
.B(n_4529),
.C(n_4526),
.D(n_4515),
.Y(n_4532)
);

OAI221xp5_ASAP7_75t_L g4533 ( 
.A1(n_4532),
.A2(n_4531),
.B1(n_307),
.B2(n_308),
.C(n_310),
.Y(n_4533)
);

XOR2xp5_ASAP7_75t_L g4534 ( 
.A(n_4533),
.B(n_305),
.Y(n_4534)
);

AO22x2_ASAP7_75t_L g4535 ( 
.A1(n_4534),
.A2(n_312),
.B1(n_313),
.B2(n_316),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4535),
.B(n_320),
.Y(n_4536)
);

AND3x4_ASAP7_75t_L g4537 ( 
.A(n_4536),
.B(n_323),
.C(n_324),
.Y(n_4537)
);

AO21x2_ASAP7_75t_L g4538 ( 
.A1(n_4537),
.A2(n_328),
.B(n_329),
.Y(n_4538)
);

OAI321xp33_ASAP7_75t_L g4539 ( 
.A1(n_4538),
.A2(n_332),
.A3(n_334),
.B1(n_335),
.B2(n_336),
.C(n_337),
.Y(n_4539)
);

AOI22xp5_ASAP7_75t_SL g4540 ( 
.A1(n_4539),
.A2(n_338),
.B1(n_345),
.B2(n_347),
.Y(n_4540)
);

AO21x2_ASAP7_75t_L g4541 ( 
.A1(n_4540),
.A2(n_348),
.B(n_352),
.Y(n_4541)
);

OAI221xp5_ASAP7_75t_R g4542 ( 
.A1(n_4541),
.A2(n_366),
.B1(n_369),
.B2(n_370),
.C(n_372),
.Y(n_4542)
);

AOI21xp5_ASAP7_75t_L g4543 ( 
.A1(n_4542),
.A2(n_1467),
.B(n_1457),
.Y(n_4543)
);

AOI211xp5_ASAP7_75t_L g4544 ( 
.A1(n_4543),
.A2(n_375),
.B(n_381),
.C(n_388),
.Y(n_4544)
);


endmodule