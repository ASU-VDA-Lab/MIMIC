module fake_jpeg_30765_n_82 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_7),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_11),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_27),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_20),
.Y(n_37)
);

XNOR2x1_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_19),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_12),
.B(n_15),
.C(n_20),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_44),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_15),
.C(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_14),
.B1(n_10),
.B2(n_2),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_57),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_44),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_46),
.B1(n_41),
.B2(n_39),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_48),
.C(n_43),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_65),
.C(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_63),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_49),
.C(n_10),
.Y(n_65)
);

NOR2xp67_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_61),
.B1(n_70),
.B2(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_76),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_72),
.C(n_77),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_81),
.B(n_6),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_73),
.C(n_74),
.Y(n_81)
);


endmodule