module real_jpeg_24302_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_71),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_2),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_3),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_66),
.C(n_88),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_5),
.B(n_60),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_5),
.A2(n_102),
.B1(n_172),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_5),
.B(n_98),
.Y(n_211)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_77),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_8),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_47),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_9),
.A2(n_47),
.B1(n_65),
.B2(n_66),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_9),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_198)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_10),
.B(n_29),
.C(n_32),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_59),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_59),
.B1(n_65),
.B2(n_66),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_15),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_136),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_19),
.B(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_100),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_20),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_61),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_44),
.C(n_82),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_38),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_79),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_25),
.A2(n_41),
.B1(n_98),
.B2(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_27),
.A2(n_30),
.B(n_79),
.C(n_81),
.Y(n_78)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_29),
.B(n_51),
.C(n_55),
.Y(n_190)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g189 ( 
.A(n_30),
.B(n_80),
.CON(n_189),
.SN(n_189)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_38),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_42),
.B(n_80),
.CON(n_79),
.SN(n_79)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_57),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_49),
.B1(n_60),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_48),
.A2(n_53),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_49),
.A2(n_58),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_49),
.A2(n_60),
.B1(n_189),
.B2(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_52),
.A2(n_54),
.B(n_188),
.C(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_132),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_55),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_55),
.B(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_78),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_62),
.A2(n_63),
.B1(n_78),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_76),
.Y(n_63)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_64),
.B(n_105),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_64),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_66),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_65),
.B(n_178),
.Y(n_177)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_70),
.A2(n_119),
.B(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_75),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_78),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_80),
.B(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_80),
.B(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_83),
.B(n_100),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.C(n_97),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_84),
.B(n_95),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_122),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_85),
.A2(n_122),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_86),
.A2(n_90),
.B1(n_150),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_86),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_91),
.B(n_122),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_97),
.B(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_115),
.B(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_102),
.A2(n_164),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_102),
.A2(n_104),
.B(n_118),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_133),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_125),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_120),
.B2(n_124),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_238),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_234),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_224),
.B(n_233),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_201),
.B(n_223),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_183),
.B(n_200),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_160),
.B(n_182),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_147),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_155),
.C(n_158),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_168),
.B(n_181),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_167),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_180),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_199),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_193),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_194),
.C(n_196),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_215),
.B2(n_216),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_218),
.C(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_210),
.C(n_213),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_232),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_229),
.C(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);


endmodule