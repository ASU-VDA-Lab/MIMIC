module real_aes_15417_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1800;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_SL g1489 ( .A1(n_0), .A2(n_262), .B1(n_527), .B2(n_1490), .Y(n_1489) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_0), .A2(n_161), .B1(n_431), .B2(n_1523), .Y(n_1526) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_1), .A2(n_61), .B1(n_694), .B2(n_1326), .Y(n_1325) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_1), .Y(n_1344) );
INVx1_ASAP7_75t_L g1274 ( .A(n_2), .Y(n_1274) );
INVx1_ASAP7_75t_L g969 ( .A(n_3), .Y(n_969) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_4), .A2(n_251), .B1(n_532), .B2(n_1341), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_4), .A2(n_339), .B1(n_399), .B2(n_1022), .Y(n_1392) );
INVx1_ASAP7_75t_L g376 ( .A(n_5), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_5), .B(n_386), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_6), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_7), .A2(n_247), .B1(n_532), .B2(n_928), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_7), .A2(n_190), .B1(n_434), .B2(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g1177 ( .A(n_8), .Y(n_1177) );
INVx1_ASAP7_75t_L g1504 ( .A(n_9), .Y(n_1504) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_9), .A2(n_181), .B1(n_891), .B2(n_936), .Y(n_1514) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_10), .A2(n_60), .B1(n_378), .B2(n_752), .Y(n_1059) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_10), .A2(n_60), .B1(n_707), .B2(n_731), .Y(n_1098) );
OAI22xp33_ASAP7_75t_SL g837 ( .A1(n_11), .A2(n_346), .B1(n_482), .B2(n_838), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_11), .A2(n_172), .B1(n_444), .B2(n_465), .Y(n_853) );
INVx1_ASAP7_75t_L g919 ( .A(n_12), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_12), .A2(n_247), .B1(n_404), .B2(n_948), .Y(n_954) );
INVx1_ASAP7_75t_L g1281 ( .A(n_13), .Y(n_1281) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_14), .A2(n_200), .B1(n_1547), .B2(n_1561), .Y(n_1573) );
INVx1_ASAP7_75t_L g1510 ( .A(n_15), .Y(n_1510) );
INVx1_ASAP7_75t_L g1306 ( .A(n_16), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g1782 ( .A(n_17), .Y(n_1782) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_18), .A2(n_45), .B1(n_707), .B2(n_731), .Y(n_730) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_18), .A2(n_45), .B1(n_378), .B2(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_19), .A2(n_94), .B1(n_1547), .B2(n_1549), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_20), .A2(n_113), .B1(n_527), .B2(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1521 ( .A(n_20), .Y(n_1521) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_21), .Y(n_862) );
XOR2x2_ASAP7_75t_L g1396 ( .A(n_22), .B(n_1397), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_22), .A2(n_341), .B1(n_1539), .B2(n_1544), .Y(n_1632) );
OAI22xp5_ASAP7_75t_L g1757 ( .A1(n_23), .A2(n_319), .B1(n_747), .B2(n_1031), .Y(n_1757) );
OAI22xp5_ASAP7_75t_L g1760 ( .A1(n_23), .A2(n_319), .B1(n_721), .B2(n_722), .Y(n_1760) );
INVx2_ASAP7_75t_L g425 ( .A(n_24), .Y(n_425) );
INVx1_ASAP7_75t_L g456 ( .A(n_25), .Y(n_456) );
INVx1_ASAP7_75t_L g450 ( .A(n_26), .Y(n_450) );
XNOR2xp5_ASAP7_75t_L g1297 ( .A(n_27), .B(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g645 ( .A(n_28), .Y(n_645) );
INVx1_ASAP7_75t_L g589 ( .A(n_29), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_30), .A2(n_87), .B1(n_412), .B2(n_416), .C(n_421), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_30), .A2(n_43), .B1(n_543), .B2(n_546), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g1581 ( .A1(n_31), .A2(n_209), .B1(n_1539), .B2(n_1544), .Y(n_1581) );
INVx1_ASAP7_75t_L g1211 ( .A(n_32), .Y(n_1211) );
INVx1_ASAP7_75t_L g637 ( .A(n_33), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_34), .A2(n_687), .B(n_690), .C(n_696), .Y(n_686) );
INVx1_ASAP7_75t_L g719 ( .A(n_34), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_35), .A2(n_86), .B1(n_446), .B2(n_465), .C(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g997 ( .A(n_35), .Y(n_997) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_36), .Y(n_371) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_36), .B(n_369), .Y(n_1540) );
AOI22xp33_ASAP7_75t_L g1630 ( .A1(n_37), .A2(n_186), .B1(n_1547), .B2(n_1631), .Y(n_1630) );
XOR2xp5_ASAP7_75t_L g1798 ( .A(n_38), .B(n_1799), .Y(n_1798) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_39), .A2(n_199), .B1(n_1547), .B2(n_1549), .Y(n_1570) );
OAI22xp33_ASAP7_75t_SL g1163 ( .A1(n_40), .A2(n_162), .B1(n_747), .B2(n_1031), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_40), .A2(n_162), .B1(n_721), .B2(n_1042), .Y(n_1166) );
AOI22xp33_ASAP7_75t_SL g1431 ( .A1(n_41), .A2(n_258), .B1(n_532), .B2(n_1427), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_41), .A2(n_151), .B1(n_946), .B2(n_1434), .Y(n_1437) );
INVx1_ASAP7_75t_L g1125 ( .A(n_42), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_43), .A2(n_76), .B1(n_412), .B2(n_416), .C(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_SL g1324 ( .A(n_44), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_44), .A2(n_61), .B1(n_845), .B2(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1011 ( .A(n_46), .Y(n_1011) );
INVx1_ASAP7_75t_L g1077 ( .A(n_47), .Y(n_1077) );
INVx1_ASAP7_75t_L g1234 ( .A(n_48), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_48), .A2(n_352), .B1(n_699), .B2(n_701), .Y(n_1242) );
INVx1_ASAP7_75t_L g757 ( .A(n_49), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_50), .A2(n_295), .B1(n_492), .B2(n_493), .Y(n_1366) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_50), .A2(n_295), .B1(n_446), .B2(n_467), .Y(n_1369) );
AOI22xp5_ASAP7_75t_L g1546 ( .A1(n_51), .A2(n_158), .B1(n_1547), .B2(n_1549), .Y(n_1546) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_52), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_53), .Y(n_915) );
INVx1_ASAP7_75t_L g435 ( .A(n_54), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_54), .A2(n_252), .B1(n_527), .B2(n_532), .Y(n_526) );
INVx1_ASAP7_75t_L g1475 ( .A(n_55), .Y(n_1475) );
INVx1_ASAP7_75t_L g972 ( .A(n_56), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_57), .A2(n_255), .B1(n_1323), .B2(n_1377), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_57), .A2(n_93), .B1(n_416), .B2(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1203 ( .A(n_58), .Y(n_1203) );
XNOR2xp5_ASAP7_75t_L g1254 ( .A(n_59), .B(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g604 ( .A(n_62), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_63), .B(n_424), .Y(n_984) );
INVxp67_ASAP7_75t_SL g993 ( .A(n_63), .Y(n_993) );
OAI211xp5_ASAP7_75t_SL g732 ( .A1(n_64), .A2(n_712), .B(n_713), .C(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g745 ( .A(n_64), .Y(n_745) );
OAI211xp5_ASAP7_75t_L g830 ( .A1(n_65), .A2(n_560), .B(n_831), .C(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g852 ( .A(n_65), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_66), .A2(n_167), .B1(n_721), .B2(n_722), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_66), .A2(n_167), .B1(n_747), .B2(n_748), .Y(n_746) );
OAI22xp33_ASAP7_75t_L g1446 ( .A1(n_67), .A2(n_227), .B1(n_446), .B2(n_722), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_67), .A2(n_227), .B1(n_700), .B2(n_1459), .Y(n_1458) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_68), .Y(n_799) );
INVx1_ASAP7_75t_L g1328 ( .A(n_69), .Y(n_1328) );
INVx1_ASAP7_75t_L g1472 ( .A(n_70), .Y(n_1472) );
OAI222xp33_ASAP7_75t_L g903 ( .A1(n_71), .A2(n_175), .B1(n_483), .B2(n_836), .C1(n_904), .C2(n_905), .Y(n_903) );
OAI222xp33_ASAP7_75t_L g934 ( .A1(n_71), .A2(n_175), .B1(n_215), .B2(n_935), .C1(n_936), .C2(n_937), .Y(n_934) );
OAI211xp5_ASAP7_75t_L g1026 ( .A1(n_72), .A2(n_739), .B(n_742), .C(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1040 ( .A(n_72), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1145 ( .A1(n_73), .A2(n_305), .B1(n_378), .B2(n_752), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_73), .A2(n_305), .B1(n_731), .B2(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g695 ( .A(n_74), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g711 ( .A1(n_74), .A2(n_712), .B(n_713), .C(n_714), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_75), .A2(n_179), .B1(n_444), .B2(n_988), .Y(n_987) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_75), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_76), .A2(n_87), .B1(n_535), .B2(n_537), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_77), .Y(n_871) );
INVx1_ASAP7_75t_L g1329 ( .A(n_78), .Y(n_1329) );
INVx1_ASAP7_75t_L g770 ( .A(n_79), .Y(n_770) );
INVx1_ASAP7_75t_L g1319 ( .A(n_80), .Y(n_1319) );
INVx1_ASAP7_75t_L g1487 ( .A(n_81), .Y(n_1487) );
OAI211xp5_ASAP7_75t_L g1362 ( .A1(n_82), .A2(n_511), .B(n_918), .C(n_1363), .Y(n_1362) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_82), .A2(n_197), .B1(n_800), .B2(n_1346), .C(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1260 ( .A(n_83), .Y(n_1260) );
OAI211xp5_ASAP7_75t_L g1267 ( .A1(n_83), .A2(n_712), .B(n_713), .C(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g971 ( .A(n_84), .Y(n_971) );
INVx1_ASAP7_75t_L g1188 ( .A(n_85), .Y(n_1188) );
OAI22xp33_ASAP7_75t_L g999 ( .A1(n_86), .A2(n_179), .B1(n_482), .B2(n_568), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_88), .A2(n_187), .B1(n_444), .B2(n_446), .Y(n_443) );
INVx1_ASAP7_75t_L g480 ( .A(n_88), .Y(n_480) );
INVx1_ASAP7_75t_L g650 ( .A(n_89), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_90), .A2(n_268), .B1(n_482), .B2(n_493), .Y(n_881) );
OAI22xp5_ASAP7_75t_SL g889 ( .A1(n_90), .A2(n_126), .B1(n_444), .B2(n_467), .Y(n_889) );
INVx1_ASAP7_75t_L g769 ( .A(n_91), .Y(n_769) );
INVx1_ASAP7_75t_L g986 ( .A(n_92), .Y(n_986) );
AOI22xp33_ASAP7_75t_SL g1380 ( .A1(n_93), .A2(n_351), .B1(n_532), .B2(n_1381), .Y(n_1380) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_95), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_96), .Y(n_860) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_97), .A2(n_153), .B1(n_378), .B2(n_568), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_97), .A2(n_153), .B1(n_707), .B2(n_709), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_98), .Y(n_798) );
OAI211xp5_ASAP7_75t_L g1447 ( .A1(n_99), .A2(n_453), .B(n_667), .C(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1456 ( .A(n_99), .Y(n_1456) );
INVx1_ASAP7_75t_L g460 ( .A(n_100), .Y(n_460) );
OAI22xp33_ASAP7_75t_SL g1065 ( .A1(n_101), .A2(n_267), .B1(n_699), .B2(n_1066), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_101), .A2(n_267), .B1(n_722), .B2(n_1044), .Y(n_1102) );
XOR2xp5_ASAP7_75t_L g793 ( .A(n_102), .B(n_794), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g1555 ( .A1(n_102), .A2(n_208), .B1(n_1539), .B2(n_1544), .Y(n_1555) );
XNOR2x2_ASAP7_75t_SL g1443 ( .A(n_103), .B(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1308 ( .A(n_104), .Y(n_1308) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_104), .A2(n_293), .B1(n_1335), .B2(n_1341), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_105), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_106), .A2(n_218), .B1(n_936), .B2(n_1406), .Y(n_1405) );
INVxp67_ASAP7_75t_SL g1416 ( .A(n_106), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_107), .A2(n_291), .B1(n_532), .B2(n_1427), .Y(n_1426) );
AOI22xp33_ASAP7_75t_SL g1438 ( .A1(n_107), .A2(n_254), .B1(n_431), .B2(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1131 ( .A(n_108), .Y(n_1131) );
INVx1_ASAP7_75t_L g369 ( .A(n_109), .Y(n_369) );
INVx1_ASAP7_75t_L g1084 ( .A(n_110), .Y(n_1084) );
INVx1_ASAP7_75t_L g1315 ( .A(n_111), .Y(n_1315) );
INVxp67_ASAP7_75t_SL g1403 ( .A(n_112), .Y(n_1403) );
OAI22xp33_ASAP7_75t_L g1417 ( .A1(n_112), .A2(n_218), .B1(n_694), .B2(n_1326), .Y(n_1417) );
INVxp67_ASAP7_75t_SL g1525 ( .A(n_113), .Y(n_1525) );
XOR2xp5_ASAP7_75t_L g895 ( .A(n_114), .B(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g1277 ( .A(n_115), .Y(n_1277) );
INVx1_ASAP7_75t_L g1161 ( .A(n_116), .Y(n_1161) );
INVx1_ASAP7_75t_L g1505 ( .A(n_117), .Y(n_1505) );
INVx1_ASAP7_75t_L g1118 ( .A(n_118), .Y(n_1118) );
INVx1_ASAP7_75t_L g1063 ( .A(n_119), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g1559 ( .A1(n_120), .A2(n_318), .B1(n_1539), .B2(n_1544), .Y(n_1559) );
INVx1_ASAP7_75t_L g1304 ( .A(n_121), .Y(n_1304) );
INVx1_ASAP7_75t_L g1180 ( .A(n_122), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_123), .A2(n_183), .B1(n_573), .B2(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1050 ( .A(n_123), .Y(n_1050) );
INVx1_ASAP7_75t_L g597 ( .A(n_124), .Y(n_597) );
OAI22xp33_ASAP7_75t_SL g886 ( .A1(n_125), .A2(n_126), .B1(n_492), .B2(n_568), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_125), .A2(n_131), .B1(n_850), .B2(n_851), .Y(n_893) );
INVx1_ASAP7_75t_L g774 ( .A(n_127), .Y(n_774) );
INVx1_ASAP7_75t_L g602 ( .A(n_128), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_129), .A2(n_211), .B1(n_1547), .B2(n_1549), .Y(n_1580) );
CKINVDCx5p33_ASAP7_75t_R g1778 ( .A(n_130), .Y(n_1778) );
INVx1_ASAP7_75t_L g885 ( .A(n_131), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_132), .A2(n_345), .B1(n_444), .B2(n_1452), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_132), .A2(n_345), .B1(n_482), .B2(n_752), .Y(n_1460) );
INVx1_ASAP7_75t_L g1474 ( .A(n_133), .Y(n_1474) );
INVx1_ASAP7_75t_L g599 ( .A(n_134), .Y(n_599) );
AOI31xp33_ASAP7_75t_L g396 ( .A1(n_135), .A2(n_397), .A3(n_442), .B(n_478), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g520 ( .A(n_135), .B(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_135), .Y(n_549) );
INVx1_ASAP7_75t_L g1488 ( .A(n_136), .Y(n_1488) );
AOI22xp5_ASAP7_75t_L g1574 ( .A1(n_137), .A2(n_221), .B1(n_1539), .B2(n_1544), .Y(n_1574) );
INVx1_ASAP7_75t_L g639 ( .A(n_138), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g1781 ( .A(n_139), .Y(n_1781) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_140), .Y(n_865) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_141), .A2(n_739), .B(n_742), .C(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1170 ( .A(n_141), .Y(n_1170) );
INVx1_ASAP7_75t_L g1162 ( .A(n_142), .Y(n_1162) );
OAI211xp5_ASAP7_75t_L g1167 ( .A1(n_142), .A2(n_453), .B(n_1168), .C(n_1169), .Y(n_1167) );
INVx1_ASAP7_75t_L g763 ( .A(n_143), .Y(n_763) );
INVx1_ASAP7_75t_L g734 ( .A(n_144), .Y(n_734) );
INVx1_ASAP7_75t_L g652 ( .A(n_145), .Y(n_652) );
INVx1_ASAP7_75t_L g1471 ( .A(n_146), .Y(n_1471) );
INVx1_ASAP7_75t_L g1178 ( .A(n_147), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_148), .Y(n_802) );
OAI211xp5_ASAP7_75t_L g1140 ( .A1(n_149), .A2(n_741), .B(n_742), .C(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1152 ( .A(n_149), .Y(n_1152) );
CKINVDCx20_ASAP7_75t_R g1284 ( .A(n_150), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_151), .A2(n_332), .B1(n_1422), .B2(n_1425), .Y(n_1421) );
INVx1_ASAP7_75t_L g1142 ( .A(n_152), .Y(n_1142) );
INVx1_ASAP7_75t_L g967 ( .A(n_154), .Y(n_967) );
INVx1_ASAP7_75t_L g595 ( .A(n_155), .Y(n_595) );
INVx1_ASAP7_75t_L g1259 ( .A(n_156), .Y(n_1259) );
INVx1_ASAP7_75t_L g1064 ( .A(n_157), .Y(n_1064) );
OAI211xp5_ASAP7_75t_L g1099 ( .A1(n_157), .A2(n_712), .B(n_713), .C(n_1100), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_159), .A2(n_290), .B1(n_747), .B2(n_1031), .Y(n_1144) );
OAI22xp33_ASAP7_75t_L g1153 ( .A1(n_159), .A2(n_290), .B1(n_721), .B2(n_1042), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g1492 ( .A(n_160), .Y(n_1492) );
AOI22xp33_ASAP7_75t_SL g1522 ( .A1(n_160), .A2(n_262), .B1(n_983), .B2(n_1523), .Y(n_1522) );
INVxp67_ASAP7_75t_SL g1493 ( .A(n_161), .Y(n_1493) );
CKINVDCx5p33_ASAP7_75t_R g809 ( .A(n_163), .Y(n_809) );
XNOR2xp5_ASAP7_75t_L g1483 ( .A(n_164), .B(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1187 ( .A(n_165), .Y(n_1187) );
INVx1_ASAP7_75t_L g1130 ( .A(n_166), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_168), .A2(n_245), .B1(n_699), .B2(n_1066), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_168), .A2(n_245), .B1(n_1265), .B2(n_1266), .Y(n_1264) );
INVx1_ASAP7_75t_L g735 ( .A(n_169), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_169), .A2(n_739), .B(n_742), .C(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g1283 ( .A(n_170), .Y(n_1283) );
INVx1_ASAP7_75t_L g1075 ( .A(n_171), .Y(n_1075) );
OAI22xp33_ASAP7_75t_SL g840 ( .A1(n_172), .A2(n_306), .B1(n_700), .B2(n_752), .Y(n_840) );
INVx1_ASAP7_75t_L g1071 ( .A(n_173), .Y(n_1071) );
INVx1_ASAP7_75t_L g1111 ( .A(n_174), .Y(n_1111) );
INVx1_ASAP7_75t_L g581 ( .A(n_176), .Y(n_581) );
INVx2_ASAP7_75t_L g1542 ( .A(n_177), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_177), .B(n_1543), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_177), .B(n_302), .Y(n_1550) );
AOI22xp5_ASAP7_75t_L g1538 ( .A1(n_178), .A2(n_271), .B1(n_1539), .B2(n_1544), .Y(n_1538) );
INVx1_ASAP7_75t_L g1082 ( .A(n_180), .Y(n_1082) );
INVx1_ASAP7_75t_L g1507 ( .A(n_181), .Y(n_1507) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_182), .Y(n_867) );
INVx1_ASAP7_75t_L g1054 ( .A(n_183), .Y(n_1054) );
INVx1_ASAP7_75t_L g1280 ( .A(n_184), .Y(n_1280) );
INVx1_ASAP7_75t_L g759 ( .A(n_185), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_187), .A2(n_278), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g1360 ( .A(n_188), .Y(n_1360) );
AOI22xp5_ASAP7_75t_L g1560 ( .A1(n_189), .A2(n_309), .B1(n_1547), .B2(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g920 ( .A(n_190), .Y(n_920) );
XOR2xp5_ASAP7_75t_L g955 ( .A(n_191), .B(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g1236 ( .A(n_192), .Y(n_1236) );
OAI22xp33_ASAP7_75t_L g1247 ( .A1(n_192), .A2(n_223), .B1(n_482), .B2(n_752), .Y(n_1247) );
XNOR2x2_ASAP7_75t_L g631 ( .A(n_193), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g961 ( .A(n_194), .Y(n_961) );
INVx1_ASAP7_75t_L g565 ( .A(n_195), .Y(n_565) );
INVx1_ASAP7_75t_L g1028 ( .A(n_196), .Y(n_1028) );
INVx1_ASAP7_75t_L g1365 ( .A(n_197), .Y(n_1365) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_198), .A2(n_254), .B1(n_535), .B2(n_1425), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_198), .A2(n_291), .B1(n_431), .B2(n_1022), .Y(n_1435) );
OAI211xp5_ASAP7_75t_L g898 ( .A1(n_201), .A2(n_899), .B(n_900), .C(n_909), .Y(n_898) );
INVx1_ASAP7_75t_L g941 ( .A(n_201), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g1755 ( .A(n_202), .Y(n_1755) );
INVx1_ASAP7_75t_L g1119 ( .A(n_203), .Y(n_1119) );
INVx1_ASAP7_75t_L g964 ( .A(n_204), .Y(n_964) );
OAI22xp33_ASAP7_75t_L g1158 ( .A1(n_205), .A2(n_292), .B1(n_378), .B2(n_752), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g1171 ( .A1(n_205), .A2(n_292), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
INVx2_ASAP7_75t_L g423 ( .A(n_206), .Y(n_423) );
INVx1_ASAP7_75t_L g440 ( .A(n_206), .Y(n_440) );
INVx1_ASAP7_75t_L g1465 ( .A(n_207), .Y(n_1465) );
XNOR2xp5_ASAP7_75t_L g1056 ( .A(n_209), .B(n_1057), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_210), .A2(n_277), .B1(n_492), .B2(n_493), .Y(n_554) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_210), .A2(n_237), .B1(n_444), .B2(n_446), .Y(n_570) );
INVx1_ASAP7_75t_L g1213 ( .A(n_212), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_213), .A2(n_311), .B1(n_1539), .B2(n_1544), .Y(n_1564) );
INVx1_ASAP7_75t_L g908 ( .A(n_214), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_214), .A2(n_242), .B1(n_446), .B2(n_467), .Y(n_938) );
INVx1_ASAP7_75t_L g901 ( .A(n_215), .Y(n_901) );
INVx1_ASAP7_75t_L g1230 ( .A(n_216), .Y(n_1230) );
OA211x2_ASAP7_75t_L g1243 ( .A1(n_216), .A2(n_556), .B(n_1244), .C(n_1245), .Y(n_1243) );
BUFx3_ASAP7_75t_L g403 ( .A(n_217), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_219), .A2(n_349), .B1(n_378), .B2(n_752), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_219), .A2(n_349), .B1(n_731), .B2(n_1034), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g1779 ( .A(n_220), .Y(n_1779) );
OAI22xp5_ASAP7_75t_SL g1197 ( .A1(n_221), .A2(n_1198), .B1(n_1240), .B2(n_1249), .Y(n_1197) );
NAND4xp25_ASAP7_75t_L g1198 ( .A(n_221), .B(n_1199), .C(n_1215), .D(n_1224), .Y(n_1198) );
XOR2xp5_ASAP7_75t_L g1106 ( .A(n_222), .B(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1233 ( .A(n_223), .Y(n_1233) );
INVx1_ASAP7_75t_L g1029 ( .A(n_224), .Y(n_1029) );
OAI211xp5_ASAP7_75t_L g1036 ( .A1(n_224), .A2(n_713), .B(n_1037), .C(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g1311 ( .A(n_225), .Y(n_1311) );
INVx1_ASAP7_75t_L g1756 ( .A(n_226), .Y(n_1756) );
OAI211xp5_ASAP7_75t_L g1761 ( .A1(n_226), .A2(n_453), .B(n_1762), .C(n_1764), .Y(n_1761) );
INVx1_ASAP7_75t_L g913 ( .A(n_228), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_228), .B(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g1401 ( .A(n_229), .Y(n_1401) );
INVx1_ASAP7_75t_L g1114 ( .A(n_230), .Y(n_1114) );
INVx1_ASAP7_75t_L g1206 ( .A(n_231), .Y(n_1206) );
OAI22xp33_ASAP7_75t_L g1262 ( .A1(n_232), .A2(n_321), .B1(n_378), .B2(n_752), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1270 ( .A1(n_232), .A2(n_321), .B1(n_707), .B2(n_731), .Y(n_1270) );
INVx1_ASAP7_75t_L g1181 ( .A(n_233), .Y(n_1181) );
INVx1_ASAP7_75t_L g1364 ( .A(n_234), .Y(n_1364) );
AOI22xp5_ASAP7_75t_L g1556 ( .A1(n_235), .A2(n_261), .B1(n_1547), .B2(n_1549), .Y(n_1556) );
INVx1_ASAP7_75t_L g562 ( .A(n_236), .Y(n_562) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_237), .A2(n_280), .B1(n_482), .B2(n_568), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g1776 ( .A(n_238), .Y(n_1776) );
INVx1_ASAP7_75t_L g1314 ( .A(n_239), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_239), .A2(n_303), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
XOR2xp5_ASAP7_75t_L g855 ( .A(n_240), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g1278 ( .A(n_241), .Y(n_1278) );
INVx1_ASAP7_75t_L g910 ( .A(n_242), .Y(n_910) );
BUFx3_ASAP7_75t_L g386 ( .A(n_243), .Y(n_386) );
INVx1_ASAP7_75t_L g487 ( .A(n_243), .Y(n_487) );
INVx1_ASAP7_75t_L g692 ( .A(n_244), .Y(n_692) );
XOR2x2_ASAP7_75t_L g727 ( .A(n_246), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g960 ( .A(n_248), .Y(n_960) );
INVx1_ASAP7_75t_L g1229 ( .A(n_249), .Y(n_1229) );
INVx1_ASAP7_75t_L g1214 ( .A(n_250), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_251), .A2(n_301), .B1(n_1014), .B2(n_1384), .Y(n_1383) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_252), .A2(n_284), .B1(n_399), .B2(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g1449 ( .A(n_253), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_255), .A2(n_351), .B1(n_1386), .B2(n_1388), .Y(n_1385) );
XNOR2x1_ASAP7_75t_L g1004 ( .A(n_256), .B(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g660 ( .A(n_257), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_258), .A2(n_332), .B1(n_946), .B2(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1012 ( .A(n_259), .Y(n_1012) );
OAI211xp5_ASAP7_75t_L g1060 ( .A1(n_260), .A2(n_696), .B(n_1061), .C(n_1062), .Y(n_1060) );
INVx1_ASAP7_75t_L g1101 ( .A(n_260), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_263), .A2(n_353), .B1(n_983), .B2(n_1014), .Y(n_1013) );
INVxp33_ASAP7_75t_SL g1049 ( .A(n_263), .Y(n_1049) );
OAI211xp5_ASAP7_75t_L g555 ( .A1(n_264), .A2(n_556), .B(n_560), .C(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g575 ( .A(n_264), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_265), .Y(n_807) );
INVx1_ASAP7_75t_L g1509 ( .A(n_266), .Y(n_1509) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_268), .B(n_446), .Y(n_888) );
INVx1_ASAP7_75t_L g1464 ( .A(n_269), .Y(n_1464) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_270), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_272), .Y(n_812) );
INVx1_ASAP7_75t_L g1450 ( .A(n_273), .Y(n_1450) );
OAI211xp5_ASAP7_75t_L g1454 ( .A1(n_273), .A2(n_598), .B(n_1244), .C(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1400 ( .A(n_274), .Y(n_1400) );
INVx1_ASAP7_75t_L g1210 ( .A(n_275), .Y(n_1210) );
XOR2x2_ASAP7_75t_L g1155 ( .A(n_276), .B(n_1156), .Y(n_1155) );
OAI22xp33_ASAP7_75t_L g576 ( .A1(n_277), .A2(n_280), .B1(n_465), .B2(n_467), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_278), .A2(n_322), .B1(n_465), .B2(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g402 ( .A(n_279), .Y(n_402) );
INVx1_ASAP7_75t_L g410 ( .A(n_279), .Y(n_410) );
INVx1_ASAP7_75t_L g659 ( .A(n_281), .Y(n_659) );
INVx1_ASAP7_75t_L g643 ( .A(n_282), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_283), .A2(n_340), .B1(n_747), .B2(n_1031), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_283), .A2(n_340), .B1(n_1042), .B2(n_1044), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_284), .A2(n_325), .B1(n_535), .B2(n_537), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_285), .A2(n_342), .B1(n_699), .B2(n_701), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_285), .A2(n_342), .B1(n_721), .B2(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g1207 ( .A(n_286), .Y(n_1207) );
INVx1_ASAP7_75t_L g1469 ( .A(n_287), .Y(n_1469) );
INVx1_ASAP7_75t_L g1018 ( .A(n_288), .Y(n_1018) );
INVx1_ASAP7_75t_L g1500 ( .A(n_289), .Y(n_1500) );
INVx1_ASAP7_75t_L g1312 ( .A(n_293), .Y(n_1312) );
INVx1_ASAP7_75t_L g833 ( .A(n_294), .Y(n_833) );
OAI211xp5_ASAP7_75t_SL g844 ( .A1(n_294), .A2(n_713), .B(n_845), .C(n_847), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g1758 ( .A1(n_296), .A2(n_298), .B1(n_378), .B2(n_752), .Y(n_1758) );
OAI22xp33_ASAP7_75t_L g1766 ( .A1(n_296), .A2(n_298), .B1(n_731), .B2(n_1172), .Y(n_1766) );
INVx1_ASAP7_75t_L g765 ( .A(n_297), .Y(n_765) );
INVx1_ASAP7_75t_L g963 ( .A(n_299), .Y(n_963) );
INVx1_ASAP7_75t_L g1468 ( .A(n_300), .Y(n_1468) );
AOI22xp33_ASAP7_75t_SL g1379 ( .A1(n_301), .A2(n_339), .B1(n_902), .B2(n_1377), .Y(n_1379) );
INVx1_ASAP7_75t_L g1543 ( .A(n_302), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_302), .B(n_1542), .Y(n_1548) );
INVx1_ASAP7_75t_L g1301 ( .A(n_303), .Y(n_1301) );
INVx1_ASAP7_75t_L g1408 ( .A(n_304), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_306), .A2(n_346), .B1(n_446), .B2(n_467), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g1770 ( .A(n_307), .Y(n_1770) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_308), .A2(n_347), .B1(n_1539), .B2(n_1544), .Y(n_1571) );
INVx1_ASAP7_75t_L g1318 ( .A(n_310), .Y(n_1318) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_312), .Y(n_922) );
OAI211xp5_ASAP7_75t_SL g882 ( .A1(n_313), .A2(n_560), .B(n_831), .C(n_883), .Y(n_882) );
OAI211xp5_ASAP7_75t_SL g890 ( .A1(n_313), .A2(n_713), .B(n_891), .C(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g587 ( .A(n_314), .Y(n_587) );
INVx1_ASAP7_75t_L g985 ( .A(n_315), .Y(n_985) );
INVx1_ASAP7_75t_L g1019 ( .A(n_316), .Y(n_1019) );
INVx1_ASAP7_75t_L g1080 ( .A(n_317), .Y(n_1080) );
XOR2x2_ASAP7_75t_L g551 ( .A(n_318), .B(n_552), .Y(n_551) );
OAI211xp5_ASAP7_75t_L g1753 ( .A1(n_320), .A2(n_741), .B(n_1244), .C(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1765 ( .A(n_320), .Y(n_1765) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_322), .Y(n_484) );
INVx1_ASAP7_75t_L g1501 ( .A(n_323), .Y(n_1501) );
INVx1_ASAP7_75t_L g1143 ( .A(n_324), .Y(n_1143) );
OAI211xp5_ASAP7_75t_L g1150 ( .A1(n_324), .A2(n_453), .B(n_1037), .C(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g432 ( .A(n_325), .Y(n_432) );
INVx1_ASAP7_75t_L g1070 ( .A(n_326), .Y(n_1070) );
OAI211xp5_ASAP7_75t_SL g1257 ( .A1(n_327), .A2(n_687), .B(n_1244), .C(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1269 ( .A(n_327), .Y(n_1269) );
INVx1_ASAP7_75t_L g1275 ( .A(n_328), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_329), .Y(n_815) );
INVx1_ASAP7_75t_L g1359 ( .A(n_330), .Y(n_1359) );
CKINVDCx5p33_ASAP7_75t_R g1772 ( .A(n_331), .Y(n_1772) );
INVx1_ASAP7_75t_L g1202 ( .A(n_333), .Y(n_1202) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
INVx1_ASAP7_75t_L g1184 ( .A(n_335), .Y(n_1184) );
INVx1_ASAP7_75t_L g1124 ( .A(n_336), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g1775 ( .A(n_337), .Y(n_1775) );
OA22x2_ASAP7_75t_L g1355 ( .A1(n_338), .A2(n_1356), .B1(n_1394), .B2(n_1395), .Y(n_1355) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_338), .Y(n_1395) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_343), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_344), .Y(n_864) );
XOR2x2_ASAP7_75t_L g1750 ( .A(n_347), .B(n_1751), .Y(n_1750) );
AOI22xp5_ASAP7_75t_L g1796 ( .A1(n_347), .A2(n_1797), .B1(n_1800), .B2(n_1803), .Y(n_1796) );
INVx2_ASAP7_75t_L g427 ( .A(n_348), .Y(n_427) );
INVx1_ASAP7_75t_L g477 ( .A(n_348), .Y(n_477) );
INVx1_ASAP7_75t_L g679 ( .A(n_348), .Y(n_679) );
INVx1_ASAP7_75t_L g1074 ( .A(n_350), .Y(n_1074) );
INVx1_ASAP7_75t_L g1237 ( .A(n_352), .Y(n_1237) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_353), .Y(n_1053) );
INVx1_ASAP7_75t_L g1409 ( .A(n_354), .Y(n_1409) );
INVx1_ASAP7_75t_L g1185 ( .A(n_355), .Y(n_1185) );
AOI21xp33_ASAP7_75t_L g924 ( .A1(n_356), .A2(n_535), .B(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g944 ( .A(n_356), .Y(n_944) );
INVx1_ASAP7_75t_L g773 ( .A(n_357), .Y(n_773) );
INVx1_ASAP7_75t_L g1231 ( .A(n_358), .Y(n_1231) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_359), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_387), .B(n_1530), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx4f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_372), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g1795 ( .A(n_366), .B(n_375), .Y(n_1795) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g1802 ( .A(n_368), .B(n_371), .Y(n_1802) );
INVx1_ASAP7_75t_L g1805 ( .A(n_368), .Y(n_1805) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g1808 ( .A(n_371), .B(n_1805), .Y(n_1808) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g514 ( .A(n_375), .B(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_SL g897 ( .A1(n_375), .A2(n_898), .B(n_911), .Y(n_897) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g541 ( .A(n_376), .B(n_386), .Y(n_541) );
AND2x4_ASAP7_75t_L g926 ( .A(n_376), .B(n_385), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_377), .A2(n_485), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
AOI22xp5_ASAP7_75t_L g1358 ( .A1(n_377), .A2(n_485), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AOI22xp33_ASAP7_75t_SL g1508 ( .A1(n_377), .A2(n_485), .B1(n_1509), .B2(n_1510), .Y(n_1508) );
AND2x4_ASAP7_75t_SL g1794 ( .A(n_377), .B(n_1795), .Y(n_1794) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
OR2x2_ASAP7_75t_L g492 ( .A(n_379), .B(n_486), .Y(n_492) );
OR2x6_ASAP7_75t_L g700 ( .A(n_379), .B(n_486), .Y(n_700) );
INVx1_ASAP7_75t_L g827 ( .A(n_379), .Y(n_827) );
BUFx4f_ASAP7_75t_L g914 ( .A(n_379), .Y(n_914) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g483 ( .A(n_380), .Y(n_483) );
BUFx4f_ASAP7_75t_L g583 ( .A(n_380), .Y(n_583) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g488 ( .A(n_382), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g497 ( .A(n_382), .Y(n_497) );
INVx1_ASAP7_75t_L g504 ( .A(n_382), .Y(n_504) );
AND2x2_ASAP7_75t_L g510 ( .A(n_382), .B(n_383), .Y(n_510) );
INVx2_ASAP7_75t_L g530 ( .A(n_382), .Y(n_530) );
NAND2x1_ASAP7_75t_L g559 ( .A(n_382), .B(n_383), .Y(n_559) );
INVx2_ASAP7_75t_L g489 ( .A(n_383), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_383), .B(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g501 ( .A(n_383), .Y(n_501) );
INVx1_ASAP7_75t_L g531 ( .A(n_383), .Y(n_531) );
AND2x2_ASAP7_75t_L g533 ( .A(n_383), .B(n_497), .Y(n_533) );
OR2x2_ASAP7_75t_L g592 ( .A(n_383), .B(n_530), .Y(n_592) );
OR2x6_ASAP7_75t_L g482 ( .A(n_384), .B(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_384), .A2(n_906), .B1(n_907), .B2(n_908), .Y(n_905) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g494 ( .A(n_385), .Y(n_494) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g502 ( .A(n_386), .B(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g564 ( .A(n_386), .Y(n_564) );
XNOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_1000), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
XOR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_790), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_629), .B2(n_789), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
XNOR2x1_ASAP7_75t_L g394 ( .A(n_395), .B(n_551), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_517), .Y(n_395) );
INVx1_ASAP7_75t_L g519 ( .A(n_397), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_411), .B(n_428), .Y(n_397) );
AOI222xp33_ASAP7_75t_L g1228 ( .A1(n_399), .A2(n_457), .B1(n_718), .B2(n_1229), .C1(n_1230), .C2(n_1231), .Y(n_1228) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g431 ( .A(n_400), .Y(n_431) );
INVx2_ASAP7_75t_L g452 ( .A(n_400), .Y(n_452) );
AND2x4_ASAP7_75t_L g454 ( .A(n_400), .B(n_441), .Y(n_454) );
BUFx2_ASAP7_75t_L g573 ( .A(n_400), .Y(n_573) );
BUFx2_ASAP7_75t_L g948 ( .A(n_400), .Y(n_948) );
BUFx2_ASAP7_75t_L g983 ( .A(n_400), .Y(n_983) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_400), .Y(n_1404) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g463 ( .A(n_402), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_402), .B(n_403), .Y(n_469) );
INVx2_ASAP7_75t_L g407 ( .A(n_403), .Y(n_407) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
OR2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_409), .Y(n_445) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx8_ASAP7_75t_L g1022 ( .A(n_405), .Y(n_1022) );
INVx3_ASAP7_75t_L g1523 ( .A(n_405), .Y(n_1523) );
INVx8_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_406), .Y(n_1015) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
AND2x4_ASAP7_75t_L g414 ( .A(n_407), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g415 ( .A(n_410), .Y(n_415) );
INVx1_ASAP7_75t_L g1290 ( .A(n_412), .Y(n_1290) );
INVx1_ASAP7_75t_L g1789 ( .A(n_412), .Y(n_1789) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g466 ( .A(n_413), .B(n_447), .Y(n_466) );
INVx2_ASAP7_75t_L g621 ( .A(n_413), .Y(n_621) );
AND2x4_ASAP7_75t_L g710 ( .A(n_413), .B(n_447), .Y(n_710) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_413), .Y(n_946) );
INVx2_ASAP7_75t_L g1387 ( .A(n_413), .Y(n_1387) );
INVx1_ASAP7_75t_L g1391 ( .A(n_413), .Y(n_1391) );
INVx2_ASAP7_75t_L g1791 ( .A(n_413), .Y(n_1791) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_414), .Y(n_616) );
BUFx8_ASAP7_75t_L g804 ( .A(n_414), .Y(n_804) );
INVx2_ASAP7_75t_L g953 ( .A(n_414), .Y(n_953) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_R g1388 ( .A(n_417), .Y(n_1388) );
INVx5_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g950 ( .A(n_418), .Y(n_950) );
BUFx12f_ASAP7_75t_L g1434 ( .A(n_418), .Y(n_1434) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
BUFx2_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_419), .B(n_463), .Y(n_613) );
INVx2_ASAP7_75t_L g851 ( .A(n_419), .Y(n_851) );
INVx1_ASAP7_75t_L g849 ( .A(n_420), .Y(n_849) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI33xp33_ASAP7_75t_L g1382 ( .A1(n_422), .A2(n_1383), .A3(n_1385), .B1(n_1389), .B2(n_1392), .B3(n_1393), .Y(n_1382) );
NAND3xp33_ASAP7_75t_L g1432 ( .A(n_422), .B(n_1433), .C(n_1435), .Y(n_1432) );
AND3x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .C(n_426), .Y(n_422) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_423), .Y(n_472) );
NAND2xp33_ASAP7_75t_SL g608 ( .A(n_423), .B(n_425), .Y(n_608) );
INVx3_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
AND2x2_ASAP7_75t_L g848 ( .A(n_424), .B(n_849), .Y(n_848) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g441 ( .A(n_425), .Y(n_441) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g438 ( .A(n_427), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_433), .B2(n_435), .C(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI211xp5_ASAP7_75t_L g1343 ( .A1(n_431), .A2(n_454), .B(n_1344), .C(n_1345), .Y(n_1343) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI33xp33_ASAP7_75t_L g958 ( .A1(n_437), .A2(n_755), .A3(n_959), .B1(n_962), .B2(n_965), .B3(n_970), .Y(n_958) );
OAI33xp33_ASAP7_75t_L g1200 ( .A1(n_437), .A2(n_755), .A3(n_1201), .B1(n_1204), .B2(n_1208), .B3(n_1212), .Y(n_1200) );
INVx1_ASAP7_75t_L g1393 ( .A(n_437), .Y(n_1393) );
OAI33xp33_ASAP7_75t_L g1462 ( .A1(n_437), .A2(n_755), .A3(n_1463), .B1(n_1467), .B2(n_1470), .B3(n_1473), .Y(n_1462) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
AND2x4_ASAP7_75t_L g524 ( .A(n_438), .B(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g623 ( .A(n_438), .B(n_439), .Y(n_623) );
INVx1_ASAP7_75t_L g930 ( .A(n_438), .Y(n_930) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND3x1_ASAP7_75t_L g677 ( .A(n_440), .B(n_441), .C(n_678), .Y(n_677) );
OR2x4_ASAP7_75t_L g444 ( .A(n_441), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_441), .Y(n_447) );
OR2x6_ASAP7_75t_L g467 ( .A(n_441), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_442), .B(n_478), .Y(n_518) );
OAI31xp33_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_448), .A3(n_464), .B(n_470), .Y(n_442) );
INVx2_ASAP7_75t_SL g708 ( .A(n_444), .Y(n_708) );
INVx1_ASAP7_75t_L g940 ( .A(n_444), .Y(n_940) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_444), .Y(n_1035) );
INVx1_ASAP7_75t_L g1149 ( .A(n_444), .Y(n_1149) );
OR2x4_ASAP7_75t_L g446 ( .A(n_445), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g611 ( .A(n_445), .Y(n_611) );
BUFx4f_ASAP7_75t_L g625 ( .A(n_445), .Y(n_625) );
BUFx3_ASAP7_75t_L g666 ( .A(n_445), .Y(n_666) );
BUFx3_ASAP7_75t_L g758 ( .A(n_445), .Y(n_758) );
BUFx3_ASAP7_75t_L g721 ( .A(n_446), .Y(n_721) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_446), .Y(n_1045) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_446), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1518 ( .A(n_446), .Y(n_1518) );
NAND3xp33_ASAP7_75t_SL g448 ( .A(n_449), .B(n_453), .C(n_455), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_450), .A2(n_456), .B1(n_500), .B2(n_502), .Y(n_499) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g1384 ( .A(n_452), .Y(n_1384) );
INVx2_ASAP7_75t_L g1513 ( .A(n_452), .Y(n_1513) );
NAND3xp33_ASAP7_75t_SL g571 ( .A(n_453), .B(n_572), .C(n_574), .Y(n_571) );
CKINVDCx8_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
CKINVDCx8_ASAP7_75t_R g713 ( .A(n_454), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g933 ( .A(n_454), .B(n_934), .C(n_938), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g1226 ( .A(n_454), .B(n_1227), .Y(n_1226) );
NOR3xp33_ASAP7_75t_L g1368 ( .A(n_454), .B(n_1369), .C(n_1370), .Y(n_1368) );
AOI211xp5_ASAP7_75t_L g1402 ( .A1(n_454), .A2(n_1403), .B(n_1404), .C(n_1405), .Y(n_1402) );
AOI211xp5_ASAP7_75t_L g1512 ( .A1(n_454), .A2(n_1505), .B(n_1513), .C(n_1514), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_460), .B2(n_461), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_457), .A2(n_461), .B1(n_562), .B2(n_575), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_457), .A2(n_848), .B1(n_884), .B2(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g936 ( .A(n_457), .Y(n_936) );
AOI222xp33_ASAP7_75t_L g982 ( .A1(n_457), .A2(n_461), .B1(n_983), .B2(n_984), .C1(n_985), .C2(n_986), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_457), .B(n_1364), .Y(n_1371) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AND2x2_ASAP7_75t_L g461 ( .A(n_458), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g716 ( .A(n_458), .B(n_459), .Y(n_716) );
AND2x4_ASAP7_75t_L g718 ( .A(n_458), .B(n_462), .Y(n_718) );
AND2x4_ASAP7_75t_L g846 ( .A(n_458), .B(n_459), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_460), .B(n_506), .Y(n_505) );
AOI32xp33_ASAP7_75t_L g847 ( .A1(n_461), .A2(n_834), .A3(n_848), .B1(n_850), .B2(n_852), .Y(n_847) );
INVxp67_ASAP7_75t_L g891 ( .A(n_461), .Y(n_891) );
INVxp67_ASAP7_75t_L g937 ( .A(n_461), .Y(n_937) );
INVx1_ASAP7_75t_L g1406 ( .A(n_461), .Y(n_1406) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_466), .A2(n_906), .B1(n_940), .B2(n_941), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_466), .A2(n_723), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g723 ( .A(n_467), .Y(n_723) );
INVx2_ASAP7_75t_L g989 ( .A(n_467), .Y(n_989) );
INVx1_ASAP7_75t_L g1043 ( .A(n_467), .Y(n_1043) );
BUFx3_ASAP7_75t_L g674 ( .A(n_468), .Y(n_674) );
INVx1_ASAP7_75t_L g806 ( .A(n_468), .Y(n_806) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g619 ( .A(n_469), .Y(n_619) );
OAI31xp33_ASAP7_75t_SL g569 ( .A1(n_470), .A2(n_570), .A3(n_571), .B(n_576), .Y(n_569) );
INVx1_ASAP7_75t_L g1373 ( .A(n_470), .Y(n_1373) );
OAI31xp33_ASAP7_75t_L g1445 ( .A1(n_470), .A2(n_1446), .A3(n_1447), .B(n_1451), .Y(n_1445) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_471), .B(n_473), .Y(n_725) );
AND2x2_ASAP7_75t_L g854 ( .A(n_471), .B(n_473), .Y(n_854) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_471), .B(n_473), .Y(n_1154) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_471), .B(n_473), .Y(n_1239) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_475), .B(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g607 ( .A(n_475), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g656 ( .A(n_475), .Y(n_656) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g516 ( .A(n_476), .Y(n_516) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AO21x1_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_490), .B(n_513), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_484), .B2(n_485), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g1412 ( .A(n_482), .Y(n_1412) );
BUFx3_ASAP7_75t_L g658 ( .A(n_483), .Y(n_658) );
BUFx3_ASAP7_75t_L g874 ( .A(n_483), .Y(n_874) );
BUFx6f_ASAP7_75t_L g979 ( .A(n_483), .Y(n_979) );
INVx2_ASAP7_75t_SL g1479 ( .A(n_483), .Y(n_1479) );
INVx4_ASAP7_75t_L g568 ( .A(n_485), .Y(n_568) );
CKINVDCx16_ASAP7_75t_R g752 ( .A(n_485), .Y(n_752) );
INVx3_ASAP7_75t_SL g899 ( .A(n_485), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_485), .A2(n_1400), .B1(n_1401), .B2(n_1412), .Y(n_1411) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
BUFx3_ASAP7_75t_L g1424 ( .A(n_488), .Y(n_1424) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_498), .Y(n_490) );
INVx1_ASAP7_75t_L g998 ( .A(n_493), .Y(n_998) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
AND2x2_ASAP7_75t_L g500 ( .A(n_494), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g512 ( .A(n_494), .B(n_508), .Y(n_512) );
AND2x2_ASAP7_75t_L g697 ( .A(n_494), .B(n_538), .Y(n_697) );
INVx8_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
OR2x2_ASAP7_75t_L g703 ( .A(n_495), .B(n_564), .Y(n_703) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_495), .Y(n_1219) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .C(n_511), .Y(n_498) );
INVx1_ASAP7_75t_L g904 ( .A(n_500), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g1363 ( .A1(n_500), .A2(n_835), .B1(n_1364), .B2(n_1365), .Y(n_1363) );
AOI22xp5_ASAP7_75t_L g1503 ( .A1(n_500), .A2(n_835), .B1(n_1504), .B2(n_1505), .Y(n_1503) );
AND2x4_ASAP7_75t_L g563 ( .A(n_501), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g744 ( .A(n_501), .B(n_564), .Y(n_744) );
BUFx3_ASAP7_75t_L g566 ( .A(n_502), .Y(n_566) );
INVx2_ASAP7_75t_L g694 ( .A(n_502), .Y(n_694) );
INVx2_ASAP7_75t_L g836 ( .A(n_502), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_502), .A2(n_744), .B1(n_1028), .B2(n_1029), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_502), .A2(n_563), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g1415 ( .A(n_509), .Y(n_1415) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_510), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g1502 ( .A(n_511), .B(n_1503), .C(n_1506), .Y(n_1502) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g560 ( .A(n_512), .Y(n_560) );
AOI211xp5_ASAP7_75t_L g1413 ( .A1(n_512), .A2(n_1414), .B(n_1416), .C(n_1417), .Y(n_1413) );
AOI31xp33_ASAP7_75t_SL g1316 ( .A1(n_513), .A2(n_1317), .A3(n_1320), .B(n_1327), .Y(n_1316) );
AO21x1_ASAP7_75t_L g1357 ( .A1(n_513), .A2(n_1358), .B(n_1361), .Y(n_1357) );
AOI21xp33_ASAP7_75t_L g1498 ( .A1(n_513), .A2(n_1499), .B(n_1508), .Y(n_1498) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI31xp33_ASAP7_75t_L g553 ( .A1(n_514), .A2(n_554), .A3(n_555), .B(n_567), .Y(n_553) );
BUFx3_ASAP7_75t_L g704 ( .A(n_514), .Y(n_704) );
BUFx2_ASAP7_75t_L g841 ( .A(n_514), .Y(n_841) );
OAI31xp33_ASAP7_75t_L g880 ( .A1(n_514), .A2(n_881), .A3(n_882), .B(n_886), .Y(n_880) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_514), .A2(n_991), .B(n_999), .Y(n_990) );
BUFx2_ASAP7_75t_SL g1164 ( .A(n_514), .Y(n_1164) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .A3(n_520), .B(n_548), .Y(n_517) );
INVx1_ASAP7_75t_L g550 ( .A(n_521), .Y(n_550) );
AOI33xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_526), .A3(n_534), .B1(n_539), .B2(n_540), .B3(n_542), .Y(n_521) );
INVx1_ASAP7_75t_L g1217 ( .A(n_522), .Y(n_1217) );
AOI33xp33_ASAP7_75t_L g1374 ( .A1(n_522), .A2(n_540), .A3(n_1375), .B1(n_1376), .B2(n_1379), .B3(n_1380), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_522), .Y(n_1428) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
OAI33xp33_ASAP7_75t_L g1272 ( .A1(n_523), .A2(n_653), .A3(n_1273), .B1(n_1276), .B2(n_1279), .B3(n_1282), .Y(n_1272) );
OAI33xp33_ASAP7_75t_L g1476 ( .A1(n_523), .A2(n_600), .A3(n_1477), .B1(n_1480), .B2(n_1481), .B3(n_1482), .Y(n_1476) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
INVx2_ASAP7_75t_L g635 ( .A(n_524), .Y(n_635) );
INVx2_ASAP7_75t_L g817 ( .A(n_524), .Y(n_817) );
INVx1_ASAP7_75t_L g1773 ( .A(n_524), .Y(n_1773) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g928 ( .A(n_528), .Y(n_928) );
INVx2_ASAP7_75t_L g1334 ( .A(n_528), .Y(n_1334) );
INVx1_ASAP7_75t_L g1427 ( .A(n_528), .Y(n_1427) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_529), .Y(n_545) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g547 ( .A(n_533), .Y(n_547) );
BUFx6f_ASAP7_75t_L g1336 ( .A(n_533), .Y(n_1336) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g1378 ( .A(n_536), .Y(n_1378) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g902 ( .A(n_538), .Y(n_902) );
BUFx6f_ASAP7_75t_L g1323 ( .A(n_538), .Y(n_1323) );
BUFx3_ASAP7_75t_L g1425 ( .A(n_538), .Y(n_1425) );
INVx2_ASAP7_75t_L g600 ( .A(n_540), .Y(n_600) );
INVx2_ASAP7_75t_L g828 ( .A(n_540), .Y(n_828) );
AND2x4_ASAP7_75t_L g654 ( .A(n_541), .B(n_655), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_541), .A2(n_780), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g1497 ( .A(n_541), .B(n_655), .Y(n_1497) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g1381 ( .A(n_544), .Y(n_1381) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g996 ( .A(n_545), .B(n_564), .Y(n_996) );
BUFx6f_ASAP7_75t_L g1341 ( .A(n_545), .Y(n_1341) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g1490 ( .A(n_547), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND3xp33_ASAP7_75t_SL g552 ( .A(n_553), .B(n_569), .C(n_577), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_556), .A2(n_647), .B1(n_1074), .B2(n_1077), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_556), .A2(n_1071), .B1(n_1084), .B2(n_1090), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_556), .A2(n_1135), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_556), .A2(n_644), .B1(n_1277), .B2(n_1278), .Y(n_1276) );
INVx5_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_558), .A2(n_643), .B1(n_644), .B2(n_645), .Y(n_642) );
BUFx2_ASAP7_75t_SL g651 ( .A(n_558), .Y(n_651) );
BUFx3_ASAP7_75t_L g741 ( .A(n_558), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_558), .A2(n_647), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_559), .Y(n_594) );
NAND3xp33_ASAP7_75t_SL g991 ( .A(n_560), .B(n_992), .C(n_994), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_565), .B2(n_566), .Y(n_561) );
BUFx3_ASAP7_75t_L g691 ( .A(n_563), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_563), .A2(n_566), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_563), .A2(n_835), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_563), .A2(n_693), .B1(n_1229), .B2(n_1231), .Y(n_1245) );
INVx1_ASAP7_75t_L g1326 ( .A(n_563), .Y(n_1326) );
O2A1O1Ixp33_ASAP7_75t_L g900 ( .A1(n_564), .A2(n_901), .B(n_902), .C(n_903), .Y(n_900) );
INVx1_ASAP7_75t_L g907 ( .A(n_564), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_565), .B(n_573), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g992 ( .A1(n_566), .A2(n_744), .B1(n_902), .B2(n_985), .C1(n_986), .C2(n_993), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_566), .A2(n_691), .B1(n_1259), .B2(n_1260), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_605), .Y(n_577) );
OAI33xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .A3(n_588), .B1(n_596), .B2(n_600), .B3(n_601), .Y(n_578) );
OAI33xp33_ASAP7_75t_L g872 ( .A1(n_579), .A2(n_828), .A3(n_873), .B1(n_875), .B2(n_876), .B3(n_879), .Y(n_872) );
BUFx6f_ASAP7_75t_L g1047 ( .A(n_579), .Y(n_1047) );
OAI33xp33_ASAP7_75t_L g1085 ( .A1(n_579), .A2(n_653), .A3(n_1086), .B1(n_1088), .B2(n_1089), .B3(n_1092), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_584), .B2(n_587), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_581), .A2(n_597), .B1(n_610), .B2(n_612), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_582), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_582), .A2(n_798), .B1(n_814), .B2(n_819), .Y(n_818) );
INVx4_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g638 ( .A(n_583), .Y(n_638) );
BUFx6f_ASAP7_75t_L g1094 ( .A(n_583), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_584), .A2(n_860), .B1(n_870), .B2(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_584), .A2(n_964), .B1(n_969), .B2(n_979), .Y(n_978) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_SL g603 ( .A(n_586), .Y(n_603) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_586), .Y(n_641) );
INVx4_ASAP7_75t_L g819 ( .A(n_586), .Y(n_819) );
INVx1_ASAP7_75t_L g1087 ( .A(n_586), .Y(n_1087) );
INVx1_ASAP7_75t_L g1096 ( .A(n_586), .Y(n_1096) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_587), .A2(n_599), .B1(n_625), .B2(n_626), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_593), .B2(n_595), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_589), .A2(n_602), .B1(n_615), .B2(n_617), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_590), .A2(n_597), .B1(n_598), .B2(n_599), .Y(n_596) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g644 ( .A(n_591), .Y(n_644) );
BUFx2_ASAP7_75t_L g781 ( .A(n_591), .Y(n_781) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g649 ( .A(n_592), .Y(n_649) );
INVx1_ASAP7_75t_L g822 ( .A(n_592), .Y(n_822) );
BUFx3_ASAP7_75t_L g877 ( .A(n_592), .Y(n_877) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_592), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_593), .A2(n_961), .B1(n_972), .B2(n_977), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g1491 ( .A1(n_593), .A2(n_647), .B1(n_1492), .B2(n_1493), .C(n_1494), .Y(n_1491) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx4f_ASAP7_75t_L g598 ( .A(n_594), .Y(n_598) );
BUFx4f_ASAP7_75t_L g689 ( .A(n_594), .Y(n_689) );
INVx4_ASAP7_75t_L g783 ( .A(n_594), .Y(n_783) );
BUFx4f_ASAP7_75t_L g831 ( .A(n_594), .Y(n_831) );
BUFx4f_ASAP7_75t_L g923 ( .A(n_594), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_595), .A2(n_604), .B1(n_621), .B2(n_622), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_598), .A2(n_821), .B1(n_864), .B2(n_867), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g1486 ( .A1(n_598), .A2(n_977), .B1(n_1487), .B2(n_1488), .C(n_1489), .Y(n_1486) );
OAI33xp33_ASAP7_75t_L g1216 ( .A1(n_600), .A2(n_1217), .A3(n_1218), .B1(n_1220), .B2(n_1222), .B3(n_1223), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_603), .A2(n_914), .B1(n_1207), .B2(n_1211), .Y(n_1223) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_603), .A2(n_1469), .B1(n_1472), .B2(n_1478), .Y(n_1482) );
OAI33xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .A3(n_614), .B1(n_620), .B2(n_623), .B3(n_624), .Y(n_605) );
OAI33xp33_ASAP7_75t_L g796 ( .A1(n_606), .A2(n_623), .A3(n_797), .B1(n_801), .B2(n_808), .B3(n_813), .Y(n_796) );
OAI33xp33_ASAP7_75t_L g858 ( .A1(n_606), .A2(n_623), .A3(n_859), .B1(n_863), .B2(n_866), .B3(n_869), .Y(n_858) );
BUFx3_ASAP7_75t_L g1016 ( .A(n_606), .Y(n_1016) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_606), .A2(n_675), .A3(n_1069), .B1(n_1073), .B2(n_1076), .B3(n_1081), .Y(n_1068) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx4f_ASAP7_75t_L g662 ( .A(n_607), .Y(n_662) );
BUFx2_ASAP7_75t_L g755 ( .A(n_607), .Y(n_755) );
BUFx8_ASAP7_75t_L g1286 ( .A(n_607), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1303 ( .A(n_610), .Y(n_1303) );
OAI22xp33_ASAP7_75t_L g1313 ( .A1(n_610), .A2(n_1083), .B1(n_1314), .B2(n_1315), .Y(n_1313) );
INVx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g1113 ( .A(n_611), .Y(n_1113) );
INVx2_ASAP7_75t_L g668 ( .A(n_612), .Y(n_668) );
OAI22xp33_ASAP7_75t_L g813 ( .A1(n_612), .A2(n_625), .B1(n_814), .B2(n_815), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_612), .A2(n_625), .B1(n_870), .B2(n_871), .Y(n_869) );
BUFx6f_ASAP7_75t_L g1083 ( .A(n_612), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1288 ( .A(n_612), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1473 ( .A1(n_612), .A2(n_1113), .B1(n_1474), .B2(n_1475), .Y(n_1473) );
BUFx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_613), .Y(n_628) );
BUFx2_ASAP7_75t_L g683 ( .A(n_613), .Y(n_683) );
INVx2_ASAP7_75t_L g768 ( .A(n_615), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_615), .A2(n_809), .B1(n_810), .B2(n_812), .Y(n_808) );
OAI22xp33_ASAP7_75t_SL g1117 ( .A1(n_615), .A2(n_1118), .B1(n_1119), .B2(n_1120), .Y(n_1117) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx5_ASAP7_75t_L g670 ( .A(n_616), .Y(n_670) );
INVx2_ASAP7_75t_SL g673 ( .A(n_616), .Y(n_673) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_616), .Y(n_1307) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_617), .A2(n_621), .B1(n_864), .B2(n_865), .Y(n_863) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g622 ( .A(n_618), .Y(n_622) );
CKINVDCx8_ASAP7_75t_R g671 ( .A(n_618), .Y(n_671) );
INVx3_ASAP7_75t_L g968 ( .A(n_618), .Y(n_968) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g811 ( .A(n_619), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_621), .A2(n_674), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1291 ( .A1(n_621), .A2(n_674), .B1(n_1278), .B2(n_1284), .Y(n_1291) );
OAI221xp5_ASAP7_75t_L g1524 ( .A1(n_621), .A2(n_622), .B1(n_1488), .B2(n_1525), .C(n_1526), .Y(n_1524) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_622), .A2(n_673), .B1(n_867), .B2(n_868), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_625), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_625), .A2(n_860), .B1(n_861), .B2(n_862), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g959 ( .A1(n_625), .A2(n_935), .B1(n_960), .B2(n_961), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_625), .A2(n_800), .B1(n_971), .B2(n_972), .Y(n_970) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g712 ( .A(n_627), .Y(n_712) );
INVx2_ASAP7_75t_L g935 ( .A(n_627), .Y(n_935) );
INVx1_ASAP7_75t_L g1037 ( .A(n_627), .Y(n_1037) );
INVx1_ASAP7_75t_L g1072 ( .A(n_627), .Y(n_1072) );
INVx4_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g761 ( .A(n_628), .Y(n_761) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_628), .Y(n_800) );
OA21x2_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_726), .B(n_788), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g789 ( .A1(n_630), .A2(n_726), .B(n_788), .Y(n_789) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g788 ( .A(n_631), .B(n_727), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_684), .C(n_705), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_661), .Y(n_633) );
OAI33xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .A3(n_642), .B1(n_646), .B2(n_653), .B3(n_657), .Y(n_634) );
OAI33xp33_ASAP7_75t_L g775 ( .A1(n_635), .A2(n_776), .A3(n_779), .B1(n_784), .B2(n_786), .B3(n_787), .Y(n_775) );
OAI22xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_637), .A2(n_650), .B1(n_664), .B2(n_667), .Y(n_663) );
INVx2_ASAP7_75t_SL g778 ( .A(n_638), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_639), .A2(n_652), .B1(n_664), .B2(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_640), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_640), .A2(n_757), .B1(n_773), .B2(n_777), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_640), .A2(n_765), .B1(n_770), .B2(n_777), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_640), .A2(n_658), .B1(n_1012), .B2(n_1019), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_640), .A2(n_658), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
OAI22xp33_ASAP7_75t_L g1769 ( .A1(n_640), .A2(n_1770), .B1(n_1771), .B2(n_1772), .Y(n_1769) );
OAI22xp33_ASAP7_75t_L g1780 ( .A1(n_640), .A2(n_1771), .B1(n_1781), .B2(n_1782), .Y(n_1780) );
INVx6_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx5_ASAP7_75t_L g916 ( .A(n_641), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_643), .A2(n_659), .B1(n_670), .B2(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g1091 ( .A(n_644), .Y(n_1091) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_644), .A2(n_741), .B1(n_1306), .B2(n_1311), .C(n_1333), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_645), .A2(n_660), .B1(n_673), .B2(n_674), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_647), .A2(n_651), .B1(n_1011), .B2(n_1018), .Y(n_1051) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx4_ASAP7_75t_L g1135 ( .A(n_648), .Y(n_1135) );
INVx4_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI33xp33_ASAP7_75t_L g1132 ( .A1(n_653), .A2(n_1047), .A3(n_1133), .B1(n_1134), .B2(n_1136), .B3(n_1137), .Y(n_1132) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_654), .Y(n_786) );
NAND3xp33_ASAP7_75t_L g1429 ( .A(n_654), .B(n_1430), .C(n_1431), .Y(n_1429) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI33xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .A3(n_669), .B1(n_672), .B2(n_675), .B3(n_680), .Y(n_661) );
OAI33xp33_ASAP7_75t_L g1109 ( .A1(n_662), .A2(n_1110), .A3(n_1117), .B1(n_1122), .B2(n_1126), .B3(n_1129), .Y(n_1109) );
OAI33xp33_ASAP7_75t_L g1189 ( .A1(n_662), .A2(n_771), .A3(n_1190), .B1(n_1191), .B2(n_1192), .B3(n_1193), .Y(n_1189) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_664), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1069) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g1294 ( .A(n_666), .Y(n_1294) );
INVx1_ASAP7_75t_L g1786 ( .A(n_666), .Y(n_1786) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx3_ASAP7_75t_L g764 ( .A(n_670), .Y(n_764) );
INVx8_ASAP7_75t_L g1079 ( .A(n_670), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_670), .A2(n_671), .B1(n_1181), .B2(n_1188), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_671), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g951 ( .A1(n_671), .A2(n_915), .B1(n_922), .B2(n_952), .C(n_954), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_671), .A2(n_1123), .B1(n_1124), .B2(n_1125), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_673), .A2(n_1120), .B1(n_1180), .B2(n_1187), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_674), .A2(n_767), .B1(n_769), .B2(n_770), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_674), .A2(n_1009), .B1(n_1011), .B2(n_1012), .C(n_1013), .Y(n_1008) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_674), .A2(n_945), .B1(n_1018), .B2(n_1019), .C(n_1020), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_674), .A2(n_1077), .B1(n_1078), .B2(n_1080), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_674), .A2(n_1277), .B1(n_1283), .B2(n_1290), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g1520 ( .A1(n_674), .A2(n_1387), .B1(n_1487), .B2(n_1521), .C(n_1522), .Y(n_1520) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_676), .Y(n_771) );
INVx2_ASAP7_75t_L g1023 ( .A(n_676), .Y(n_1023) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g1128 ( .A(n_677), .Y(n_1128) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g772 ( .A1(n_681), .A2(n_758), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_681), .A2(n_1112), .B1(n_1177), .B2(n_1184), .Y(n_1190) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g1116 ( .A(n_683), .Y(n_1116) );
OAI31xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .A3(n_698), .B(n_704), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g1777 ( .A1(n_689), .A2(n_977), .B1(n_1778), .B2(n_1779), .Y(n_1777) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_693), .B2(n_695), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_691), .A2(n_835), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_692), .A2(n_715), .B1(n_717), .B2(n_719), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_693), .A2(n_734), .B1(n_744), .B2(n_745), .Y(n_743) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g1457 ( .A(n_694), .Y(n_1457) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g742 ( .A(n_697), .Y(n_742) );
INVx3_ASAP7_75t_L g1244 ( .A(n_697), .Y(n_1244) );
AOI211xp5_ASAP7_75t_L g1320 ( .A1(n_697), .A2(n_1321), .B(n_1324), .C(n_1325), .Y(n_1320) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g747 ( .A(n_700), .Y(n_747) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g1031 ( .A(n_702), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_702), .A2(n_996), .B1(n_1408), .B2(n_1409), .Y(n_1418) );
INVxp67_ASAP7_75t_SL g1459 ( .A(n_702), .Y(n_1459) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g750 ( .A(n_703), .Y(n_750) );
INVx1_ASAP7_75t_L g839 ( .A(n_703), .Y(n_839) );
OAI31xp33_ASAP7_75t_L g737 ( .A1(n_704), .A2(n_738), .A3(n_746), .B(n_751), .Y(n_737) );
OAI31xp33_ASAP7_75t_L g1058 ( .A1(n_704), .A2(n_1059), .A3(n_1060), .B(n_1065), .Y(n_1058) );
OAI31xp33_ASAP7_75t_SL g1139 ( .A1(n_704), .A2(n_1140), .A3(n_1144), .B(n_1145), .Y(n_1139) );
OAI31xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_711), .A3(n_720), .B(n_724), .Y(n_705) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_708), .A2(n_710), .B1(n_1509), .B2(n_1510), .Y(n_1515) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g731 ( .A(n_710), .Y(n_731) );
INVx1_ASAP7_75t_L g1173 ( .A(n_710), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_710), .A2(n_1035), .B1(n_1318), .B2(n_1319), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_710), .A2(n_1035), .B1(n_1359), .B2(n_1360), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_710), .A2(n_1035), .B1(n_1400), .B2(n_1401), .Y(n_1399) );
INVx2_ASAP7_75t_L g1452 ( .A(n_710), .Y(n_1452) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_712), .A2(n_1112), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_712), .A2(n_1275), .B1(n_1281), .B2(n_1293), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1792 ( .A1(n_712), .A2(n_1293), .B1(n_1772), .B2(n_1779), .Y(n_1792) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_715), .A2(n_717), .B1(n_734), .B2(n_735), .Y(n_733) );
BUFx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_716), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_717), .A2(n_1028), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_717), .A2(n_1039), .B1(n_1063), .B2(n_1101), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g1268 ( .A1(n_717), .A2(n_1039), .B1(n_1259), .B2(n_1269), .Y(n_1268) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g1151 ( .A1(n_718), .A2(n_846), .B1(n_1142), .B2(n_1152), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_718), .A2(n_846), .B1(n_1161), .B2(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1346 ( .A(n_718), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_718), .A2(n_846), .B1(n_1449), .B2(n_1450), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1764 ( .A1(n_718), .A2(n_846), .B1(n_1755), .B2(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI31xp33_ASAP7_75t_L g729 ( .A1(n_724), .A2(n_730), .A3(n_732), .B(n_736), .Y(n_729) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g931 ( .A1(n_725), .A2(n_932), .B(n_942), .Y(n_931) );
OAI31xp33_ASAP7_75t_L g1032 ( .A1(n_725), .A2(n_1033), .A3(n_1036), .B(n_1041), .Y(n_1032) );
OAI31xp33_ASAP7_75t_L g1097 ( .A1(n_725), .A2(n_1098), .A3(n_1099), .B(n_1102), .Y(n_1097) );
OAI31xp33_ASAP7_75t_L g1263 ( .A1(n_725), .A2(n_1264), .A3(n_1267), .B(n_1270), .Y(n_1263) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_725), .A2(n_1164), .B1(n_1398), .B2(n_1410), .C(n_1419), .Y(n_1397) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_737), .C(n_753), .Y(n_728) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g1061 ( .A(n_741), .Y(n_1061) );
OAI221xp5_ASAP7_75t_L g1337 ( .A1(n_741), .A2(n_1304), .B1(n_1315), .B2(n_1338), .C(n_1340), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1480 ( .A1(n_741), .A2(n_1221), .B1(n_1468), .B2(n_1471), .Y(n_1480) );
OAI22xp5_ASAP7_75t_L g1481 ( .A1(n_741), .A2(n_1221), .B1(n_1465), .B2(n_1475), .Y(n_1481) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_744), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_744), .A2(n_1449), .B1(n_1456), .B2(n_1457), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1754 ( .A1(n_744), .A2(n_1457), .B1(n_1755), .B2(n_1756), .Y(n_1754) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_749), .A2(n_996), .B1(n_1500), .B2(n_1501), .C(n_1502), .Y(n_1499) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_750), .Y(n_1066) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_775), .Y(n_753) );
OAI33xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .A3(n_762), .B1(n_766), .B2(n_771), .B3(n_772), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_755), .A2(n_771), .B1(n_943), .B2(n_951), .Y(n_942) );
OAI22xp33_ASAP7_75t_L g1519 ( .A1(n_755), .A2(n_1520), .B1(n_1524), .B2(n_1527), .Y(n_1519) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_758), .A2(n_1082), .B1(n_1083), .B2(n_1084), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1212 ( .A1(n_758), .A2(n_800), .B1(n_1213), .B2(n_1214), .Y(n_1212) );
OAI22xp33_ASAP7_75t_L g1287 ( .A1(n_758), .A2(n_1274), .B1(n_1280), .B2(n_1288), .Y(n_1287) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_759), .A2(n_774), .B1(n_780), .B2(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx3_ASAP7_75t_L g861 ( .A(n_761), .Y(n_861) );
INVx2_ASAP7_75t_L g1787 ( .A(n_761), .Y(n_1787) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_763), .A2(n_769), .B1(n_780), .B2(n_782), .Y(n_779) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI33xp33_ASAP7_75t_L g1285 ( .A1(n_771), .A2(n_1286), .A3(n_1287), .B1(n_1289), .B2(n_1291), .B3(n_1292), .Y(n_1285) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_777), .A2(n_1070), .B1(n_1082), .B2(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_780), .A2(n_831), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_780), .A2(n_918), .B1(n_1203), .B2(n_1214), .Y(n_1222) );
INVx4_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_783), .Y(n_785) );
INVx2_ASAP7_75t_L g823 ( .A(n_783), .Y(n_823) );
INVx2_ASAP7_75t_L g878 ( .A(n_783), .Y(n_878) );
INVx1_ASAP7_75t_L g918 ( .A(n_783), .Y(n_918) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_785), .A2(n_1118), .B1(n_1124), .B2(n_1135), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1774 ( .A1(n_785), .A2(n_977), .B1(n_1775), .B2(n_1776), .Y(n_1774) );
OA33x2_ASAP7_75t_L g1046 ( .A1(n_786), .A2(n_1047), .A3(n_1048), .B1(n_1051), .B2(n_1052), .B3(n_1055), .Y(n_1046) );
OAI33xp33_ASAP7_75t_L g1175 ( .A1(n_786), .A2(n_1047), .A3(n_1176), .B1(n_1179), .B2(n_1182), .B3(n_1186), .Y(n_1175) );
OAI22xp5_ASAP7_75t_SL g1331 ( .A1(n_786), .A2(n_817), .B1(n_1332), .B2(n_1337), .Y(n_1331) );
OAI33xp33_ASAP7_75t_L g1768 ( .A1(n_786), .A2(n_1769), .A3(n_1773), .B1(n_1774), .B2(n_1777), .B3(n_1780), .Y(n_1768) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
XNOR2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_894), .Y(n_791) );
XNOR2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_855), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_829), .C(n_842), .Y(n_794) );
NOR2xp33_ASAP7_75t_SL g795 ( .A(n_796), .B(n_816), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_799), .A2(n_815), .B1(n_821), .B2(n_823), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g1300 ( .A1(n_800), .A2(n_1301), .B1(n_1302), .B2(n_1304), .Y(n_1300) );
INVx1_ASAP7_75t_L g1763 ( .A(n_800), .Y(n_1763) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B1(n_805), .B2(n_807), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_802), .A2(n_809), .B1(n_821), .B2(n_823), .Y(n_820) );
INVx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx3_ASAP7_75t_L g966 ( .A(n_804), .Y(n_966) );
INVx3_ASAP7_75t_L g1209 ( .A(n_804), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1310 ( .A(n_804), .Y(n_1310) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_806), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_807), .A2(n_812), .B1(n_819), .B2(n_826), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_810), .A2(n_952), .B1(n_963), .B2(n_964), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_810), .A2(n_1205), .B1(n_1206), .B2(n_1207), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_810), .A2(n_1209), .B1(n_1210), .B2(n_1211), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_810), .A2(n_1310), .B1(n_1311), .B2(n_1312), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1470 ( .A1(n_810), .A2(n_1310), .B1(n_1471), .B2(n_1472), .Y(n_1470) );
BUFx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI33xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .A3(n_820), .B1(n_824), .B2(n_825), .B3(n_828), .Y(n_816) );
OAI33xp33_ASAP7_75t_L g973 ( .A1(n_817), .A2(n_828), .A3(n_974), .B1(n_975), .B2(n_976), .B3(n_978), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_819), .A2(n_865), .B1(n_868), .B2(n_874), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_819), .A2(n_874), .B1(n_960), .B2(n_971), .Y(n_974) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g977 ( .A(n_822), .Y(n_977) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI31xp33_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_837), .A3(n_840), .B(n_841), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_831), .A2(n_877), .B1(n_963), .B2(n_967), .Y(n_975) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g1330 ( .A(n_838), .Y(n_1330) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_SL g909 ( .A(n_839), .B(n_910), .Y(n_909) );
OAI31xp33_ASAP7_75t_SL g1024 ( .A1(n_841), .A2(n_1025), .A3(n_1026), .B(n_1030), .Y(n_1024) );
INVx1_ASAP7_75t_L g1248 ( .A(n_841), .Y(n_1248) );
OAI31xp33_ASAP7_75t_L g1256 ( .A1(n_841), .A2(n_1257), .A3(n_1261), .B(n_1262), .Y(n_1256) );
OAI31xp33_ASAP7_75t_SL g842 ( .A1(n_843), .A2(n_844), .A3(n_853), .B(n_854), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx3_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
OAI31xp33_ASAP7_75t_SL g887 ( .A1(n_854), .A2(n_888), .A3(n_889), .B(n_890), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g980 ( .A1(n_854), .A2(n_981), .B(n_987), .Y(n_980) );
NAND3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_880), .C(n_887), .Y(n_856) );
NOR2xp33_ASAP7_75t_SL g857 ( .A(n_858), .B(n_872), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g1201 ( .A1(n_861), .A2(n_1113), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_862), .A2(n_871), .B1(n_877), .B2(n_878), .Y(n_876) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_877), .Y(n_1183) );
INVx2_ASAP7_75t_L g1339 ( .A(n_877), .Y(n_1339) );
XOR2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_955), .Y(n_894) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_929), .B(n_931), .Y(n_896) );
OAI21xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_917), .B(n_921), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_914), .A2(n_916), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1133 ( .A1(n_914), .A2(n_916), .B1(n_1111), .B2(n_1130), .Y(n_1133) );
OAI22xp33_ASAP7_75t_L g1176 ( .A1(n_914), .A2(n_916), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
OAI22xp33_ASAP7_75t_L g1218 ( .A1(n_914), .A2(n_1202), .B1(n_1213), .B2(n_1219), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_916), .A2(n_1119), .B1(n_1125), .B2(n_1138), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_916), .A2(n_1138), .B1(n_1187), .B2(n_1188), .Y(n_1186) );
OAI22xp5_ASAP7_75t_SL g1220 ( .A1(n_918), .A2(n_1206), .B1(n_1210), .B2(n_1221), .Y(n_1220) );
OAI211xp5_ASAP7_75t_SL g921 ( .A1(n_922), .A2(n_923), .B(n_924), .C(n_927), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_923), .A2(n_1114), .B1(n_1131), .B2(n_1135), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g1182 ( .A1(n_923), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1182) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
BUFx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NAND2xp5_ASAP7_75t_SL g932 ( .A(n_933), .B(n_939), .Y(n_932) );
INVx1_ASAP7_75t_L g1172 ( .A(n_940), .Y(n_1172) );
OAI211xp5_ASAP7_75t_L g943 ( .A1(n_944), .A2(n_945), .B(n_947), .C(n_949), .Y(n_943) );
INVx2_ASAP7_75t_SL g945 ( .A(n_946), .Y(n_945) );
BUFx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx3_ASAP7_75t_L g1010 ( .A(n_953), .Y(n_1010) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_953), .Y(n_1205) );
NAND3xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_980), .C(n_990), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_958), .B(n_973), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_968), .A2(n_1306), .B1(n_1307), .B2(n_1308), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g1467 ( .A1(n_968), .A2(n_1009), .B1(n_1468), .B2(n_1469), .Y(n_1467) );
INVx2_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1266 ( .A(n_989), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_989), .A2(n_1045), .B1(n_1328), .B2(n_1329), .Y(n_1348) );
AOI22xp5_ASAP7_75t_L g1516 ( .A1(n_989), .A2(n_1500), .B1(n_1501), .B2(n_1517), .Y(n_1516) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_996), .A2(n_1328), .B1(n_1329), .B2(n_1330), .Y(n_1327) );
XNOR2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1351), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1250), .B1(n_1349), .B2(n_1350), .Y(n_1001) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1002), .Y(n_1349) );
XOR2xp5_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1103), .Y(n_1002) );
XNOR2x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1056), .Y(n_1003) );
NAND4xp75_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1024), .C(n_1032), .D(n_1046), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1016), .B1(n_1017), .B2(n_1023), .Y(n_1007) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1015), .Y(n_1440) );
OAI33xp33_ASAP7_75t_L g1299 ( .A1(n_1016), .A2(n_1126), .A3(n_1300), .B1(n_1305), .B2(n_1309), .B3(n_1313), .Y(n_1299) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
OAI33xp33_ASAP7_75t_L g1783 ( .A1(n_1023), .A2(n_1286), .A3(n_1784), .B1(n_1788), .B2(n_1790), .B3(n_1792), .Y(n_1783) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_1035), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_1037), .Y(n_1168) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_1037), .A2(n_1112), .B1(n_1178), .B2(n_1185), .Y(n_1193) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1407 ( .A1(n_1043), .A2(n_1045), .B1(n_1408), .B2(n_1409), .Y(n_1407) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_1045), .A2(n_1149), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
OAI22xp33_ASAP7_75t_L g1485 ( .A1(n_1047), .A2(n_1486), .B1(n_1491), .B2(n_1497), .Y(n_1485) );
AND3x1_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1067), .C(n_1097), .Y(n_1057) );
NOR2xp33_ASAP7_75t_SL g1067 ( .A(n_1068), .B(n_1085), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_1075), .A2(n_1080), .B1(n_1093), .B2(n_1095), .Y(n_1092) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1079), .Y(n_1123) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1282 ( .A1(n_1093), .A2(n_1095), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1094), .Y(n_1138) );
INVx3_ASAP7_75t_L g1771 ( .A(n_1094), .Y(n_1771) );
BUFx3_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
XNOR2xp5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1196), .Y(n_1103) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1155), .B1(n_1194), .B2(n_1195), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1106), .Y(n_1195) );
NAND3xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1139), .C(n_1146), .Y(n_1107) );
NOR2xp33_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1132), .Y(n_1108) );
OAI22xp33_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1112), .B1(n_1114), .B2(n_1115), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1463 ( .A1(n_1112), .A2(n_1464), .B1(n_1465), .B2(n_1466), .Y(n_1463) );
BUFx4f_ASAP7_75t_SL g1112 ( .A(n_1113), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1115 ( .A(n_1116), .Y(n_1115) );
INVxp67_ASAP7_75t_SL g1466 ( .A(n_1116), .Y(n_1466) );
OAI22xp5_ASAP7_75t_L g1788 ( .A1(n_1120), .A2(n_1775), .B1(n_1781), .B2(n_1789), .Y(n_1788) );
OAI22xp5_ASAP7_75t_L g1790 ( .A1(n_1120), .A2(n_1776), .B1(n_1782), .B2(n_1791), .Y(n_1790) );
INVx3_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g1436 ( .A(n_1127), .B(n_1437), .C(n_1438), .Y(n_1436) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1528 ( .A(n_1128), .Y(n_1528) );
OAI31xp33_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1150), .A3(n_1153), .B(n_1154), .Y(n_1146) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI31xp33_ASAP7_75t_L g1165 ( .A1(n_1154), .A2(n_1166), .A3(n_1167), .B(n_1171), .Y(n_1165) );
OAI31xp33_ASAP7_75t_L g1759 ( .A1(n_1154), .A2(n_1760), .A3(n_1761), .B(n_1766), .Y(n_1759) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1155), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1165), .C(n_1174), .Y(n_1156) );
OAI31xp33_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .A3(n_1163), .B(n_1164), .Y(n_1157) );
OAI31xp33_ASAP7_75t_L g1453 ( .A1(n_1164), .A2(n_1454), .A3(n_1458), .B(n_1460), .Y(n_1453) );
OAI31xp33_ASAP7_75t_L g1752 ( .A1(n_1164), .A2(n_1753), .A3(n_1757), .B(n_1758), .Y(n_1752) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1189), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVxp67_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NOR4xp25_ASAP7_75t_L g1249 ( .A(n_1200), .B(n_1216), .C(n_1225), .D(n_1240), .Y(n_1249) );
INVxp67_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1477 ( .A1(n_1219), .A2(n_1464), .B1(n_1474), .B2(n_1478), .Y(n_1477) );
INVxp67_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
AOI31xp33_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1232), .A3(n_1235), .B(n_1238), .Y(n_1225) );
INVxp67_ASAP7_75t_SL g1227 ( .A(n_1228), .Y(n_1227) );
AOI31xp33_ASAP7_75t_L g1342 ( .A1(n_1238), .A2(n_1343), .A3(n_1347), .B(n_1348), .Y(n_1342) );
CKINVDCx14_ASAP7_75t_R g1238 ( .A(n_1239), .Y(n_1238) );
AOI31xp67_ASAP7_75t_SL g1240 ( .A1(n_1241), .A2(n_1243), .A3(n_1246), .B(n_1248), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
INVxp67_ASAP7_75t_SL g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1250), .Y(n_1350) );
AOI22xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1252), .B1(n_1295), .B2(n_1296), .Y(n_1250) );
INVxp67_ASAP7_75t_SL g1251 ( .A(n_1252), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1263), .C(n_1271), .Y(n_1255) );
NOR2xp33_ASAP7_75t_SL g1271 ( .A(n_1272), .B(n_1285), .Y(n_1271) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
NOR4xp25_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1316), .C(n_1331), .D(n_1342), .Y(n_1298) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1323), .B(n_1507), .Y(n_1506) );
BUFx2_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1336), .Y(n_1496) );
INVx3_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
BUFx2_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
AOI22xp5_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1441), .B1(n_1442), .B2(n_1529), .Y(n_1353) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1354), .Y(n_1529) );
XNOR2xp5_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1396), .Y(n_1354) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1356), .Y(n_1394) );
NAND4xp75_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1367), .C(n_1374), .D(n_1382), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1366), .Y(n_1361) );
AO21x1_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1372), .B(n_1373), .Y(n_1367) );
AOI31xp33_ASAP7_75t_L g1511 ( .A1(n_1373), .A2(n_1512), .A3(n_1515), .B(n_1516), .Y(n_1511) );
INVx2_ASAP7_75t_SL g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1398 ( .A(n_1399), .B(n_1402), .C(n_1407), .Y(n_1398) );
NAND3xp33_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1413), .C(n_1418), .Y(n_1410) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
NAND4xp25_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1429), .C(n_1432), .D(n_1436), .Y(n_1419) );
NAND3xp33_ASAP7_75t_L g1420 ( .A(n_1421), .B(n_1426), .C(n_1428), .Y(n_1420) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
XNOR2xp5_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1483), .Y(n_1442) );
NAND3xp33_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1453), .C(n_1461), .Y(n_1444) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1476), .Y(n_1461) );
INVx2_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
NOR4xp25_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1498), .C(n_1511), .D(n_1519), .Y(n_1484) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
OAI221xp5_ASAP7_75t_SL g1530 ( .A1(n_1531), .A2(n_1747), .B1(n_1750), .B2(n_1793), .C(n_1796), .Y(n_1530) );
AND5x1_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1680), .C(n_1695), .D(n_1724), .E(n_1732), .Y(n_1531) );
AOI21xp5_ASAP7_75t_L g1532 ( .A1(n_1533), .A2(n_1629), .B(n_1633), .Y(n_1532) );
NAND5xp2_ASAP7_75t_L g1533 ( .A(n_1534), .B(n_1584), .C(n_1599), .D(n_1612), .E(n_1627), .Y(n_1533) );
AOI21xp5_ASAP7_75t_L g1534 ( .A1(n_1535), .A2(n_1566), .B(n_1575), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1551), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1536), .B(n_1553), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1536), .B(n_1569), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1536), .B(n_1601), .Y(n_1628) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1536), .B(n_1658), .Y(n_1657) );
CKINVDCx14_ASAP7_75t_R g1689 ( .A(n_1536), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1536), .B(n_1607), .Y(n_1714) );
NAND2xp5_ASAP7_75t_L g1723 ( .A(n_1536), .B(n_1610), .Y(n_1723) );
NOR2xp33_ASAP7_75t_L g1739 ( .A(n_1536), .B(n_1606), .Y(n_1739) );
INVx3_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1537), .B(n_1590), .Y(n_1589) );
CKINVDCx5p33_ASAP7_75t_R g1596 ( .A(n_1537), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1537), .B(n_1597), .Y(n_1604) );
AOI311xp33_ASAP7_75t_L g1612 ( .A1(n_1537), .A2(n_1613), .A3(n_1615), .B(n_1617), .C(n_1621), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1537), .B(n_1554), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1537), .B(n_1665), .Y(n_1664) );
OR2x2_ASAP7_75t_L g1678 ( .A(n_1537), .B(n_1667), .Y(n_1678) );
AND2x4_ASAP7_75t_SL g1537 ( .A(n_1538), .B(n_1546), .Y(n_1537) );
AND2x4_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1541), .Y(n_1539) );
AND2x6_ASAP7_75t_L g1544 ( .A(n_1540), .B(n_1545), .Y(n_1544) );
AND2x6_ASAP7_75t_L g1547 ( .A(n_1540), .B(n_1548), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1540), .B(n_1550), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1540), .B(n_1550), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1540), .B(n_1550), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1540), .B(n_1541), .Y(n_1749) );
HB1xp67_ASAP7_75t_L g1806 ( .A(n_1541), .Y(n_1806) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1543), .Y(n_1541) );
A2O1A1Ixp33_ASAP7_75t_L g1680 ( .A1(n_1551), .A2(n_1655), .B(n_1681), .C(n_1692), .Y(n_1680) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
NOR2xp33_ASAP7_75t_L g1712 ( .A(n_1552), .B(n_1713), .Y(n_1712) );
NOR2xp33_ASAP7_75t_L g1731 ( .A(n_1552), .B(n_1642), .Y(n_1731) );
OR2x2_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1557), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1553), .B(n_1597), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1553), .B(n_1563), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1553), .B(n_1558), .Y(n_1654) );
NOR2xp33_ASAP7_75t_L g1662 ( .A(n_1553), .B(n_1663), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1553), .B(n_1610), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1553), .B(n_1625), .Y(n_1690) );
OR2x2_ASAP7_75t_L g1699 ( .A(n_1553), .B(n_1591), .Y(n_1699) );
OR2x2_ASAP7_75t_L g1734 ( .A(n_1553), .B(n_1723), .Y(n_1734) );
INVx2_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1554), .B(n_1595), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1616 ( .A(n_1554), .B(n_1563), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1554), .B(n_1598), .Y(n_1619) );
OR2x2_ASAP7_75t_L g1667 ( .A(n_1554), .B(n_1558), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1668 ( .A(n_1554), .B(n_1558), .Y(n_1668) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1554), .B(n_1597), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1711 ( .A(n_1554), .B(n_1604), .Y(n_1711) );
OR2x2_ASAP7_75t_L g1720 ( .A(n_1554), .B(n_1591), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1556), .Y(n_1554) );
NOR2xp33_ASAP7_75t_L g1575 ( .A(n_1557), .B(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1557), .Y(n_1625) );
OR2x2_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1562), .Y(n_1557) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1558), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1558), .B(n_1563), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1560), .Y(n_1558) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
OR2x2_ASAP7_75t_L g1591 ( .A(n_1563), .B(n_1592), .Y(n_1591) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1563), .Y(n_1598) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1563), .Y(n_1742) );
NAND2x1_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
AOI322xp5_ASAP7_75t_L g1660 ( .A1(n_1566), .A2(n_1628), .A3(n_1635), .B1(n_1661), .B2(n_1662), .C1(n_1666), .C2(n_1670), .Y(n_1660) );
OAI21xp33_ASAP7_75t_L g1721 ( .A1(n_1566), .A2(n_1719), .B(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1567), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1572), .Y(n_1567) );
INVx2_ASAP7_75t_L g1614 ( .A(n_1568), .Y(n_1614) );
AOI321xp33_ASAP7_75t_L g1671 ( .A1(n_1568), .A2(n_1652), .A3(n_1672), .B1(n_1673), .B2(n_1675), .C(n_1677), .Y(n_1671) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1569), .B(n_1583), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1602 ( .A(n_1569), .B(n_1572), .Y(n_1602) );
INVx2_ASAP7_75t_SL g1607 ( .A(n_1569), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1569), .B(n_1641), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1571), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_1572), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1572), .B(n_1578), .Y(n_1593) );
HB1xp67_ASAP7_75t_SL g1691 ( .A(n_1572), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1572), .B(n_1579), .Y(n_1728) );
AND2x4_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1574), .Y(n_1572) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1576), .Y(n_1649) );
OR2x2_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1582), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1577), .B(n_1656), .Y(n_1655) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1578), .B(n_1587), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1578), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1578), .B(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1578), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_1578), .B(n_1629), .Y(n_1674) );
NAND3xp33_ASAP7_75t_L g1746 ( .A(n_1578), .B(n_1590), .C(n_1714), .Y(n_1746) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1579), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1579), .B(n_1583), .Y(n_1652) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1579), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1581), .Y(n_1579) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1582), .Y(n_1694) );
OR2x2_ASAP7_75t_L g1606 ( .A(n_1583), .B(n_1607), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1583), .B(n_1669), .Y(n_1670) );
OAI32xp33_ASAP7_75t_L g1700 ( .A1(n_1583), .A2(n_1595), .A3(n_1644), .B1(n_1656), .B2(n_1701), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1583), .B(n_1629), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1583), .B(n_1656), .Y(n_1715) );
AOI211xp5_ASAP7_75t_L g1716 ( .A1(n_1583), .A2(n_1614), .B(n_1629), .C(n_1717), .Y(n_1716) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_1585), .A2(n_1588), .B1(n_1593), .B2(n_1594), .Y(n_1584) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
OAI311xp33_ASAP7_75t_L g1650 ( .A1(n_1589), .A2(n_1629), .A3(n_1651), .B1(n_1653), .C1(n_1659), .Y(n_1650) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1590), .B(n_1637), .Y(n_1636) );
OAI211xp5_ASAP7_75t_L g1653 ( .A1(n_1590), .A2(n_1654), .B(n_1655), .C(n_1657), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1661 ( .A(n_1590), .B(n_1625), .Y(n_1661) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1592), .B(n_1598), .Y(n_1597) );
NAND3xp33_ASAP7_75t_L g1659 ( .A(n_1593), .B(n_1614), .C(n_1624), .Y(n_1659) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1593), .Y(n_1679) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1594), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1597), .Y(n_1595) );
OR2x2_ASAP7_75t_L g1647 ( .A(n_1596), .B(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1596), .Y(n_1686) );
OAI32xp33_ASAP7_75t_L g1724 ( .A1(n_1596), .A2(n_1601), .A3(n_1725), .B1(n_1729), .B2(n_1731), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1596), .B(n_1619), .Y(n_1745) );
AOI21xp5_ASAP7_75t_L g1599 ( .A1(n_1600), .A2(n_1603), .B(n_1605), .Y(n_1599) );
AOI22xp5_ASAP7_75t_L g1681 ( .A1(n_1601), .A2(n_1682), .B1(n_1687), .B2(n_1691), .Y(n_1681) );
INVx2_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1603), .Y(n_1735) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1608), .Y(n_1605) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1606), .Y(n_1623) );
OAI21xp33_ASAP7_75t_L g1696 ( .A1(n_1606), .A2(n_1697), .B(n_1700), .Y(n_1696) );
INVx2_ASAP7_75t_L g1658 ( .A(n_1607), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1607), .B(n_1688), .Y(n_1687) );
NOR2xp33_ASAP7_75t_L g1710 ( .A(n_1607), .B(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1608), .Y(n_1641) );
OR2x2_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1611), .Y(n_1608) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1610), .B(n_1628), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1610), .B(n_1626), .Y(n_1676) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1611), .Y(n_1637) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1613), .Y(n_1736) );
A2O1A1Ixp33_ASAP7_75t_L g1634 ( .A1(n_1614), .A2(n_1635), .B(n_1638), .C(n_1642), .Y(n_1634) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1614), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1614), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1620), .Y(n_1618) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
AOI21xp5_ASAP7_75t_L g1692 ( .A1(n_1623), .A2(n_1693), .B(n_1694), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
INVx3_ASAP7_75t_L g1656 ( .A(n_1629), .Y(n_1656) );
NOR3xp33_ASAP7_75t_L g1677 ( .A(n_1629), .B(n_1678), .C(n_1679), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1632), .Y(n_1629) );
NAND4xp25_ASAP7_75t_SL g1633 ( .A(n_1634), .B(n_1643), .C(n_1660), .D(n_1671), .Y(n_1633) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1640), .B(n_1641), .Y(n_1639) );
O2A1O1Ixp33_ASAP7_75t_L g1643 ( .A1(n_1644), .A2(n_1646), .B(n_1649), .C(n_1650), .Y(n_1643) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
OAI21xp5_ASAP7_75t_SL g1732 ( .A1(n_1656), .A2(n_1733), .B(n_1737), .Y(n_1732) );
NOR2xp33_ASAP7_75t_L g1683 ( .A(n_1658), .B(n_1684), .Y(n_1683) );
OAI221xp5_ASAP7_75t_L g1708 ( .A1(n_1658), .A2(n_1709), .B1(n_1716), .B2(n_1718), .C(n_1721), .Y(n_1708) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
AOI21xp33_ASAP7_75t_L g1666 ( .A1(n_1667), .A2(n_1668), .B(n_1669), .Y(n_1666) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1669), .Y(n_1740) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1670), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1672), .B(n_1686), .Y(n_1685) );
NOR2xp33_ASAP7_75t_L g1697 ( .A(n_1672), .B(n_1698), .Y(n_1697) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
OAI311xp33_ASAP7_75t_L g1695 ( .A1(n_1674), .A2(n_1696), .A3(n_1702), .B1(n_1707), .C1(n_1708), .Y(n_1695) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1678), .Y(n_1717) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
NOR4xp25_ASAP7_75t_L g1709 ( .A(n_1685), .B(n_1710), .C(n_1712), .D(n_1715), .Y(n_1709) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1687), .Y(n_1707) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1688), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1689), .B(n_1719), .Y(n_1718) );
INVx2_ASAP7_75t_L g1726 ( .A(n_1690), .Y(n_1726) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1694), .Y(n_1703) );
INVx2_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
OAI21xp33_ASAP7_75t_SL g1702 ( .A1(n_1703), .A2(n_1704), .B(n_1706), .Y(n_1702) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
AOI21xp33_ASAP7_75t_L g1725 ( .A1(n_1706), .A2(n_1726), .B(n_1727), .Y(n_1725) );
AOI21xp33_ASAP7_75t_L g1729 ( .A1(n_1706), .A2(n_1727), .B(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
AOI21xp33_ASAP7_75t_L g1733 ( .A1(n_1734), .A2(n_1735), .B(n_1736), .Y(n_1733) );
OAI321xp33_ASAP7_75t_L g1737 ( .A1(n_1738), .A2(n_1740), .A3(n_1741), .B1(n_1743), .B2(n_1744), .C(n_1746), .Y(n_1737) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
CKINVDCx20_ASAP7_75t_R g1747 ( .A(n_1748), .Y(n_1747) );
CKINVDCx5p33_ASAP7_75t_R g1748 ( .A(n_1749), .Y(n_1748) );
HB1xp67_ASAP7_75t_L g1799 ( .A(n_1751), .Y(n_1799) );
NAND3xp33_ASAP7_75t_SL g1751 ( .A(n_1752), .B(n_1759), .C(n_1767), .Y(n_1751) );
INVx2_ASAP7_75t_SL g1762 ( .A(n_1763), .Y(n_1762) );
NOR2xp33_ASAP7_75t_SL g1767 ( .A(n_1768), .B(n_1783), .Y(n_1767) );
OAI22xp33_ASAP7_75t_L g1784 ( .A1(n_1770), .A2(n_1778), .B1(n_1785), .B2(n_1787), .Y(n_1784) );
INVx2_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
CKINVDCx5p33_ASAP7_75t_R g1793 ( .A(n_1794), .Y(n_1793) );
INVxp33_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
HB1xp67_ASAP7_75t_SL g1800 ( .A(n_1801), .Y(n_1800) );
BUFx3_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
HB1xp67_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
OAI21xp5_ASAP7_75t_L g1804 ( .A1(n_1805), .A2(n_1806), .B(n_1807), .Y(n_1804) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
endmodule