module fake_jpeg_5283_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_8),
.B(n_14),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_32),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_48),
.B(n_57),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_29),
.B1(n_25),
.B2(n_21),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_18),
.B1(n_34),
.B2(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_24),
.B1(n_20),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_24),
.B1(n_20),
.B2(n_35),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_21),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_66),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_27),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_71),
.B1(n_68),
.B2(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_35),
.B1(n_39),
.B2(n_18),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_76),
.Y(n_104)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_34),
.B1(n_39),
.B2(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_87),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_85),
.B1(n_75),
.B2(n_66),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_39),
.B1(n_34),
.B2(n_27),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_39),
.B1(n_34),
.B2(n_27),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_88),
.C(n_44),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_16),
.B1(n_17),
.B2(n_22),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_40),
.C(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_105),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_86),
.B1(n_81),
.B2(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_47),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_61),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_44),
.B1(n_52),
.B2(n_48),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_81),
.B1(n_75),
.B2(n_54),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_65),
.B(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_70),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_122),
.C(n_135),
.Y(n_160)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_130),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_54),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_127),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_98),
.B(n_104),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_139),
.Y(n_147)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_40),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_54),
.C(n_40),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_92),
.B(n_12),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_23),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_93),
.B(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_142),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_31),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_40),
.B1(n_72),
.B2(n_76),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_89),
.B1(n_95),
.B2(n_94),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_113),
.B(n_108),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_146),
.B(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_155),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_99),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_119),
.A3(n_139),
.B1(n_136),
.B2(n_142),
.C1(n_127),
.C2(n_116),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_104),
.B(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_166),
.B1(n_146),
.B2(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_97),
.B1(n_110),
.B2(n_109),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_165),
.B1(n_141),
.B2(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_102),
.B(n_112),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_22),
.B1(n_31),
.B2(n_28),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_110),
.B1(n_107),
.B2(n_72),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_169),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_87),
.C(n_31),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_170),
.C(n_135),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_117),
.B(n_23),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_185),
.C(n_164),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_144),
.C(n_170),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_183),
.C(n_195),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_190),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_147),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_123),
.B1(n_87),
.B2(n_22),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_138),
.C(n_31),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_23),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_28),
.B(n_26),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_194),
.C(n_169),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_155),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_138),
.B(n_28),
.C(n_26),
.D(n_3),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_28),
.C(n_26),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_147),
.C(n_165),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_209),
.C(n_210),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_194),
.B(n_192),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_217),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_158),
.B1(n_143),
.B2(n_163),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_212),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_175),
.C(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_159),
.C(n_163),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_172),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_178),
.C(n_195),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_171),
.C(n_153),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_197),
.A2(n_177),
.B1(n_188),
.B2(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_233),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_177),
.B1(n_174),
.B2(n_196),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_204),
.B1(n_201),
.B2(n_198),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_226),
.A2(n_7),
.B(n_13),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_191),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_200),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_172),
.B1(n_153),
.B2(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_241),
.C(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_198),
.C(n_1),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_222),
.B(n_231),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_7),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_8),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_221),
.C(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_247),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_223),
.B(n_224),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_251),
.B(n_255),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_254),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_225),
.B(n_228),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_236),
.C(n_244),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_260),
.B(n_10),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_230),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_219),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_234),
.B1(n_235),
.B2(n_238),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_219),
.A3(n_9),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_256),
.B(n_11),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_259),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_10),
.B(n_13),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_9),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_258),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_10),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_271),
.C(n_11),
.Y(n_276)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_275),
.A3(n_11),
.B1(n_2),
.B2(n_6),
.C1(n_12),
.C2(n_15),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_277),
.A2(n_6),
.B(n_15),
.C(n_0),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_1),
.Y(n_279)
);


endmodule