module fake_ibex_604_n_3712 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3712);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3712;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_641;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_2333;
wire n_715;
wire n_1910;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2806;
wire n_2283;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_709;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2451;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_3054;
wire n_2924;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_1036;
wire n_974;
wire n_1831;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2910;
wire n_2552;
wire n_3331;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_705;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_847;
wire n_2699;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1599;
wire n_712;
wire n_1539;
wire n_1400;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_650;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2698;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_648;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_3162;
wire n_2732;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_768;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2348;
wire n_2093;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_631;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2816;
wire n_2803;
wire n_2433;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2653;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_665;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_720;
wire n_1390;
wire n_710;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_759;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_3015;
wire n_2588;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_635;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2148;
wire n_949;
wire n_2357;
wire n_704;
wire n_2104;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2349;
wire n_2100;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

INVx1_ASAP7_75t_L g629 ( 
.A(n_442),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_502),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_123),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_505),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_424),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_8),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_487),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_624),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_601),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_552),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_608),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_244),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_137),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_293),
.Y(n_643)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_197),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_526),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_609),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_186),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_317),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_365),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_520),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_398),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_596),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_380),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_34),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_432),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_286),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_391),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_171),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_470),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_22),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_272),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_319),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_330),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_517),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_612),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_53),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_298),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_333),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_48),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_490),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_143),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_485),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_589),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_563),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_152),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_331),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_96),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_448),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_329),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_92),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_558),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_122),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_621),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_506),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_559),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_568),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_597),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_494),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_184),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_342),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_514),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_207),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_0),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_69),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_219),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_131),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_389),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_459),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_307),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_230),
.Y(n_700)
);

INVxp33_ASAP7_75t_R g701 ( 
.A(n_81),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_489),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_346),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_488),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_221),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_416),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_583),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_313),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_595),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_478),
.Y(n_710)
);

BUFx2_ASAP7_75t_SL g711 ( 
.A(n_549),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_577),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_594),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_451),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_399),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_566),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_570),
.Y(n_717)
);

BUFx5_ASAP7_75t_L g718 ( 
.A(n_272),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_551),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_28),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_579),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_264),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_150),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_301),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_290),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_288),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_282),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_51),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_553),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_592),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_456),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_507),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_273),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_113),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_581),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_354),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_585),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_161),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_530),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_344),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_344),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_274),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_511),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_169),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_92),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_160),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_288),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_53),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_550),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_183),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_188),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_320),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_259),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_324),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_442),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_572),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_195),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_616),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_593),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_10),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_332),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_223),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_407),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_543),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_250),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_94),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_498),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_452),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_394),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_266),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_460),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_7),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_411),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_391),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_357),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_70),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_41),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_576),
.Y(n_778)
);

CKINVDCx14_ASAP7_75t_R g779 ( 
.A(n_610),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_279),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_93),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_160),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_569),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_195),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_306),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_617),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_64),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_424),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_409),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_333),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_231),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_499),
.Y(n_792)
);

INVxp33_ASAP7_75t_L g793 ( 
.A(n_28),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_546),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_512),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_421),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_375),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_82),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_121),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_402),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_386),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_573),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_100),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_243),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_76),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_197),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_65),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_31),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_582),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_544),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_76),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_87),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_574),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_510),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_364),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_351),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_440),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_562),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_116),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_353),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_547),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_325),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_148),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_208),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_555),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_347),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_425),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_30),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_289),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_21),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_253),
.Y(n_831)
);

CKINVDCx14_ASAP7_75t_R g832 ( 
.A(n_627),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_152),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_584),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_140),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_348),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_414),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_149),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_163),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_432),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_103),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_109),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_205),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_177),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_229),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_557),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_249),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_298),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_591),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_397),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_375),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_5),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_540),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_182),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_429),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_34),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_542),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_352),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_345),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_388),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_412),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_611),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_126),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_367),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_605),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_454),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_541),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_245),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_388),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_516),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_15),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_263),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_110),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_423),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_451),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_561),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_380),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_93),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_538),
.Y(n_879)
);

CKINVDCx16_ASAP7_75t_R g880 ( 
.A(n_119),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_599),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_165),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_497),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_349),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_238),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_310),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_71),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_345),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_477),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_327),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_156),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_440),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_534),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_491),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_284),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_586),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_191),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_118),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_134),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_103),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_357),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_509),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_450),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_513),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_613),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_130),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_252),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_330),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_495),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_290),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_620),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_443),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_37),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_548),
.Y(n_914)
);

BUFx10_ASAP7_75t_L g915 ( 
.A(n_332),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_157),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_564),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_607),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_5),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_405),
.Y(n_920)
);

CKINVDCx16_ASAP7_75t_R g921 ( 
.A(n_580),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_112),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_253),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_503),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_571),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_369),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_602),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_455),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_397),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_25),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_82),
.Y(n_931)
);

BUFx5_ASAP7_75t_L g932 ( 
.A(n_554),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_4),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_587),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_468),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_604),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_588),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_619),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_296),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_463),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_68),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_387),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_565),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_80),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_521),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_208),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_88),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_450),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_257),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_188),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_600),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_372),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_426),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_43),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_373),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_282),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_614),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_90),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_111),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_598),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_59),
.Y(n_961)
);

BUFx8_ASAP7_75t_SL g962 ( 
.A(n_177),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_311),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_444),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_189),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_545),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_415),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_228),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_216),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_10),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_144),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_255),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_289),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_247),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_189),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_87),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_383),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_307),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_590),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_351),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_27),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_164),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_172),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_147),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_49),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_293),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_193),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_575),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_54),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_146),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_147),
.Y(n_991)
);

BUFx5_ASAP7_75t_L g992 ( 
.A(n_201),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_110),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_271),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_303),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_238),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_411),
.Y(n_997)
);

CKINVDCx14_ASAP7_75t_R g998 ( 
.A(n_415),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_389),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_81),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_18),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_216),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_295),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_578),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_169),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_615),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_221),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_473),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_623),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_402),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_567),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_122),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_146),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_48),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_254),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_196),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_144),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_153),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_508),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_606),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_618),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_209),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_365),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_331),
.Y(n_1024)
);

BUFx8_ASAP7_75t_SL g1025 ( 
.A(n_240),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_245),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_273),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_308),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_560),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_107),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_219),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_556),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_266),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_0),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_379),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_3),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_206),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_11),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_77),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_267),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_30),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_176),
.Y(n_1042)
);

CKINVDCx14_ASAP7_75t_R g1043 ( 
.A(n_26),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_60),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_369),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_622),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_9),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_96),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_303),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_341),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_603),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_271),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_682),
.Y(n_1053)
);

BUFx8_ASAP7_75t_SL g1054 ( 
.A(n_962),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_672),
.B(n_1),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_672),
.B(n_1),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_893),
.B(n_2),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_635),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_660),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_655),
.B(n_2),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_745),
.B(n_968),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_635),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_635),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_793),
.B(n_3),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_635),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_756),
.B(n_745),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_640),
.Y(n_1067)
);

INVx5_ASAP7_75t_L g1068 ( 
.A(n_640),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_640),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_900),
.B(n_4),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_640),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_805),
.B(n_6),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_718),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_968),
.B(n_6),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_754),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_984),
.B(n_7),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_793),
.B(n_8),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_984),
.B(n_9),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_754),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_644),
.B(n_880),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_754),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_921),
.B(n_457),
.Y(n_1082)
);

AND2x6_ASAP7_75t_L g1083 ( 
.A(n_698),
.B(n_628),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_718),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_718),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_998),
.B(n_11),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_688),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_671),
.B(n_12),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_754),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_893),
.B(n_12),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_705),
.B(n_13),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_630),
.B(n_13),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_656),
.B(n_14),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_718),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_682),
.Y(n_1095)
);

BUFx12f_ASAP7_75t_L g1096 ( 
.A(n_682),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1043),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_785),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_671),
.B(n_690),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_688),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_656),
.B(n_14),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_785),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_785),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_688),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_718),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_658),
.B(n_661),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_822),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_822),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_690),
.B(n_15),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_658),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_785),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_718),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_734),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_718),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_822),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_632),
.B(n_16),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_915),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_972),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_740),
.Y(n_1119)
);

BUFx8_ASAP7_75t_SL g1120 ( 
.A(n_962),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_L g1121 ( 
.A(n_734),
.B(n_16),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_915),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_740),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_972),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_698),
.B(n_458),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_972),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_629),
.B(n_17),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_972),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_915),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_740),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_762),
.B(n_17),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_767),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1025),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_950),
.B(n_767),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_740),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_661),
.B(n_662),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_662),
.B(n_18),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_991),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_740),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_740),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_950),
.B(n_19),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_950),
.B(n_19),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_667),
.B(n_668),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_991),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_667),
.B(n_20),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_740),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_992),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_638),
.B(n_20),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_762),
.B(n_21),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_767),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_916),
.B(n_22),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_992),
.Y(n_1152)
);

BUFx8_ASAP7_75t_L g1153 ( 
.A(n_992),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_636),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_645),
.B(n_23),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_916),
.B(n_23),
.Y(n_1156)
);

BUFx8_ASAP7_75t_SL g1157 ( 
.A(n_1025),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_991),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_647),
.B(n_24),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_668),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_669),
.B(n_24),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_992),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_669),
.B(n_25),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_766),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_991),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_985),
.B(n_26),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1034),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1034),
.Y(n_1168)
);

BUFx12f_ASAP7_75t_L g1169 ( 
.A(n_766),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_985),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_673),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_992),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_1034),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_646),
.B(n_27),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1005),
.B(n_29),
.Y(n_1175)
);

INVxp33_ASAP7_75t_SL g1176 ( 
.A(n_877),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1005),
.B(n_29),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1018),
.B(n_31),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1100),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1176),
.A2(n_1024),
.B1(n_1027),
.B2(n_877),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1078),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_R g1182 ( 
.A1(n_1059),
.A2(n_701),
.B1(n_720),
.B2(n_654),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1097),
.B(n_779),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1150),
.B(n_832),
.Y(n_1184)
);

OAI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1159),
.A2(n_1027),
.B1(n_1031),
.B2(n_1024),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1080),
.A2(n_1033),
.B1(n_1035),
.B2(n_1031),
.Y(n_1186)
);

AO22x2_ASAP7_75t_L g1187 ( 
.A1(n_1078),
.A2(n_807),
.B1(n_841),
.B2(n_748),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1100),
.Y(n_1188)
);

OA22x2_ASAP7_75t_L g1189 ( 
.A1(n_1133),
.A2(n_1035),
.B1(n_1036),
.B2(n_1033),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1170),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1088),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1088),
.Y(n_1192)
);

AO22x2_ASAP7_75t_L g1193 ( 
.A1(n_1109),
.A2(n_946),
.B1(n_931),
.B2(n_1048),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1171),
.A2(n_679),
.B1(n_787),
.B2(n_746),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1106),
.A2(n_1036),
.B1(n_870),
.B2(n_934),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1136),
.A2(n_870),
.B1(n_934),
.B2(n_673),
.Y(n_1196)
);

OAI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1082),
.A2(n_633),
.B1(n_634),
.B2(n_631),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_1053),
.B(n_711),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1150),
.B(n_707),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1170),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1134),
.B(n_1018),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1109),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1100),
.B(n_1029),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1110),
.B(n_1113),
.Y(n_1204)
);

AO22x2_ASAP7_75t_L g1205 ( 
.A1(n_1131),
.A2(n_1044),
.B1(n_1042),
.B2(n_648),
.Y(n_1205)
);

AO22x2_ASAP7_75t_L g1206 ( 
.A1(n_1131),
.A2(n_663),
.B1(n_666),
.B2(n_657),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1082),
.A2(n_679),
.B1(n_787),
.B2(n_746),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1143),
.A2(n_988),
.B1(n_1046),
.B2(n_960),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1099),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1064),
.A2(n_988),
.B1(n_1046),
.B2(n_960),
.Y(n_1210)
);

AO22x2_ASAP7_75t_L g1211 ( 
.A1(n_1149),
.A2(n_1151),
.B1(n_1178),
.B2(n_1066),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1077),
.A2(n_642),
.B1(n_649),
.B2(n_643),
.Y(n_1212)
);

NAND3x1_ASAP7_75t_L g1213 ( 
.A(n_1054),
.B(n_826),
.C(n_796),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1149),
.A2(n_1178),
.B1(n_1151),
.B2(n_1096),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1104),
.B(n_731),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1104),
.B(n_918),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1099),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1095),
.A2(n_651),
.B1(n_677),
.B2(n_676),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1066),
.A2(n_694),
.B1(n_695),
.B2(n_675),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1107),
.A2(n_1129),
.B1(n_1117),
.B2(n_1115),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1060),
.A2(n_826),
.B1(n_828),
.B2(n_796),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1070),
.A2(n_854),
.B1(n_886),
.B2(n_828),
.Y(n_1222)
);

AO22x2_ASAP7_75t_L g1223 ( 
.A1(n_1061),
.A2(n_700),
.B1(n_722),
.B2(n_699),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1160),
.A2(n_680),
.B1(n_689),
.B2(n_678),
.Y(n_1224)
);

AOI22x1_ASAP7_75t_L g1225 ( 
.A1(n_1073),
.A2(n_862),
.B1(n_650),
.B2(n_665),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1072),
.A2(n_886),
.B1(n_913),
.B2(n_854),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1108),
.B(n_641),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1164),
.A2(n_693),
.B1(n_696),
.B2(n_692),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1061),
.Y(n_1229)
);

AO22x2_ASAP7_75t_L g1230 ( 
.A1(n_1141),
.A2(n_726),
.B1(n_728),
.B2(n_725),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1165),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1156),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1166),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1169),
.A2(n_1086),
.B1(n_1177),
.B2(n_1175),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1108),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1122),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1074),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1122),
.B(n_992),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1076),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1084),
.Y(n_1240)
);

NOR2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1087),
.B(n_760),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1165),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1154),
.B(n_1029),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1104),
.B(n_992),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1093),
.A2(n_703),
.B1(n_714),
.B2(n_697),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1132),
.B(n_652),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_1142),
.A2(n_757),
.B1(n_763),
.B2(n_744),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1165),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1173),
.Y(n_1249)
);

AO22x2_ASAP7_75t_L g1250 ( 
.A1(n_1101),
.A2(n_773),
.B1(n_775),
.B2(n_769),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1132),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1120),
.B(n_641),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1137),
.A2(n_923),
.B1(n_975),
.B2(n_913),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1132),
.B(n_652),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1173),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1145),
.A2(n_975),
.B1(n_990),
.B2(n_923),
.Y(n_1256)
);

AND2x6_ASAP7_75t_L g1257 ( 
.A(n_1121),
.B(n_849),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1157),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1121),
.B(n_653),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1084),
.Y(n_1260)
);

AO22x2_ASAP7_75t_L g1261 ( 
.A1(n_1161),
.A2(n_1163),
.B1(n_1127),
.B2(n_784),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1127),
.A2(n_1030),
.B1(n_990),
.B2(n_790),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1091),
.A2(n_723),
.B1(n_724),
.B2(n_715),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1154),
.B(n_664),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1153),
.A2(n_733),
.B1(n_736),
.B2(n_727),
.Y(n_1265)
);

NAND3x1_ASAP7_75t_L g1266 ( 
.A(n_1092),
.B(n_1030),
.C(n_791),
.Y(n_1266)
);

AO22x2_ASAP7_75t_L g1267 ( 
.A1(n_1085),
.A2(n_803),
.B1(n_808),
.B2(n_777),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1055),
.A2(n_738),
.B1(n_742),
.B2(n_741),
.Y(n_1268)
);

AND2x6_ASAP7_75t_L g1269 ( 
.A(n_1056),
.B(n_849),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1085),
.B(n_664),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1105),
.B(n_1147),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1105),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1112),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1153),
.B(n_670),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1094),
.Y(n_1275)
);

BUFx10_ASAP7_75t_L g1276 ( 
.A(n_1057),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1090),
.A2(n_750),
.B1(n_751),
.B2(n_747),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1116),
.A2(n_753),
.B1(n_755),
.B2(n_752),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1112),
.A2(n_765),
.B1(n_768),
.B2(n_761),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1148),
.A2(n_772),
.B1(n_774),
.B2(n_770),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1155),
.A2(n_776),
.B1(n_781),
.B2(n_780),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1119),
.B(n_670),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1083),
.B(n_782),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1119),
.B(n_653),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1123),
.B(n_706),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1173),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_SL g1287 ( 
.A(n_1123),
.B(n_788),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1174),
.B(n_815),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1083),
.A2(n_798),
.B1(n_799),
.B2(n_789),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1083),
.A2(n_801),
.B1(n_804),
.B2(n_800),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1114),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1139),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1139),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1140),
.B(n_706),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1083),
.A2(n_811),
.B1(n_812),
.B2(n_806),
.Y(n_1295)
);

AO22x2_ASAP7_75t_L g1296 ( 
.A1(n_1140),
.A2(n_1037),
.B1(n_820),
.B2(n_829),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1125),
.A2(n_819),
.B1(n_823),
.B2(n_816),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1146),
.A2(n_831),
.B1(n_833),
.B2(n_817),
.Y(n_1298)
);

AO22x2_ASAP7_75t_L g1299 ( 
.A1(n_1146),
.A2(n_837),
.B1(n_842),
.B2(n_835),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1130),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1147),
.B(n_708),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1135),
.A2(n_830),
.B1(n_836),
.B2(n_824),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1172),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1152),
.B(n_1026),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1162),
.B(n_691),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1075),
.A2(n_839),
.B1(n_840),
.B2(n_838),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1125),
.A2(n_844),
.B1(n_845),
.B2(n_843),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1063),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1125),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1125),
.Y(n_1310)
);

INVx8_ASAP7_75t_L g1311 ( 
.A(n_1063),
.Y(n_1311)
);

AO22x2_ASAP7_75t_L g1312 ( 
.A1(n_1063),
.A2(n_855),
.B1(n_858),
.B2(n_850),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1075),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1065),
.B(n_708),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1065),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1075),
.A2(n_851),
.B1(n_852),
.B2(n_847),
.Y(n_1316)
);

AO22x2_ASAP7_75t_L g1317 ( 
.A1(n_1065),
.A2(n_860),
.B1(n_861),
.B2(n_859),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1068),
.B(n_659),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1079),
.A2(n_864),
.B1(n_869),
.B2(n_856),
.Y(n_1319)
);

OR2x6_ASAP7_75t_L g1320 ( 
.A(n_1079),
.B(n_1002),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1068),
.Y(n_1321)
);

AO22x2_ASAP7_75t_L g1322 ( 
.A1(n_1068),
.A2(n_866),
.B1(n_868),
.B2(n_863),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1079),
.Y(n_1323)
);

AO22x2_ASAP7_75t_L g1324 ( 
.A1(n_1081),
.A2(n_875),
.B1(n_878),
.B2(n_874),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1081),
.B(n_797),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1081),
.B(n_674),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1089),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1089),
.A2(n_872),
.B1(n_882),
.B2(n_871),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1089),
.A2(n_885),
.B1(n_888),
.B2(n_887),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1098),
.A2(n_891),
.B1(n_897),
.B2(n_884),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1098),
.A2(n_892),
.B1(n_895),
.B2(n_890),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1098),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1102),
.B(n_683),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1102),
.A2(n_901),
.B1(n_907),
.B2(n_898),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1102),
.A2(n_920),
.B1(n_922),
.B2(n_910),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1103),
.B(n_681),
.Y(n_1336)
);

AOI22x1_ASAP7_75t_L g1337 ( 
.A1(n_1058),
.A2(n_862),
.B1(n_687),
.B2(n_704),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1103),
.A2(n_903),
.B1(n_906),
.B2(n_899),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1103),
.A2(n_933),
.B1(n_939),
.B2(n_926),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1111),
.A2(n_944),
.B1(n_947),
.B2(n_941),
.Y(n_1340)
);

AO22x2_ASAP7_75t_L g1341 ( 
.A1(n_1111),
.A2(n_912),
.B1(n_919),
.B2(n_908),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1111),
.A2(n_952),
.B1(n_954),
.B2(n_949),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1118),
.A2(n_942),
.B1(n_948),
.B2(n_930),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1118),
.Y(n_1344)
);

AND2x2_ASAP7_75t_SL g1345 ( 
.A(n_1118),
.B(n_797),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1124),
.B(n_827),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1124),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1124),
.A2(n_956),
.B1(n_958),
.B2(n_953),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1126),
.A2(n_959),
.B1(n_964),
.B2(n_955),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1126),
.B(n_827),
.Y(n_1350)
);

AO22x2_ASAP7_75t_L g1351 ( 
.A1(n_1126),
.A2(n_963),
.B1(n_971),
.B2(n_961),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1128),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1128),
.B(n_1038),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1128),
.A2(n_978),
.B1(n_983),
.B2(n_974),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1138),
.B(n_1039),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1138),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1138),
.B(n_1040),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1144),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1144),
.B(n_848),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1144),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1158),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1158),
.B(n_848),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1158),
.A2(n_967),
.B1(n_969),
.B2(n_965),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1167),
.B(n_873),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1167),
.B(n_716),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1167),
.A2(n_973),
.B1(n_976),
.B2(n_970),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1168),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1168),
.A2(n_981),
.B1(n_982),
.B2(n_977),
.Y(n_1368)
);

AO22x2_ASAP7_75t_L g1369 ( 
.A1(n_1168),
.A2(n_1023),
.B1(n_989),
.B2(n_993),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_R g1370 ( 
.A1(n_1058),
.A2(n_995),
.B1(n_1001),
.B2(n_986),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1058),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1062),
.B(n_873),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1062),
.A2(n_1014),
.B1(n_1015),
.B2(n_1003),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1062),
.Y(n_1374)
);

AO22x2_ASAP7_75t_L g1375 ( 
.A1(n_1067),
.A2(n_1016),
.B1(n_980),
.B2(n_1002),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1067),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1067),
.B(n_684),
.Y(n_1377)
);

AO22x1_ASAP7_75t_SL g1378 ( 
.A1(n_1069),
.A2(n_980),
.B1(n_1026),
.B2(n_929),
.Y(n_1378)
);

AO22x2_ASAP7_75t_L g1379 ( 
.A1(n_1069),
.A2(n_1028),
.B1(n_929),
.B2(n_721),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1069),
.B(n_1028),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1071),
.A2(n_1041),
.B1(n_1045),
.B2(n_1022),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1071),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1071),
.A2(n_1049),
.B1(n_1050),
.B2(n_1047),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1080),
.A2(n_994),
.B1(n_996),
.B2(n_987),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1080),
.A2(n_999),
.B1(n_1000),
.B2(n_997),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1078),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1059),
.A2(n_1010),
.B1(n_1012),
.B2(n_1007),
.Y(n_1387)
);

OA22x2_ASAP7_75t_L g1388 ( 
.A1(n_1059),
.A2(n_1017),
.B1(n_1052),
.B2(n_1013),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1059),
.A2(n_1034),
.B1(n_737),
.B2(n_743),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1170),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1059),
.A2(n_758),
.B1(n_786),
.B2(n_717),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1059),
.A2(n_813),
.B1(n_821),
.B2(n_818),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1176),
.A2(n_834),
.B1(n_846),
.B2(n_825),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1209),
.Y(n_1394)
);

XNOR2xp5_ASAP7_75t_L g1395 ( 
.A(n_1210),
.B(n_1196),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1217),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1204),
.B(n_879),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_SL g1398 ( 
.A(n_1283),
.B(n_637),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1227),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1314),
.Y(n_1400)
);

AND2x6_ASAP7_75t_L g1401 ( 
.A(n_1289),
.B(n_879),
.Y(n_1401)
);

INVx8_ASAP7_75t_L g1402 ( 
.A(n_1198),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1258),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1237),
.B(n_979),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1238),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1239),
.B(n_809),
.Y(n_1406)
);

INVxp33_ASAP7_75t_L g1407 ( 
.A(n_1194),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1183),
.B(n_867),
.Y(n_1408)
);

XNOR2x2_ASAP7_75t_L g1409 ( 
.A(n_1187),
.B(n_857),
.Y(n_1409)
);

XOR2x2_ASAP7_75t_L g1410 ( 
.A(n_1213),
.B(n_32),
.Y(n_1410)
);

XOR2xp5_ASAP7_75t_L g1411 ( 
.A(n_1208),
.B(n_32),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1229),
.Y(n_1412)
);

NAND2xp33_ASAP7_75t_R g1413 ( 
.A(n_1198),
.B(n_639),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1235),
.B(n_883),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1190),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1200),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1270),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1390),
.Y(n_1418)
);

XNOR2xp5_ASAP7_75t_L g1419 ( 
.A(n_1195),
.B(n_33),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1236),
.B(n_905),
.Y(n_1420)
);

AND2x6_ASAP7_75t_L g1421 ( 
.A(n_1290),
.B(n_1020),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1304),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1220),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1309),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1181),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1386),
.Y(n_1426)
);

INVxp33_ASAP7_75t_L g1427 ( 
.A(n_1329),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1284),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1285),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1186),
.B(n_1184),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1294),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1346),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1230),
.B(n_1247),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1301),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1375),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1282),
.B(n_909),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1375),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1230),
.B(n_685),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1262),
.B(n_33),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1247),
.B(n_686),
.Y(n_1440)
);

INVxp67_ASAP7_75t_L g1441 ( 
.A(n_1324),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1325),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1350),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1243),
.B(n_911),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1252),
.B(n_914),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1223),
.B(n_702),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1267),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1264),
.B(n_924),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1267),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1296),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1296),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1226),
.B(n_35),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1299),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1199),
.B(n_709),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1299),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1223),
.B(n_710),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1201),
.B(n_712),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1359),
.Y(n_1458)
);

XOR2xp5_ASAP7_75t_L g1459 ( 
.A(n_1207),
.B(n_35),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1324),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1338),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1219),
.B(n_713),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1362),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1187),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1338),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1219),
.B(n_719),
.Y(n_1466)
);

CKINVDCx14_ASAP7_75t_R g1467 ( 
.A(n_1252),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1341),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1271),
.A2(n_1260),
.B(n_1240),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1341),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1351),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1351),
.Y(n_1472)
);

INVxp33_ASAP7_75t_SL g1473 ( 
.A(n_1265),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1369),
.Y(n_1474)
);

CKINVDCx14_ASAP7_75t_R g1475 ( 
.A(n_1224),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1272),
.A2(n_940),
.B(n_935),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_SL g1477 ( 
.A(n_1310),
.B(n_729),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1369),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1218),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1311),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1311),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1379),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_R g1483 ( 
.A(n_1287),
.B(n_730),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1273),
.A2(n_1008),
.B(n_1006),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1214),
.B(n_1032),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1384),
.B(n_732),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1292),
.A2(n_932),
.B(n_739),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1364),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1211),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1211),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1191),
.B(n_1051),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1192),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1202),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1353),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_R g1495 ( 
.A(n_1274),
.B(n_735),
.Y(n_1495)
);

XOR2x2_ASAP7_75t_L g1496 ( 
.A(n_1266),
.B(n_36),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1355),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1372),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1357),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1379),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1244),
.Y(n_1501)
);

INVxp33_ASAP7_75t_SL g1502 ( 
.A(n_1385),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1212),
.B(n_1021),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1380),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1332),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1250),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1232),
.B(n_749),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1231),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1250),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1205),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1261),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1242),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1228),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1261),
.B(n_1019),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1205),
.B(n_759),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1345),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1234),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1206),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1206),
.B(n_1011),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1233),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1259),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1320),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1278),
.B(n_764),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1320),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_1316),
.B(n_1319),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1312),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1312),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1246),
.B(n_1009),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1317),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1317),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1193),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_R g1532 ( 
.A(n_1254),
.B(n_771),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_SL g1533 ( 
.A(n_1197),
.B(n_1004),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1322),
.Y(n_1534)
);

AND2x6_ASAP7_75t_L g1535 ( 
.A(n_1295),
.B(n_1297),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1280),
.B(n_778),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1248),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1249),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1193),
.B(n_966),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1322),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1245),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1378),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1288),
.B(n_783),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1179),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1188),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1293),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1251),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1373),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1255),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1331),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1330),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1279),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1241),
.B(n_36),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1306),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1343),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1203),
.B(n_792),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_SL g1557 ( 
.A(n_1257),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1348),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1354),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_SL g1560 ( 
.A(n_1257),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1298),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1326),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1334),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1286),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1333),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1225),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1221),
.B(n_37),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1277),
.B(n_794),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1257),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1335),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1318),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1370),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1377),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1363),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1263),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1328),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1368),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1180),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1389),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1388),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1276),
.B(n_957),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1339),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1307),
.B(n_795),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1340),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1393),
.B(n_951),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1349),
.Y(n_1586)
);

XNOR2xp5_ASAP7_75t_L g1587 ( 
.A(n_1253),
.B(n_38),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1366),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1269),
.B(n_802),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1315),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1268),
.B(n_1302),
.Y(n_1591)
);

AND2x2_ASAP7_75t_SL g1592 ( 
.A(n_1182),
.B(n_38),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1342),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1275),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1303),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1189),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1256),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1215),
.B(n_810),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1308),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1269),
.B(n_814),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1269),
.B(n_853),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1336),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1321),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1365),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1381),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1383),
.Y(n_1606)
);

INVxp33_ASAP7_75t_L g1607 ( 
.A(n_1216),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1281),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1300),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1291),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1391),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1185),
.B(n_945),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1392),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1305),
.B(n_865),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1337),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1358),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1387),
.B(n_943),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1352),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1367),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1347),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1222),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1313),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1327),
.B(n_39),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1356),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_R g1625 ( 
.A(n_1360),
.B(n_876),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1361),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1323),
.B(n_938),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1344),
.B(n_39),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1371),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1374),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_SL g1631 ( 
.A(n_1376),
.B(n_937),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1382),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1209),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1209),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1209),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1209),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1209),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1209),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1237),
.B(n_881),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1209),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1209),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1309),
.Y(n_1642)
);

XNOR2xp5_ASAP7_75t_L g1643 ( 
.A(n_1210),
.B(n_40),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1346),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1204),
.B(n_936),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1209),
.Y(n_1646)
);

NAND2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1184),
.B(n_889),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1209),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1204),
.B(n_894),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1209),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1209),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1209),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1209),
.Y(n_1653)
);

AOI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1240),
.A2(n_932),
.B(n_739),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1209),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1183),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1209),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1209),
.Y(n_1658)
);

XNOR2xp5_ASAP7_75t_L g1659 ( 
.A(n_1210),
.B(n_40),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1237),
.B(n_896),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1184),
.B(n_41),
.Y(n_1661)
);

XOR2xp5_ASAP7_75t_L g1662 ( 
.A(n_1196),
.B(n_42),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1209),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1237),
.B(n_902),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1209),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1190),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1209),
.Y(n_1667)
);

INVxp33_ASAP7_75t_SL g1668 ( 
.A(n_1195),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1209),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1271),
.A2(n_917),
.B(n_904),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1204),
.B(n_925),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1237),
.B(n_927),
.Y(n_1672)
);

XOR2xp5_ASAP7_75t_L g1673 ( 
.A(n_1196),
.B(n_42),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1258),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1209),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1209),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1209),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1258),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1209),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1214),
.B(n_928),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1209),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1209),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1209),
.Y(n_1683)
);

NAND2xp33_ASAP7_75t_R g1684 ( 
.A(n_1198),
.B(n_43),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1204),
.B(n_932),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1489),
.B(n_44),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1404),
.B(n_44),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1490),
.B(n_45),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1520),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1610),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1609),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1417),
.B(n_1510),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1406),
.B(n_45),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1424),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1398),
.B(n_739),
.Y(n_1695)
);

AND2x2_ASAP7_75t_SL g1696 ( 
.A(n_1540),
.B(n_46),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1417),
.B(n_739),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1546),
.B(n_739),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1546),
.B(n_739),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1511),
.B(n_739),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1639),
.B(n_932),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1476),
.A2(n_932),
.B(n_462),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1487),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1654),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1476),
.A2(n_932),
.B(n_464),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1639),
.B(n_932),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1424),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1394),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1518),
.B(n_46),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1396),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1633),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1416),
.Y(n_1712)
);

INVxp33_ASAP7_75t_L g1713 ( 
.A(n_1645),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1543),
.B(n_47),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1634),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1543),
.B(n_47),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1433),
.B(n_49),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1447),
.B(n_50),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1660),
.B(n_50),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1660),
.B(n_51),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1418),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1480),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1649),
.B(n_52),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1635),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1666),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1664),
.B(n_52),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1415),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1671),
.B(n_54),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_R g1729 ( 
.A(n_1467),
.B(n_55),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1438),
.B(n_55),
.Y(n_1730)
);

OR2x2_ASAP7_75t_SL g1731 ( 
.A(n_1452),
.B(n_1567),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1440),
.B(n_56),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1572),
.B(n_56),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1405),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1680),
.B(n_57),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1680),
.B(n_1430),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1636),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1664),
.B(n_57),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1611),
.B(n_58),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1637),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1638),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1613),
.B(n_58),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1480),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1444),
.A2(n_465),
.B(n_461),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1564),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1590),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1640),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1672),
.B(n_59),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1612),
.B(n_60),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1672),
.B(n_61),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_R g1751 ( 
.A(n_1413),
.B(n_61),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1397),
.B(n_62),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1425),
.B(n_62),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1508),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1426),
.B(n_63),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1424),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1641),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1646),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1492),
.B(n_63),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1449),
.B(n_64),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1446),
.B(n_65),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1493),
.B(n_66),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1441),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1456),
.B(n_66),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1398),
.B(n_1526),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1444),
.A2(n_467),
.B(n_466),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1512),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1500),
.B(n_67),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1412),
.B(n_67),
.Y(n_1769)
);

NOR2xp67_ASAP7_75t_L g1770 ( 
.A(n_1531),
.B(n_68),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1515),
.B(n_69),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1684),
.Y(n_1772)
);

BUFx3_ASAP7_75t_L g1773 ( 
.A(n_1481),
.Y(n_1773)
);

AND2x4_ASAP7_75t_SL g1774 ( 
.A(n_1445),
.B(n_70),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1441),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1661),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1648),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1537),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1500),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1519),
.B(n_71),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_R g1781 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1608),
.B(n_72),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1408),
.B(n_72),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1566),
.A2(n_471),
.B(n_469),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1511),
.B(n_73),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1685),
.B(n_73),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1484),
.A2(n_474),
.B(n_472),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1527),
.B(n_626),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_R g1789 ( 
.A(n_1464),
.B(n_74),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1650),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1482),
.Y(n_1791)
);

AND2x2_ASAP7_75t_SL g1792 ( 
.A(n_1460),
.B(n_74),
.Y(n_1792)
);

INVxp33_ASAP7_75t_L g1793 ( 
.A(n_1514),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1585),
.B(n_75),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1395),
.B(n_75),
.Y(n_1795)
);

AND2x2_ASAP7_75t_SL g1796 ( 
.A(n_1461),
.B(n_77),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1538),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1651),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1529),
.B(n_625),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1652),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1482),
.B(n_78),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1448),
.B(n_78),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1448),
.B(n_79),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1521),
.B(n_79),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1653),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1564),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1549),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1655),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1465),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1469),
.B(n_80),
.Y(n_1810)
);

AND2x2_ASAP7_75t_SL g1811 ( 
.A(n_1468),
.B(n_83),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1469),
.B(n_83),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1450),
.B(n_84),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1451),
.B(n_84),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1428),
.B(n_1429),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1462),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1466),
.B(n_85),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1657),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1431),
.B(n_85),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1503),
.B(n_86),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1599),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1658),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1663),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1618),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1434),
.B(n_86),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1470),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1665),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1603),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1402),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1471),
.B(n_475),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1593),
.B(n_88),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1486),
.B(n_89),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1582),
.B(n_89),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1642),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1457),
.B(n_1561),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1642),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1584),
.B(n_90),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1541),
.B(n_91),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1667),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1661),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1539),
.B(n_91),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1586),
.B(n_94),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1588),
.B(n_95),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1523),
.B(n_95),
.Y(n_1844)
);

NAND2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1472),
.B(n_1474),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1436),
.B(n_97),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1442),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1536),
.B(n_1581),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1669),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1675),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1676),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1568),
.B(n_97),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1677),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1642),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1478),
.Y(n_1855)
);

INVx3_ASAP7_75t_L g1856 ( 
.A(n_1443),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1435),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1522),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1656),
.B(n_98),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1607),
.B(n_98),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1679),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1597),
.B(n_99),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1402),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1621),
.B(n_99),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1436),
.B(n_100),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1617),
.B(n_1485),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1485),
.B(n_1579),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1458),
.Y(n_1868)
);

AND2x2_ASAP7_75t_SL g1869 ( 
.A(n_1437),
.B(n_101),
.Y(n_1869)
);

NOR2x1p5_ASAP7_75t_L g1870 ( 
.A(n_1674),
.B(n_101),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1681),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1605),
.B(n_102),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1606),
.B(n_1422),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1682),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1617),
.B(n_102),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1683),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1531),
.B(n_104),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1419),
.B(n_104),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1463),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1548),
.B(n_105),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1551),
.B(n_105),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1400),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1488),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1580),
.B(n_106),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1555),
.B(n_106),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1557),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1591),
.B(n_107),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1427),
.B(n_108),
.Y(n_1888)
);

INVx4_ASAP7_75t_L g1889 ( 
.A(n_1557),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1504),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1629),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1453),
.B(n_108),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1455),
.B(n_109),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1678),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1445),
.Y(n_1895)
);

NAND2xp33_ASAP7_75t_SL g1896 ( 
.A(n_1560),
.B(n_111),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1439),
.B(n_112),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1505),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1530),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1498),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1570),
.B(n_113),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1432),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1596),
.B(n_114),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1570),
.B(n_114),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_R g1905 ( 
.A(n_1495),
.B(n_1423),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1587),
.B(n_115),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1501),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1614),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1494),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1558),
.B(n_115),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1484),
.A2(n_479),
.B(n_476),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1445),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1497),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1499),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1569),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1506),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1630),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1509),
.B(n_116),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1644),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1644),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1507),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1643),
.B(n_117),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1399),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1659),
.B(n_117),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1594),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1407),
.B(n_1552),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1409),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1595),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1559),
.B(n_118),
.Y(n_1929)
);

INVx8_ASAP7_75t_L g1930 ( 
.A(n_1560),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1670),
.B(n_119),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1624),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1534),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1670),
.B(n_120),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1576),
.B(n_120),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1592),
.B(n_1575),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1626),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1614),
.B(n_121),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1507),
.B(n_1491),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1574),
.B(n_123),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1628),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1571),
.A2(n_481),
.B(n_480),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1491),
.B(n_124),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1632),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1578),
.B(n_124),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1535),
.B(n_125),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1577),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1550),
.B(n_125),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1535),
.B(n_126),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1459),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1411),
.B(n_127),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1550),
.B(n_127),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1615),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1662),
.B(n_128),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1553),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1622),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1562),
.A2(n_483),
.B(n_482),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1602),
.B(n_128),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1535),
.B(n_129),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1604),
.B(n_129),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1535),
.B(n_130),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1477),
.B(n_1525),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1553),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1524),
.Y(n_1964)
);

OAI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1565),
.A2(n_1573),
.B(n_1420),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1620),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1544),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1414),
.B(n_131),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1673),
.B(n_132),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1583),
.B(n_132),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1545),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1542),
.Y(n_1972)
);

OAI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1414),
.A2(n_486),
.B(n_484),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1547),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1420),
.B(n_133),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1421),
.B(n_133),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1528),
.B(n_134),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1421),
.B(n_1528),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1421),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1627),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1616),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1421),
.B(n_135),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1502),
.B(n_135),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1619),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1401),
.B(n_136),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1401),
.B(n_136),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1554),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1623),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1401),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1401),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1496),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1516),
.B(n_137),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1589),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1477),
.B(n_492),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1483),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1563),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1454),
.B(n_138),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1589),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1600),
.A2(n_496),
.B(n_493),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1600),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1601),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1516),
.B(n_1533),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1601),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1598),
.B(n_138),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1598),
.B(n_139),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1647),
.B(n_139),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1556),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1556),
.B(n_140),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1533),
.B(n_141),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1475),
.B(n_141),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1532),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1410),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1517),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1668),
.Y(n_2014)
);

INVx3_ASAP7_75t_L g2015 ( 
.A(n_1625),
.Y(n_2015)
);

OAI21xp5_ASAP7_75t_L g2016 ( 
.A1(n_1631),
.A2(n_501),
.B(n_500),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1513),
.Y(n_2017)
);

AND2x2_ASAP7_75t_SL g2018 ( 
.A(n_1631),
.B(n_142),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1473),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1479),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1424),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1404),
.B(n_142),
.Y(n_2022)
);

BUFx3_ASAP7_75t_L g2023 ( 
.A(n_1480),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_R g2024 ( 
.A(n_1467),
.B(n_143),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1609),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1572),
.B(n_145),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1736),
.B(n_145),
.Y(n_2027)
);

BUFx8_ASAP7_75t_L g2028 ( 
.A(n_1863),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1746),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1909),
.Y(n_2030)
);

NAND2x1_ASAP7_75t_L g2031 ( 
.A(n_1830),
.B(n_504),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1835),
.B(n_148),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1866),
.B(n_149),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1694),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1743),
.B(n_150),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1743),
.B(n_151),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1746),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1956),
.Y(n_2038)
);

OR2x6_ASAP7_75t_L g2039 ( 
.A(n_1930),
.B(n_151),
.Y(n_2039)
);

NAND2x1p5_ASAP7_75t_L g2040 ( 
.A(n_2023),
.B(n_153),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1694),
.Y(n_2041)
);

NAND2x1p5_ASAP7_75t_L g2042 ( 
.A(n_2023),
.B(n_154),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1913),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1956),
.Y(n_2044)
);

INVx5_ASAP7_75t_L g2045 ( 
.A(n_1694),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1914),
.B(n_154),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1815),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_1781),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1694),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1906),
.B(n_155),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1734),
.Y(n_2051)
);

NOR2xp67_ASAP7_75t_L g2052 ( 
.A(n_1895),
.B(n_155),
.Y(n_2052)
);

BUFx5_ASAP7_75t_L g2053 ( 
.A(n_1830),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1933),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1933),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_SL g2056 ( 
.A(n_1894),
.B(n_156),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1867),
.B(n_157),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1894),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1692),
.B(n_1689),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1707),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1734),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2013),
.B(n_158),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1692),
.B(n_158),
.Y(n_2063)
);

OR2x2_ASAP7_75t_L g2064 ( 
.A(n_1731),
.B(n_159),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1916),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1692),
.B(n_159),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_1795),
.B(n_161),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1691),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1921),
.B(n_162),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1776),
.B(n_162),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1947),
.B(n_163),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1916),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1707),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1773),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1983),
.B(n_164),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1707),
.Y(n_2076)
);

CKINVDCx20_ASAP7_75t_R g2077 ( 
.A(n_1781),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1819),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1983),
.B(n_1862),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2014),
.B(n_165),
.Y(n_2080)
);

NAND2x1_ASAP7_75t_L g2081 ( 
.A(n_1830),
.B(n_515),
.Y(n_2081)
);

NAND2x1_ASAP7_75t_L g2082 ( 
.A(n_1830),
.B(n_518),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1965),
.B(n_166),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1825),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1707),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1847),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1776),
.B(n_166),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1691),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1882),
.B(n_167),
.Y(n_2089)
);

BUFx4f_ASAP7_75t_L g2090 ( 
.A(n_1774),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2019),
.B(n_167),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1713),
.B(n_168),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1847),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2025),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2025),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1783),
.B(n_168),
.Y(n_2096)
);

OR2x6_ASAP7_75t_L g2097 ( 
.A(n_1930),
.B(n_1912),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1868),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1864),
.B(n_170),
.Y(n_2099)
);

NAND2x1_ASAP7_75t_L g2100 ( 
.A(n_1830),
.B(n_519),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_1898),
.Y(n_2101)
);

HB1xp67_ASAP7_75t_L g2102 ( 
.A(n_1891),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1868),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_1935),
.Y(n_2104)
);

NOR2x1_ASAP7_75t_SL g2105 ( 
.A(n_1810),
.B(n_170),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_1773),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_1840),
.B(n_171),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1897),
.B(n_172),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_2021),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_2021),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_1840),
.B(n_173),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1878),
.B(n_1848),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1809),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_2021),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1722),
.B(n_173),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1810),
.B(n_174),
.Y(n_2116)
);

OR2x2_ASAP7_75t_L g2117 ( 
.A(n_2017),
.B(n_174),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1908),
.B(n_175),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1722),
.B(n_175),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_1935),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_1791),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1900),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1812),
.B(n_176),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1809),
.Y(n_2124)
);

NAND2x1p5_ASAP7_75t_L g2125 ( 
.A(n_1756),
.B(n_178),
.Y(n_2125)
);

HB1xp67_ASAP7_75t_L g2126 ( 
.A(n_1774),
.Y(n_2126)
);

OR2x6_ASAP7_75t_L g2127 ( 
.A(n_1930),
.B(n_1886),
.Y(n_2127)
);

BUFx6f_ASAP7_75t_L g2128 ( 
.A(n_2021),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1756),
.Y(n_2129)
);

NAND2x1p5_ASAP7_75t_L g2130 ( 
.A(n_1756),
.B(n_1834),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1955),
.B(n_1886),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1812),
.B(n_178),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_1834),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1900),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_SL g2135 ( 
.A(n_1895),
.B(n_179),
.Y(n_2135)
);

AND2x6_ASAP7_75t_L g2136 ( 
.A(n_1718),
.B(n_179),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1829),
.Y(n_2137)
);

INVx6_ASAP7_75t_L g2138 ( 
.A(n_1886),
.Y(n_2138)
);

NOR2x1_ASAP7_75t_L g2139 ( 
.A(n_1889),
.B(n_180),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2017),
.B(n_180),
.Y(n_2140)
);

AND2x6_ASAP7_75t_L g2141 ( 
.A(n_1718),
.B(n_181),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1687),
.B(n_181),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1889),
.B(n_182),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1836),
.Y(n_2144)
);

AND2x2_ASAP7_75t_SL g2145 ( 
.A(n_1696),
.B(n_183),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_1763),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1917),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1889),
.B(n_184),
.Y(n_2148)
);

INVx4_ASAP7_75t_L g2149 ( 
.A(n_1829),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1693),
.B(n_185),
.Y(n_2150)
);

NAND2x1p5_ASAP7_75t_L g2151 ( 
.A(n_1836),
.B(n_185),
.Y(n_2151)
);

CKINVDCx8_ASAP7_75t_R g2152 ( 
.A(n_1930),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2022),
.B(n_186),
.Y(n_2153)
);

INVxp67_ASAP7_75t_L g2154 ( 
.A(n_1935),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1824),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1922),
.B(n_187),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_1950),
.B(n_187),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1883),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_1950),
.B(n_190),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1713),
.B(n_190),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1854),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_2018),
.B(n_191),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1963),
.B(n_192),
.Y(n_2163)
);

INVx5_ASAP7_75t_L g2164 ( 
.A(n_1985),
.Y(n_2164)
);

INVx2_ASAP7_75t_SL g2165 ( 
.A(n_1824),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_1854),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1709),
.Y(n_2167)
);

AND2x4_ASAP7_75t_L g2168 ( 
.A(n_1963),
.B(n_192),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_SL g2169 ( 
.A(n_2018),
.B(n_193),
.Y(n_2169)
);

CKINVDCx6p67_ASAP7_75t_R g2170 ( 
.A(n_1995),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1854),
.Y(n_2171)
);

INVx5_ASAP7_75t_L g2172 ( 
.A(n_1985),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1907),
.B(n_194),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2020),
.B(n_194),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_1967),
.B(n_196),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1709),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1890),
.B(n_198),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1883),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1751),
.B(n_198),
.Y(n_2179)
);

NAND2x1_ASAP7_75t_SL g2180 ( 
.A(n_1985),
.B(n_199),
.Y(n_2180)
);

NAND2x1_ASAP7_75t_SL g2181 ( 
.A(n_1990),
.B(n_199),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1987),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1917),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1924),
.B(n_200),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_SL g2185 ( 
.A(n_1696),
.B(n_200),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1735),
.B(n_201),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1709),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_1967),
.B(n_202),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1727),
.Y(n_2189)
);

BUFx3_ASAP7_75t_L g2190 ( 
.A(n_1856),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_1729),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_1971),
.B(n_202),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1708),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1718),
.Y(n_2194)
);

NAND2x1p5_ASAP7_75t_L g2195 ( 
.A(n_1979),
.B(n_203),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1793),
.B(n_203),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1842),
.B(n_204),
.Y(n_2197)
);

BUFx6f_ASAP7_75t_L g2198 ( 
.A(n_1760),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_SL g2199 ( 
.A(n_1792),
.B(n_204),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_1971),
.B(n_205),
.Y(n_2200)
);

INVx5_ASAP7_75t_L g2201 ( 
.A(n_1760),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_SL g2202 ( 
.A(n_1792),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_1974),
.B(n_206),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1760),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_SL g2205 ( 
.A(n_1796),
.B(n_207),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_1775),
.Y(n_2206)
);

BUFx6f_ASAP7_75t_L g2207 ( 
.A(n_1814),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2010),
.B(n_209),
.Y(n_2208)
);

INVxp67_ASAP7_75t_L g2209 ( 
.A(n_1958),
.Y(n_2209)
);

AO21x2_ASAP7_75t_L g2210 ( 
.A1(n_1765),
.A2(n_523),
.B(n_522),
.Y(n_2210)
);

NAND2x1p5_ASAP7_75t_L g2211 ( 
.A(n_1979),
.B(n_210),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_1729),
.Y(n_2212)
);

OR2x6_ASAP7_75t_L g2213 ( 
.A(n_1772),
.B(n_210),
.Y(n_2213)
);

OR2x6_ASAP7_75t_L g2214 ( 
.A(n_1870),
.B(n_211),
.Y(n_2214)
);

NAND2x1_ASAP7_75t_SL g2215 ( 
.A(n_1990),
.B(n_211),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1842),
.B(n_212),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1793),
.B(n_212),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1710),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1711),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_1751),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2010),
.B(n_213),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1939),
.B(n_213),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1844),
.B(n_214),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_1926),
.B(n_214),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1814),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1814),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1892),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_1794),
.B(n_215),
.Y(n_2228)
);

AND2x6_ASAP7_75t_L g2229 ( 
.A(n_1892),
.B(n_1893),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1892),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1852),
.B(n_215),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1816),
.B(n_217),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1715),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1727),
.Y(n_2234)
);

AND2x4_ASAP7_75t_L g2235 ( 
.A(n_1974),
.B(n_217),
.Y(n_2235)
);

BUFx2_ASAP7_75t_SL g2236 ( 
.A(n_1893),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_1779),
.Y(n_2237)
);

NAND2x1p5_ASAP7_75t_L g2238 ( 
.A(n_1893),
.B(n_218),
.Y(n_2238)
);

BUFx5_ASAP7_75t_L g2239 ( 
.A(n_1920),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_1899),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1932),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1724),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_1981),
.B(n_1984),
.Y(n_2243)
);

AND2x6_ASAP7_75t_L g2244 ( 
.A(n_1686),
.B(n_1688),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1856),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1826),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1932),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_1936),
.B(n_218),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1737),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1951),
.B(n_220),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_1920),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_1991),
.B(n_220),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1972),
.B(n_222),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1937),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_SL g2255 ( 
.A(n_1796),
.B(n_222),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1954),
.B(n_223),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1740),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_1899),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1741),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1820),
.B(n_224),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1826),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_1980),
.B(n_1858),
.Y(n_2262)
);

CKINVDCx6p67_ASAP7_75t_R g2263 ( 
.A(n_1958),
.Y(n_2263)
);

BUFx6f_ASAP7_75t_L g2264 ( 
.A(n_1899),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_SL g2265 ( 
.A(n_1811),
.B(n_1768),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1855),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1937),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2012),
.B(n_224),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1969),
.B(n_225),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1832),
.B(n_225),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2012),
.B(n_226),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_1858),
.B(n_226),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1723),
.B(n_227),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1728),
.B(n_227),
.Y(n_2274)
);

BUFx5_ASAP7_75t_L g2275 ( 
.A(n_1989),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_1856),
.B(n_1879),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1855),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_2024),
.Y(n_2278)
);

OR2x6_ASAP7_75t_L g2279 ( 
.A(n_1958),
.B(n_228),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_1768),
.B(n_229),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1779),
.B(n_230),
.Y(n_2281)
);

BUFx4f_ASAP7_75t_L g2282 ( 
.A(n_1811),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_1879),
.B(n_1859),
.Y(n_2283)
);

BUFx2_ASAP7_75t_L g2284 ( 
.A(n_2024),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_1686),
.B(n_231),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1754),
.Y(n_2286)
);

INVx4_ASAP7_75t_L g2287 ( 
.A(n_1918),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1875),
.B(n_232),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_1879),
.B(n_232),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1739),
.B(n_233),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_1925),
.B(n_233),
.Y(n_2291)
);

BUFx3_ASAP7_75t_L g2292 ( 
.A(n_1960),
.Y(n_2292)
);

OR2x6_ASAP7_75t_L g2293 ( 
.A(n_1960),
.B(n_234),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_1972),
.B(n_234),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_SL g2295 ( 
.A(n_1869),
.B(n_235),
.Y(n_2295)
);

BUFx2_ASAP7_75t_L g2296 ( 
.A(n_1905),
.Y(n_2296)
);

INVx5_ASAP7_75t_L g2297 ( 
.A(n_1918),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1905),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1742),
.B(n_235),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_1928),
.B(n_236),
.Y(n_2300)
);

BUFx24_ASAP7_75t_SL g2301 ( 
.A(n_1996),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1945),
.B(n_236),
.Y(n_2302)
);

INVx8_ASAP7_75t_L g2303 ( 
.A(n_1960),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_SL g2304 ( 
.A(n_1869),
.B(n_237),
.Y(n_2304)
);

INVx6_ASAP7_75t_L g2305 ( 
.A(n_2026),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_1992),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_1747),
.B(n_1757),
.Y(n_2307)
);

AND2x4_ASAP7_75t_L g2308 ( 
.A(n_1758),
.B(n_1777),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1749),
.B(n_237),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1754),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1857),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_1790),
.B(n_239),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1752),
.B(n_1798),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_1978),
.B(n_239),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1767),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1800),
.B(n_240),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_1996),
.Y(n_2317)
);

INVx4_ASAP7_75t_L g2318 ( 
.A(n_1918),
.Y(n_2318)
);

BUFx4f_ASAP7_75t_L g2319 ( 
.A(n_1686),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2011),
.B(n_241),
.Y(n_2320)
);

NAND2x1p5_ASAP7_75t_L g2321 ( 
.A(n_1688),
.B(n_2015),
.Y(n_2321)
);

INVx4_ASAP7_75t_L g2322 ( 
.A(n_1688),
.Y(n_2322)
);

OR2x6_ASAP7_75t_L g2323 ( 
.A(n_2011),
.B(n_241),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1857),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1712),
.Y(n_2325)
);

INVx6_ASAP7_75t_L g2326 ( 
.A(n_1888),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_SL g2327 ( 
.A(n_2009),
.B(n_242),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_1992),
.Y(n_2328)
);

NAND2x1p5_ASAP7_75t_L g2329 ( 
.A(n_2015),
.B(n_242),
.Y(n_2329)
);

OR2x6_ASAP7_75t_L g2330 ( 
.A(n_2009),
.B(n_243),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_1805),
.B(n_244),
.Y(n_2331)
);

OR2x6_ASAP7_75t_L g2332 ( 
.A(n_2015),
.B(n_246),
.Y(n_2332)
);

CKINVDCx11_ASAP7_75t_R g2333 ( 
.A(n_1992),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2007),
.B(n_246),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1712),
.Y(n_2335)
);

BUFx2_ASAP7_75t_L g2336 ( 
.A(n_1801),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1767),
.Y(n_2337)
);

BUFx4f_ASAP7_75t_L g2338 ( 
.A(n_1990),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1721),
.Y(n_2339)
);

INVxp67_ASAP7_75t_L g2340 ( 
.A(n_1789),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2007),
.B(n_247),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_1761),
.B(n_248),
.Y(n_2342)
);

AND2x2_ASAP7_75t_SL g2343 ( 
.A(n_1801),
.B(n_1927),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_1808),
.B(n_248),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1818),
.B(n_249),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1822),
.B(n_250),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_1823),
.B(n_251),
.Y(n_2347)
);

INVxp67_ASAP7_75t_L g2348 ( 
.A(n_1860),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1721),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_SL g2350 ( 
.A(n_1964),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_1785),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_SL g2352 ( 
.A(n_1838),
.B(n_251),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1827),
.B(n_252),
.Y(n_2353)
);

NAND2x1p5_ASAP7_75t_L g2354 ( 
.A(n_1785),
.B(n_254),
.Y(n_2354)
);

INVx6_ASAP7_75t_L g2355 ( 
.A(n_1782),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1725),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_1839),
.B(n_255),
.Y(n_2357)
);

NOR2xp67_ASAP7_75t_L g2358 ( 
.A(n_1838),
.B(n_256),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_1899),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_1849),
.B(n_256),
.Y(n_2360)
);

INVx1_ASAP7_75t_SL g2361 ( 
.A(n_1717),
.Y(n_2361)
);

BUFx3_ASAP7_75t_L g2362 ( 
.A(n_1690),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1850),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_1730),
.B(n_257),
.Y(n_2364)
);

AND2x4_ASAP7_75t_L g2365 ( 
.A(n_1851),
.B(n_258),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_SL g2366 ( 
.A(n_2016),
.B(n_258),
.Y(n_2366)
);

INVx4_ASAP7_75t_L g2367 ( 
.A(n_1745),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2003),
.Y(n_2368)
);

NOR2x1_ASAP7_75t_SL g2369 ( 
.A(n_1962),
.B(n_259),
.Y(n_2369)
);

OR2x6_ASAP7_75t_L g2370 ( 
.A(n_1764),
.B(n_260),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_1860),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1732),
.B(n_260),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1778),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_1873),
.B(n_261),
.Y(n_2374)
);

CKINVDCx14_ASAP7_75t_R g2375 ( 
.A(n_1896),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1853),
.Y(n_2376)
);

NAND2x1p5_ASAP7_75t_L g2377 ( 
.A(n_1745),
.B(n_261),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_1938),
.B(n_262),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1861),
.Y(n_2379)
);

OR2x2_ASAP7_75t_L g2380 ( 
.A(n_1902),
.B(n_262),
.Y(n_2380)
);

INVx4_ASAP7_75t_L g2381 ( 
.A(n_1745),
.Y(n_2381)
);

BUFx2_ASAP7_75t_L g2382 ( 
.A(n_1896),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1871),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_SL g2384 ( 
.A(n_1931),
.B(n_263),
.Y(n_2384)
);

HB1xp67_ASAP7_75t_L g2385 ( 
.A(n_1698),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1874),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1876),
.B(n_1993),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_1998),
.B(n_264),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1813),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2000),
.B(n_265),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_1923),
.B(n_265),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1813),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1817),
.B(n_267),
.Y(n_2393)
);

INVx5_ASAP7_75t_L g2394 ( 
.A(n_2003),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_1975),
.B(n_268),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_1975),
.B(n_268),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_1919),
.B(n_269),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_SL g2398 ( 
.A(n_1988),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1753),
.Y(n_2399)
);

INVx6_ASAP7_75t_L g2400 ( 
.A(n_1901),
.Y(n_2400)
);

INVx2_ASAP7_75t_SL g2401 ( 
.A(n_1877),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1755),
.Y(n_2402)
);

OR2x2_ASAP7_75t_L g2403 ( 
.A(n_1771),
.B(n_269),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_1780),
.B(n_270),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_SL g2405 ( 
.A(n_2002),
.B(n_270),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_1806),
.B(n_274),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_1700),
.B(n_2001),
.Y(n_2407)
);

NAND2x1_ASAP7_75t_L g2408 ( 
.A(n_1915),
.B(n_524),
.Y(n_2408)
);

CKINVDCx6p67_ASAP7_75t_R g2409 ( 
.A(n_1733),
.Y(n_2409)
);

NOR2x1_ASAP7_75t_L g2410 ( 
.A(n_1986),
.B(n_275),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_1884),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_1977),
.B(n_275),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_1904),
.B(n_276),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_1700),
.B(n_276),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_2003),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_1841),
.B(n_277),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_1759),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_1940),
.B(n_277),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2001),
.B(n_278),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_1690),
.B(n_278),
.Y(n_2420)
);

BUFx8_ASAP7_75t_L g2421 ( 
.A(n_2002),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1778),
.Y(n_2422)
);

BUFx12f_ASAP7_75t_L g2423 ( 
.A(n_1903),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1977),
.B(n_279),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1762),
.Y(n_2425)
);

INVx2_ASAP7_75t_SL g2426 ( 
.A(n_1690),
.Y(n_2426)
);

INVx5_ASAP7_75t_L g2427 ( 
.A(n_2003),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_1966),
.B(n_280),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_1946),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_1698),
.B(n_280),
.Y(n_2430)
);

NAND2x1p5_ASAP7_75t_L g2431 ( 
.A(n_1806),
.B(n_281),
.Y(n_2431)
);

OR2x6_ASAP7_75t_L g2432 ( 
.A(n_1949),
.B(n_281),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_1797),
.Y(n_2433)
);

INVx3_ASAP7_75t_L g2434 ( 
.A(n_1806),
.Y(n_2434)
);

BUFx12f_ASAP7_75t_L g2435 ( 
.A(n_1699),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_1725),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_1699),
.Y(n_2437)
);

BUFx2_ASAP7_75t_L g2438 ( 
.A(n_1941),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_1915),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1833),
.B(n_283),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_1887),
.B(n_283),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_1966),
.B(n_284),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1837),
.B(n_285),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1797),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_1959),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_1843),
.B(n_285),
.Y(n_2446)
);

OR2x2_ASAP7_75t_L g2447 ( 
.A(n_1846),
.B(n_286),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_1962),
.B(n_287),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_1941),
.B(n_287),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_1941),
.B(n_291),
.Y(n_2450)
);

AND2x4_ASAP7_75t_L g2451 ( 
.A(n_1804),
.B(n_291),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_1769),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1865),
.B(n_292),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_1807),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_SL g2455 ( 
.A(n_1787),
.B(n_292),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_1807),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1821),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1802),
.B(n_1803),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_1770),
.B(n_294),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_SL g2460 ( 
.A(n_1911),
.B(n_294),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_1976),
.Y(n_2461)
);

INVxp67_ASAP7_75t_L g2462 ( 
.A(n_1887),
.Y(n_2462)
);

AND2x4_ASAP7_75t_L g2463 ( 
.A(n_1915),
.B(n_295),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_1821),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_SL g2465 ( 
.A(n_1961),
.B(n_296),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_2229),
.Y(n_2466)
);

CKINVDCx20_ASAP7_75t_R g2467 ( 
.A(n_2077),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2047),
.Y(n_2468)
);

INVx8_ASAP7_75t_L g2469 ( 
.A(n_2303),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2030),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2034),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2028),
.Y(n_2472)
);

INVx6_ASAP7_75t_L g2473 ( 
.A(n_2028),
.Y(n_2473)
);

NAND2x1p5_ASAP7_75t_L g2474 ( 
.A(n_2319),
.B(n_1828),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2029),
.Y(n_2475)
);

AOI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2229),
.A2(n_1952),
.B1(n_1948),
.B2(n_1970),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2034),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2074),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2043),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2037),
.Y(n_2480)
);

BUFx12f_ASAP7_75t_L g2481 ( 
.A(n_2039),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2193),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2147),
.Y(n_2483)
);

INVx3_ASAP7_75t_L g2484 ( 
.A(n_2229),
.Y(n_2484)
);

CKINVDCx14_ASAP7_75t_R g2485 ( 
.A(n_2090),
.Y(n_2485)
);

BUFx4f_ASAP7_75t_SL g2486 ( 
.A(n_2263),
.Y(n_2486)
);

BUFx2_ASAP7_75t_SL g2487 ( 
.A(n_2152),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2106),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2183),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2218),
.Y(n_2490)
);

INVxp67_ASAP7_75t_SL g2491 ( 
.A(n_2319),
.Y(n_2491)
);

INVx4_ASAP7_75t_L g2492 ( 
.A(n_2090),
.Y(n_2492)
);

BUFx3_ASAP7_75t_L g2493 ( 
.A(n_2137),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2219),
.Y(n_2494)
);

INVx3_ASAP7_75t_SL g2495 ( 
.A(n_2039),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2229),
.B(n_1934),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2325),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2233),
.Y(n_2498)
);

BUFx12f_ASAP7_75t_L g2499 ( 
.A(n_2298),
.Y(n_2499)
);

AND2x6_ASAP7_75t_L g2500 ( 
.A(n_2167),
.B(n_1948),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2244),
.Y(n_2501)
);

BUFx2_ASAP7_75t_SL g2502 ( 
.A(n_2149),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_2101),
.Y(n_2503)
);

BUFx12f_ASAP7_75t_L g2504 ( 
.A(n_2317),
.Y(n_2504)
);

INVx6_ASAP7_75t_SL g2505 ( 
.A(n_2127),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2034),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2041),
.Y(n_2507)
);

INVx1_ASAP7_75t_SL g2508 ( 
.A(n_2236),
.Y(n_2508)
);

INVx1_ASAP7_75t_SL g2509 ( 
.A(n_2236),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2244),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2145),
.B(n_1952),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2242),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2041),
.Y(n_2513)
);

INVx8_ASAP7_75t_L g2514 ( 
.A(n_2303),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2170),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2249),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2244),
.Y(n_2517)
);

BUFx3_ASAP7_75t_L g2518 ( 
.A(n_2155),
.Y(n_2518)
);

BUFx3_ASAP7_75t_L g2519 ( 
.A(n_2048),
.Y(n_2519)
);

BUFx2_ASAP7_75t_L g2520 ( 
.A(n_2244),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2112),
.B(n_2079),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2041),
.Y(n_2522)
);

INVx5_ASAP7_75t_L g2523 ( 
.A(n_2136),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2389),
.B(n_1880),
.Y(n_2524)
);

INVx5_ASAP7_75t_L g2525 ( 
.A(n_2136),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2257),
.Y(n_2526)
);

BUFx2_ASAP7_75t_L g2527 ( 
.A(n_2435),
.Y(n_2527)
);

INVx5_ASAP7_75t_L g2528 ( 
.A(n_2136),
.Y(n_2528)
);

INVx8_ASAP7_75t_L g2529 ( 
.A(n_2279),
.Y(n_2529)
);

INVx4_ASAP7_75t_L g2530 ( 
.A(n_2045),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2287),
.Y(n_2531)
);

INVx3_ASAP7_75t_SL g2532 ( 
.A(n_2097),
.Y(n_2532)
);

BUFx5_ASAP7_75t_L g2533 ( 
.A(n_2325),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2138),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2259),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2343),
.B(n_1970),
.Y(n_2536)
);

BUFx2_ASAP7_75t_SL g2537 ( 
.A(n_2149),
.Y(n_2537)
);

INVx4_ASAP7_75t_L g2538 ( 
.A(n_2045),
.Y(n_2538)
);

BUFx2_ASAP7_75t_SL g2539 ( 
.A(n_2163),
.Y(n_2539)
);

INVx4_ASAP7_75t_L g2540 ( 
.A(n_2045),
.Y(n_2540)
);

INVx5_ASAP7_75t_L g2541 ( 
.A(n_2136),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2035),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2278),
.Y(n_2543)
);

INVx5_ASAP7_75t_SL g2544 ( 
.A(n_2127),
.Y(n_2544)
);

BUFx3_ASAP7_75t_L g2545 ( 
.A(n_2182),
.Y(n_2545)
);

BUFx6f_ASAP7_75t_L g2546 ( 
.A(n_2049),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_2131),
.Y(n_2547)
);

NAND2x1p5_ASAP7_75t_L g2548 ( 
.A(n_2201),
.B(n_1828),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_SL g2549 ( 
.A(n_2214),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2035),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2392),
.B(n_1881),
.Y(n_2551)
);

BUFx6f_ASAP7_75t_L g2552 ( 
.A(n_2049),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2363),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2376),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2279),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2462),
.B(n_1885),
.Y(n_2556)
);

BUFx12f_ASAP7_75t_L g2557 ( 
.A(n_2333),
.Y(n_2557)
);

BUFx2_ASAP7_75t_L g2558 ( 
.A(n_2293),
.Y(n_2558)
);

BUFx3_ASAP7_75t_L g2559 ( 
.A(n_2131),
.Y(n_2559)
);

NAND2x1p5_ASAP7_75t_L g2560 ( 
.A(n_2201),
.B(n_1944),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2049),
.Y(n_2561)
);

BUFx4f_ASAP7_75t_SL g2562 ( 
.A(n_2141),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2379),
.Y(n_2563)
);

INVx2_ASAP7_75t_SL g2564 ( 
.A(n_2138),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2383),
.Y(n_2565)
);

NAND2x1p5_ASAP7_75t_L g2566 ( 
.A(n_2201),
.B(n_1944),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2386),
.Y(n_2567)
);

INVx5_ASAP7_75t_L g2568 ( 
.A(n_2141),
.Y(n_2568)
);

NAND2x1p5_ASAP7_75t_L g2569 ( 
.A(n_2297),
.B(n_1994),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2335),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2282),
.B(n_1982),
.Y(n_2571)
);

NAND2x1p5_ASAP7_75t_L g2572 ( 
.A(n_2297),
.B(n_1994),
.Y(n_2572)
);

BUFx2_ASAP7_75t_L g2573 ( 
.A(n_2293),
.Y(n_2573)
);

CKINVDCx20_ASAP7_75t_R g2574 ( 
.A(n_2284),
.Y(n_2574)
);

AO21x2_ASAP7_75t_L g2575 ( 
.A1(n_2334),
.A2(n_1705),
.B(n_1702),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_2141),
.Y(n_2576)
);

HB1xp67_ASAP7_75t_L g2577 ( 
.A(n_2297),
.Y(n_2577)
);

BUFx8_ASAP7_75t_L g2578 ( 
.A(n_2350),
.Y(n_2578)
);

INVx4_ASAP7_75t_L g2579 ( 
.A(n_2141),
.Y(n_2579)
);

INVx4_ASAP7_75t_L g2580 ( 
.A(n_2164),
.Y(n_2580)
);

BUFx2_ASAP7_75t_L g2581 ( 
.A(n_2126),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2335),
.Y(n_2582)
);

BUFx4f_ASAP7_75t_SL g2583 ( 
.A(n_2163),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2272),
.Y(n_2584)
);

INVx1_ASAP7_75t_SL g2585 ( 
.A(n_2036),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2387),
.B(n_1910),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2097),
.Y(n_2587)
);

INVx5_ASAP7_75t_L g2588 ( 
.A(n_2076),
.Y(n_2588)
);

BUFx6f_ASAP7_75t_L g2589 ( 
.A(n_2076),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2272),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2121),
.Y(n_2591)
);

BUFx12f_ASAP7_75t_L g2592 ( 
.A(n_2296),
.Y(n_2592)
);

BUFx12f_ASAP7_75t_L g2593 ( 
.A(n_2214),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2282),
.B(n_1697),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2117),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2140),
.Y(n_2596)
);

INVx2_ASAP7_75t_SL g2597 ( 
.A(n_2036),
.Y(n_2597)
);

BUFx12f_ASAP7_75t_L g2598 ( 
.A(n_2191),
.Y(n_2598)
);

BUFx3_ASAP7_75t_L g2599 ( 
.A(n_2168),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2168),
.Y(n_2600)
);

INVx2_ASAP7_75t_SL g2601 ( 
.A(n_2165),
.Y(n_2601)
);

INVx1_ASAP7_75t_SL g2602 ( 
.A(n_2167),
.Y(n_2602)
);

CKINVDCx20_ASAP7_75t_R g2603 ( 
.A(n_2058),
.Y(n_2603)
);

BUFx12f_ASAP7_75t_L g2604 ( 
.A(n_2212),
.Y(n_2604)
);

BUFx2_ASAP7_75t_SL g2605 ( 
.A(n_2202),
.Y(n_2605)
);

BUFx3_ASAP7_75t_L g2606 ( 
.A(n_2130),
.Y(n_2606)
);

BUFx12f_ASAP7_75t_L g2607 ( 
.A(n_2143),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2385),
.B(n_1929),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2287),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2336),
.B(n_1872),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2070),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2070),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2076),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2087),
.Y(n_2614)
);

BUFx2_ASAP7_75t_R g2615 ( 
.A(n_2301),
.Y(n_2615)
);

BUFx12f_ASAP7_75t_L g2616 ( 
.A(n_2143),
.Y(n_2616)
);

CKINVDCx16_ASAP7_75t_R g2617 ( 
.A(n_2135),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2087),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2339),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2107),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2085),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2107),
.Y(n_2622)
);

BUFx3_ASAP7_75t_L g2623 ( 
.A(n_2220),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2318),
.B(n_2322),
.Y(n_2624)
);

INVx4_ASAP7_75t_L g2625 ( 
.A(n_2164),
.Y(n_2625)
);

BUFx4_ASAP7_75t_SL g2626 ( 
.A(n_2330),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2111),
.Y(n_2627)
);

AOI22xp33_ASAP7_75t_L g2628 ( 
.A1(n_2202),
.A2(n_1831),
.B1(n_1716),
.B2(n_1714),
.Y(n_2628)
);

BUFx2_ASAP7_75t_SL g2629 ( 
.A(n_2164),
.Y(n_2629)
);

INVx6_ASAP7_75t_L g2630 ( 
.A(n_2421),
.Y(n_2630)
);

INVx5_ASAP7_75t_SL g2631 ( 
.A(n_2330),
.Y(n_2631)
);

INVx1_ASAP7_75t_SL g2632 ( 
.A(n_2167),
.Y(n_2632)
);

CKINVDCx20_ASAP7_75t_R g2633 ( 
.A(n_2375),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2102),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2085),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_L g2636 ( 
.A(n_2361),
.B(n_1719),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2111),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2312),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2262),
.Y(n_2639)
);

INVx5_ASAP7_75t_L g2640 ( 
.A(n_2085),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2312),
.Y(n_2641)
);

BUFx3_ASAP7_75t_L g2642 ( 
.A(n_2129),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_2109),
.Y(n_2643)
);

NAND2x1p5_ASAP7_75t_L g2644 ( 
.A(n_2318),
.B(n_2322),
.Y(n_2644)
);

INVx3_ASAP7_75t_L g2645 ( 
.A(n_2129),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2347),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2339),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2347),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2357),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2292),
.B(n_2006),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2172),
.B(n_1720),
.Y(n_2651)
);

CKINVDCx16_ASAP7_75t_R g2652 ( 
.A(n_2056),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2176),
.Y(n_2653)
);

INVx4_ASAP7_75t_L g2654 ( 
.A(n_2172),
.Y(n_2654)
);

BUFx10_ASAP7_75t_L g2655 ( 
.A(n_2148),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2394),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2357),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2360),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2360),
.Y(n_2659)
);

INVx6_ASAP7_75t_L g2660 ( 
.A(n_2421),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_2348),
.B(n_1726),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2176),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2365),
.Y(n_2663)
);

INVxp67_ASAP7_75t_SL g2664 ( 
.A(n_2175),
.Y(n_2664)
);

INVx4_ASAP7_75t_L g2665 ( 
.A(n_2172),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2349),
.Y(n_2666)
);

INVx8_ASAP7_75t_L g2667 ( 
.A(n_2332),
.Y(n_2667)
);

INVx6_ASAP7_75t_L g2668 ( 
.A(n_2243),
.Y(n_2668)
);

INVx3_ASAP7_75t_SL g2669 ( 
.A(n_2323),
.Y(n_2669)
);

BUFx12f_ASAP7_75t_L g2670 ( 
.A(n_2148),
.Y(n_2670)
);

BUFx3_ASAP7_75t_L g2671 ( 
.A(n_2394),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2349),
.Y(n_2672)
);

INVx1_ASAP7_75t_SL g2673 ( 
.A(n_2176),
.Y(n_2673)
);

BUFx6f_ASAP7_75t_L g2674 ( 
.A(n_2109),
.Y(n_2674)
);

BUFx3_ASAP7_75t_L g2675 ( 
.A(n_2394),
.Y(n_2675)
);

INVx4_ASAP7_75t_L g2676 ( 
.A(n_2427),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2033),
.B(n_1738),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2356),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2187),
.Y(n_2679)
);

INVx1_ASAP7_75t_SL g2680 ( 
.A(n_2187),
.Y(n_2680)
);

AND2x4_ASAP7_75t_L g2681 ( 
.A(n_2307),
.B(n_1748),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2208),
.B(n_1750),
.Y(n_2682)
);

INVx3_ASAP7_75t_SL g2683 ( 
.A(n_2323),
.Y(n_2683)
);

BUFx6f_ASAP7_75t_SL g2684 ( 
.A(n_2213),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2365),
.Y(n_2685)
);

NAND2x1p5_ASAP7_75t_L g2686 ( 
.A(n_2187),
.B(n_1765),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_2213),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2356),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2427),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2262),
.Y(n_2690)
);

INVx4_ASAP7_75t_L g2691 ( 
.A(n_2427),
.Y(n_2691)
);

BUFx3_ASAP7_75t_L g2692 ( 
.A(n_2289),
.Y(n_2692)
);

BUFx3_ASAP7_75t_L g2693 ( 
.A(n_2289),
.Y(n_2693)
);

BUFx12f_ASAP7_75t_L g2694 ( 
.A(n_2332),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2109),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2291),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2146),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2350),
.Y(n_2698)
);

BUFx6f_ASAP7_75t_L g2699 ( 
.A(n_2110),
.Y(n_2699)
);

CKINVDCx5p33_ASAP7_75t_R g2700 ( 
.A(n_2409),
.Y(n_2700)
);

INVx2_ASAP7_75t_SL g2701 ( 
.A(n_2040),
.Y(n_2701)
);

INVx5_ASAP7_75t_L g2702 ( 
.A(n_2110),
.Y(n_2702)
);

INVx3_ASAP7_75t_SL g2703 ( 
.A(n_2115),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2398),
.Y(n_2704)
);

CKINVDCx16_ASAP7_75t_R g2705 ( 
.A(n_2185),
.Y(n_2705)
);

INVx2_ASAP7_75t_SL g2706 ( 
.A(n_2042),
.Y(n_2706)
);

NAND2x1p5_ASAP7_75t_L g2707 ( 
.A(n_2194),
.B(n_1788),
.Y(n_2707)
);

BUFx12f_ASAP7_75t_L g2708 ( 
.A(n_2157),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2194),
.Y(n_2709)
);

BUFx10_ASAP7_75t_L g2710 ( 
.A(n_2291),
.Y(n_2710)
);

INVxp67_ASAP7_75t_SL g2711 ( 
.A(n_2175),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2300),
.Y(n_2712)
);

BUFx3_ASAP7_75t_L g2713 ( 
.A(n_2420),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2300),
.Y(n_2714)
);

BUFx12f_ASAP7_75t_L g2715 ( 
.A(n_2159),
.Y(n_2715)
);

BUFx12f_ASAP7_75t_L g2716 ( 
.A(n_2062),
.Y(n_2716)
);

CKINVDCx11_ASAP7_75t_R g2717 ( 
.A(n_2423),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2115),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2437),
.B(n_1943),
.Y(n_2719)
);

INVx6_ASAP7_75t_L g2720 ( 
.A(n_2243),
.Y(n_2720)
);

NAND2x1p5_ASAP7_75t_L g2721 ( 
.A(n_2194),
.B(n_1788),
.Y(n_2721)
);

BUFx12f_ASAP7_75t_L g2722 ( 
.A(n_2238),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2110),
.Y(n_2723)
);

INVx4_ASAP7_75t_L g2724 ( 
.A(n_2198),
.Y(n_2724)
);

BUFx12f_ASAP7_75t_L g2725 ( 
.A(n_2064),
.Y(n_2725)
);

INVx1_ASAP7_75t_SL g2726 ( 
.A(n_2198),
.Y(n_2726)
);

BUFx2_ASAP7_75t_R g2727 ( 
.A(n_2162),
.Y(n_2727)
);

INVx1_ASAP7_75t_SL g2728 ( 
.A(n_2198),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2420),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2133),
.Y(n_2730)
);

BUFx4_ASAP7_75t_SL g2731 ( 
.A(n_2342),
.Y(n_2731)
);

BUFx6f_ASAP7_75t_L g2732 ( 
.A(n_2128),
.Y(n_2732)
);

INVx3_ASAP7_75t_SL g2733 ( 
.A(n_2119),
.Y(n_2733)
);

BUFx4_ASAP7_75t_SL g2734 ( 
.A(n_2342),
.Y(n_2734)
);

INVx3_ASAP7_75t_L g2735 ( 
.A(n_2204),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2457),
.Y(n_2736)
);

OR2x6_ASAP7_75t_L g2737 ( 
.A(n_2204),
.B(n_2207),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2204),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2133),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2207),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2307),
.B(n_2308),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2059),
.B(n_1968),
.Y(n_2742)
);

BUFx2_ASAP7_75t_SL g2743 ( 
.A(n_2119),
.Y(n_2743)
);

INVx1_ASAP7_75t_SL g2744 ( 
.A(n_2207),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2221),
.B(n_2250),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2398),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2256),
.B(n_1786),
.Y(n_2747)
);

BUFx3_ASAP7_75t_L g2748 ( 
.A(n_2144),
.Y(n_2748)
);

INVx5_ASAP7_75t_L g2749 ( 
.A(n_2128),
.Y(n_2749)
);

BUFx8_ASAP7_75t_L g2750 ( 
.A(n_2269),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2371),
.B(n_2355),
.Y(n_2751)
);

INVx1_ASAP7_75t_SL g2752 ( 
.A(n_2225),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2237),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2206),
.Y(n_2754)
);

BUFx2_ASAP7_75t_SL g2755 ( 
.A(n_2053),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2449),
.Y(n_2756)
);

INVxp67_ASAP7_75t_SL g2757 ( 
.A(n_2188),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_2144),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2125),
.Y(n_2759)
);

CKINVDCx20_ASAP7_75t_R g2760 ( 
.A(n_2370),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2351),
.B(n_1701),
.Y(n_2761)
);

BUFx12f_ASAP7_75t_L g2762 ( 
.A(n_2151),
.Y(n_2762)
);

NAND2x1p5_ASAP7_75t_L g2763 ( 
.A(n_2225),
.B(n_1799),
.Y(n_2763)
);

BUFx3_ASAP7_75t_L g2764 ( 
.A(n_2449),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2188),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2054),
.B(n_1706),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2089),
.Y(n_2767)
);

INVxp67_ASAP7_75t_SL g2768 ( 
.A(n_2192),
.Y(n_2768)
);

BUFx2_ASAP7_75t_SL g2769 ( 
.A(n_2053),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2457),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2050),
.B(n_2099),
.Y(n_2771)
);

BUFx2_ASAP7_75t_L g2772 ( 
.A(n_2463),
.Y(n_2772)
);

NAND2x1p5_ASAP7_75t_L g2773 ( 
.A(n_2225),
.B(n_1799),
.Y(n_2773)
);

BUFx12f_ASAP7_75t_L g2774 ( 
.A(n_2370),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2173),
.Y(n_2775)
);

NAND2x1p5_ASAP7_75t_L g2776 ( 
.A(n_2226),
.B(n_1695),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2177),
.Y(n_2777)
);

BUFx2_ASAP7_75t_L g2778 ( 
.A(n_2463),
.Y(n_2778)
);

CKINVDCx11_ASAP7_75t_R g2779 ( 
.A(n_2432),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2027),
.B(n_2308),
.Y(n_2780)
);

INVx2_ASAP7_75t_SL g2781 ( 
.A(n_2397),
.Y(n_2781)
);

NAND2x1p5_ASAP7_75t_L g2782 ( 
.A(n_2226),
.B(n_1695),
.Y(n_2782)
);

NAND2x1p5_ASAP7_75t_L g2783 ( 
.A(n_2226),
.B(n_2008),
.Y(n_2783)
);

INVx6_ASAP7_75t_L g2784 ( 
.A(n_2276),
.Y(n_2784)
);

INVx4_ASAP7_75t_L g2785 ( 
.A(n_2227),
.Y(n_2785)
);

BUFx4f_ASAP7_75t_SL g2786 ( 
.A(n_2382),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_2432),
.Y(n_2787)
);

BUFx3_ASAP7_75t_L g2788 ( 
.A(n_2051),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2199),
.A2(n_2004),
.B1(n_2005),
.B2(n_1845),
.Y(n_2789)
);

NAND2x1p5_ASAP7_75t_L g2790 ( 
.A(n_2227),
.B(n_2230),
.Y(n_2790)
);

BUFx4_ASAP7_75t_SL g2791 ( 
.A(n_2429),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2380),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2054),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2061),
.Y(n_2794)
);

INVxp67_ASAP7_75t_SL g2795 ( 
.A(n_2192),
.Y(n_2795)
);

HB1xp67_ASAP7_75t_L g2796 ( 
.A(n_2200),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2128),
.Y(n_2797)
);

INVx3_ASAP7_75t_L g2798 ( 
.A(n_2227),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2230),
.Y(n_2799)
);

INVxp67_ASAP7_75t_SL g2800 ( 
.A(n_2200),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2397),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2055),
.Y(n_2802)
);

INVx4_ASAP7_75t_L g2803 ( 
.A(n_2230),
.Y(n_2803)
);

OAI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_2104),
.A2(n_2120),
.B1(n_2154),
.B2(n_2203),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2326),
.Y(n_2805)
);

BUFx24_ASAP7_75t_L g2806 ( 
.A(n_2203),
.Y(n_2806)
);

BUFx5_ASAP7_75t_L g2807 ( 
.A(n_2086),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2190),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2068),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2355),
.B(n_1997),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_SL g2811 ( 
.A(n_2448),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2055),
.Y(n_2812)
);

BUFx3_ASAP7_75t_L g2813 ( 
.A(n_2245),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2088),
.Y(n_2814)
);

INVx4_ASAP7_75t_L g2815 ( 
.A(n_2235),
.Y(n_2815)
);

BUFx6f_ASAP7_75t_L g2816 ( 
.A(n_2240),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2276),
.Y(n_2817)
);

INVx1_ASAP7_75t_SL g2818 ( 
.A(n_2438),
.Y(n_2818)
);

BUFx12f_ASAP7_75t_L g2819 ( 
.A(n_2252),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2065),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2156),
.B(n_297),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2240),
.Y(n_2822)
);

AOI22xp33_ASAP7_75t_L g2823 ( 
.A1(n_2549),
.A2(n_2205),
.B1(n_2295),
.B2(n_2255),
.Y(n_2823)
);

INVx8_ASAP7_75t_L g2824 ( 
.A(n_2469),
.Y(n_2824)
);

BUFx10_ASAP7_75t_L g2825 ( 
.A(n_2473),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2468),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2470),
.Y(n_2827)
);

OAI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2583),
.A2(n_2304),
.B1(n_2169),
.B2(n_2265),
.Y(n_2828)
);

BUFx2_ASAP7_75t_L g2829 ( 
.A(n_2583),
.Y(n_2829)
);

CKINVDCx20_ASAP7_75t_R g2830 ( 
.A(n_2578),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2521),
.B(n_2075),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2479),
.Y(n_2832)
);

CKINVDCx20_ASAP7_75t_R g2833 ( 
.A(n_2578),
.Y(n_2833)
);

AOI22xp33_ASAP7_75t_SL g2834 ( 
.A1(n_2562),
.A2(n_2384),
.B1(n_2105),
.B2(n_2327),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2731),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2482),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2549),
.A2(n_2511),
.B1(n_2811),
.B2(n_2536),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2490),
.Y(n_2838)
);

AOI22xp33_ASAP7_75t_SL g2839 ( 
.A1(n_2562),
.A2(n_2105),
.B1(n_2405),
.B2(n_2352),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2579),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2497),
.Y(n_2841)
);

BUFx8_ASAP7_75t_SL g2842 ( 
.A(n_2504),
.Y(n_2842)
);

BUFx12f_ASAP7_75t_L g2843 ( 
.A(n_2473),
.Y(n_2843)
);

NAND2x1p5_ASAP7_75t_L g2844 ( 
.A(n_2472),
.B(n_2235),
.Y(n_2844)
);

INVx1_ASAP7_75t_SL g2845 ( 
.A(n_2806),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_SL g2846 ( 
.A1(n_2760),
.A2(n_2442),
.B1(n_2428),
.B2(n_2448),
.Y(n_2846)
);

CKINVDCx11_ASAP7_75t_R g2847 ( 
.A(n_2557),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2494),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2811),
.A2(n_2305),
.B1(n_2248),
.B2(n_2441),
.Y(n_2849)
);

BUFx2_ASAP7_75t_L g2850 ( 
.A(n_2505),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_2469),
.Y(n_2851)
);

CKINVDCx11_ASAP7_75t_R g2852 ( 
.A(n_2717),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2498),
.Y(n_2853)
);

AOI22xp33_ASAP7_75t_L g2854 ( 
.A1(n_2684),
.A2(n_2305),
.B1(n_2217),
.B2(n_2196),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2512),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2703),
.A2(n_2209),
.B1(n_2321),
.B2(n_2428),
.Y(n_2856)
);

OAI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2703),
.A2(n_2442),
.B1(n_2354),
.B2(n_2328),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2516),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2771),
.B(n_2745),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2570),
.Y(n_2860)
);

AOI22xp33_ASAP7_75t_SL g2861 ( 
.A1(n_2631),
.A2(n_2366),
.B1(n_2460),
.B2(n_2455),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2526),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2684),
.A2(n_2160),
.B1(n_2092),
.B2(n_2271),
.Y(n_2863)
);

AOI22xp33_ASAP7_75t_L g2864 ( 
.A1(n_2774),
.A2(n_2400),
.B1(n_2358),
.B2(n_2320),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_2545),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_L g2866 ( 
.A1(n_2529),
.A2(n_2400),
.B1(n_2184),
.B2(n_2285),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2529),
.A2(n_2326),
.B1(n_2451),
.B2(n_2306),
.Y(n_2867)
);

OAI21xp5_ASAP7_75t_SL g2868 ( 
.A1(n_2555),
.A2(n_2211),
.B(n_2195),
.Y(n_2868)
);

INVx8_ASAP7_75t_L g2869 ( 
.A(n_2469),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2493),
.Y(n_2870)
);

AOI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2529),
.A2(n_2451),
.B1(n_2253),
.B2(n_2459),
.Y(n_2871)
);

AOI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_2593),
.A2(n_2459),
.B1(n_2374),
.B2(n_2402),
.Y(n_2872)
);

OAI22xp33_ASAP7_75t_L g2873 ( 
.A1(n_2705),
.A2(n_2465),
.B1(n_2067),
.B2(n_2294),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2535),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2582),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2553),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2554),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_2527),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2563),
.Y(n_2879)
);

INVx6_ASAP7_75t_L g2880 ( 
.A(n_2514),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2619),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2565),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2567),
.Y(n_2883)
);

CKINVDCx11_ASAP7_75t_R g2884 ( 
.A(n_2717),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2647),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2666),
.Y(n_2886)
);

CKINVDCx20_ASAP7_75t_R g2887 ( 
.A(n_2467),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2741),
.B(n_2413),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2672),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2678),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2725),
.A2(n_2399),
.B1(n_2425),
.B2(n_2417),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2793),
.Y(n_2892)
);

INVx8_ASAP7_75t_L g2893 ( 
.A(n_2514),
.Y(n_2893)
);

BUFx5_ASAP7_75t_L g2894 ( 
.A(n_2656),
.Y(n_2894)
);

OAI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2664),
.A2(n_2419),
.B1(n_2081),
.B2(n_2082),
.Y(n_2895)
);

AOI22xp33_ASAP7_75t_L g2896 ( 
.A1(n_2779),
.A2(n_2452),
.B1(n_2302),
.B2(n_2216),
.Y(n_2896)
);

AOI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_2779),
.A2(n_2197),
.B1(n_2378),
.B2(n_2445),
.Y(n_2897)
);

BUFx12f_ASAP7_75t_L g2898 ( 
.A(n_2481),
.Y(n_2898)
);

INVx3_ASAP7_75t_L g2899 ( 
.A(n_2579),
.Y(n_2899)
);

BUFx10_ASAP7_75t_L g2900 ( 
.A(n_2630),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2688),
.Y(n_2901)
);

INVx1_ASAP7_75t_SL g2902 ( 
.A(n_2806),
.Y(n_2902)
);

INVx2_ASAP7_75t_SL g2903 ( 
.A(n_2514),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2667),
.A2(n_2410),
.B1(n_2414),
.B2(n_2411),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2667),
.A2(n_2414),
.B1(n_2224),
.B2(n_2078),
.Y(n_2905)
);

CKINVDCx11_ASAP7_75t_R g2906 ( 
.A(n_2495),
.Y(n_2906)
);

BUFx2_ASAP7_75t_SL g2907 ( 
.A(n_2492),
.Y(n_2907)
);

AOI22xp33_ASAP7_75t_L g2908 ( 
.A1(n_2667),
.A2(n_2084),
.B1(n_2179),
.B2(n_2458),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_SL g2909 ( 
.A1(n_2631),
.A2(n_2369),
.B1(n_2053),
.B2(n_2419),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_SL g2910 ( 
.A1(n_2631),
.A2(n_2369),
.B1(n_2053),
.B2(n_2377),
.Y(n_2910)
);

BUFx12f_ASAP7_75t_L g2911 ( 
.A(n_2698),
.Y(n_2911)
);

BUFx3_ASAP7_75t_L g2912 ( 
.A(n_2478),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_SL g2913 ( 
.A1(n_2539),
.A2(n_2406),
.B1(n_2431),
.B2(n_2329),
.Y(n_2913)
);

INVx11_ASAP7_75t_L g2914 ( 
.A(n_2722),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2736),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2770),
.Y(n_2916)
);

AOI22xp33_ASAP7_75t_L g2917 ( 
.A1(n_2694),
.A2(n_2401),
.B1(n_2228),
.B2(n_2186),
.Y(n_2917)
);

INVx4_ASAP7_75t_L g2918 ( 
.A(n_2486),
.Y(n_2918)
);

HB1xp67_ASAP7_75t_L g2919 ( 
.A(n_2634),
.Y(n_2919)
);

BUFx8_ASAP7_75t_L g2920 ( 
.A(n_2607),
.Y(n_2920)
);

INVx1_ASAP7_75t_SL g2921 ( 
.A(n_2733),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2475),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2802),
.Y(n_2923)
);

AOI22xp33_ASAP7_75t_L g2924 ( 
.A1(n_2669),
.A2(n_2364),
.B1(n_2404),
.B2(n_2372),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2480),
.Y(n_2925)
);

NAND2x1p5_ASAP7_75t_L g2926 ( 
.A(n_2492),
.B(n_2031),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_2731),
.Y(n_2927)
);

CKINVDCx20_ASAP7_75t_R g2928 ( 
.A(n_2485),
.Y(n_2928)
);

INVx4_ASAP7_75t_L g2929 ( 
.A(n_2486),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2812),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2820),
.Y(n_2931)
);

BUFx12f_ASAP7_75t_L g2932 ( 
.A(n_2700),
.Y(n_2932)
);

BUFx4_ASAP7_75t_SL g2933 ( 
.A(n_2515),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2753),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2488),
.Y(n_2935)
);

AOI22xp33_ASAP7_75t_L g2936 ( 
.A1(n_2669),
.A2(n_2416),
.B1(n_2340),
.B2(n_2314),
.Y(n_2936)
);

BUFx2_ASAP7_75t_L g2937 ( 
.A(n_2505),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2591),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2733),
.A2(n_2403),
.B1(n_2123),
.B2(n_2132),
.Y(n_2939)
);

OAI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2617),
.A2(n_2052),
.B1(n_2268),
.B2(n_2091),
.Y(n_2940)
);

INVx6_ASAP7_75t_L g2941 ( 
.A(n_2762),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2483),
.Y(n_2942)
);

INVx1_ASAP7_75t_SL g2943 ( 
.A(n_2743),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2489),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2809),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2683),
.A2(n_2281),
.B1(n_2232),
.B2(n_2391),
.Y(n_2946)
);

INVx3_ASAP7_75t_L g2947 ( 
.A(n_2474),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2814),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2533),
.Y(n_2949)
);

NAND2x1p5_ASAP7_75t_L g2950 ( 
.A(n_2676),
.B(n_2691),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2683),
.A2(n_2222),
.B1(n_2280),
.B2(n_2418),
.Y(n_2951)
);

AOI22xp33_ASAP7_75t_L g2952 ( 
.A1(n_2495),
.A2(n_2681),
.B1(n_2555),
.B2(n_2573),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2792),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2518),
.Y(n_2954)
);

INVx4_ASAP7_75t_SL g2955 ( 
.A(n_2630),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2681),
.A2(n_2083),
.B1(n_2069),
.B2(n_2032),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2533),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2533),
.Y(n_2958)
);

INVx6_ASAP7_75t_L g2959 ( 
.A(n_2598),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2595),
.Y(n_2960)
);

BUFx12f_ASAP7_75t_L g2961 ( 
.A(n_2660),
.Y(n_2961)
);

INVx6_ASAP7_75t_L g2962 ( 
.A(n_2604),
.Y(n_2962)
);

BUFx2_ASAP7_75t_L g2963 ( 
.A(n_2616),
.Y(n_2963)
);

OAI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2664),
.A2(n_2116),
.B1(n_2081),
.B2(n_2082),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2741),
.B(n_2596),
.Y(n_2965)
);

AOI22xp33_ASAP7_75t_L g2966 ( 
.A1(n_2558),
.A2(n_2288),
.B1(n_2283),
.B2(n_2440),
.Y(n_2966)
);

BUFx3_ASAP7_75t_L g2967 ( 
.A(n_2660),
.Y(n_2967)
);

OAI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2711),
.A2(n_2100),
.B1(n_2031),
.B2(n_2412),
.Y(n_2968)
);

BUFx12f_ASAP7_75t_L g2969 ( 
.A(n_2704),
.Y(n_2969)
);

BUFx4f_ASAP7_75t_L g2970 ( 
.A(n_2670),
.Y(n_2970)
);

INVx6_ASAP7_75t_L g2971 ( 
.A(n_2750),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2638),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2641),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2533),
.Y(n_2974)
);

OAI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2652),
.A2(n_2080),
.B1(n_2100),
.B2(n_2174),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2646),
.Y(n_2976)
);

BUFx3_ASAP7_75t_L g2977 ( 
.A(n_2633),
.Y(n_2977)
);

BUFx10_ASAP7_75t_L g2978 ( 
.A(n_2746),
.Y(n_2978)
);

OAI22xp5_ASAP7_75t_L g2979 ( 
.A1(n_2711),
.A2(n_2424),
.B1(n_2395),
.B2(n_2396),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2648),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2649),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2657),
.Y(n_2982)
);

BUFx6f_ASAP7_75t_L g2983 ( 
.A(n_2671),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_2547),
.Y(n_2984)
);

OAI21xp33_ASAP7_75t_L g2985 ( 
.A1(n_2661),
.A2(n_2180),
.B(n_2108),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2533),
.Y(n_2986)
);

OAI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2757),
.A2(n_2313),
.B1(n_2044),
.B2(n_2038),
.Y(n_2987)
);

BUFx2_ASAP7_75t_L g2988 ( 
.A(n_2559),
.Y(n_2988)
);

BUFx10_ASAP7_75t_L g2989 ( 
.A(n_2668),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2780),
.B(n_2118),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2658),
.Y(n_2991)
);

NAND2x1p5_ASAP7_75t_L g2992 ( 
.A(n_2676),
.B(n_2251),
.Y(n_2992)
);

CKINVDCx20_ASAP7_75t_R g2993 ( 
.A(n_2485),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2615),
.B(n_2093),
.Y(n_2994)
);

BUFx4f_ASAP7_75t_SL g2995 ( 
.A(n_2499),
.Y(n_2995)
);

AOI22xp33_ASAP7_75t_L g2996 ( 
.A1(n_2819),
.A2(n_2283),
.B1(n_2446),
.B2(n_2443),
.Y(n_2996)
);

BUFx4f_ASAP7_75t_SL g2997 ( 
.A(n_2592),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2757),
.A2(n_2430),
.B1(n_2095),
.B2(n_2189),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2734),
.Y(n_2999)
);

BUFx2_ASAP7_75t_L g3000 ( 
.A(n_2675),
.Y(n_3000)
);

CKINVDCx11_ASAP7_75t_R g3001 ( 
.A(n_2603),
.Y(n_3001)
);

HB1xp67_ASAP7_75t_L g3002 ( 
.A(n_2697),
.Y(n_3002)
);

INVx4_ASAP7_75t_L g3003 ( 
.A(n_2523),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2768),
.A2(n_2274),
.B1(n_2273),
.B2(n_2447),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2689),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2816),
.Y(n_3006)
);

INVx1_ASAP7_75t_SL g3007 ( 
.A(n_2542),
.Y(n_3007)
);

AOI22xp33_ASAP7_75t_L g3008 ( 
.A1(n_2661),
.A2(n_2139),
.B1(n_2450),
.B2(n_2309),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2659),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2610),
.B(n_2065),
.Y(n_3010)
);

OR2x2_ASAP7_75t_L g3011 ( 
.A(n_2754),
.B(n_2103),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2788),
.Y(n_3012)
);

INVx1_ASAP7_75t_SL g3013 ( 
.A(n_2542),
.Y(n_3013)
);

BUFx3_ASAP7_75t_L g3014 ( 
.A(n_2668),
.Y(n_3014)
);

INVx4_ASAP7_75t_SL g3015 ( 
.A(n_2532),
.Y(n_3015)
);

CKINVDCx11_ASAP7_75t_R g3016 ( 
.A(n_2574),
.Y(n_3016)
);

INVx3_ASAP7_75t_L g3017 ( 
.A(n_2474),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2605),
.A2(n_2231),
.B1(n_2260),
.B2(n_2223),
.Y(n_3018)
);

AOI22xp33_ASAP7_75t_SL g3019 ( 
.A1(n_2786),
.A2(n_2461),
.B1(n_1973),
.B2(n_1766),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2550),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2663),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2708),
.A2(n_2270),
.B1(n_2393),
.B2(n_2407),
.Y(n_3022)
);

OAI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2768),
.A2(n_2066),
.B1(n_2063),
.B2(n_2142),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_2715),
.A2(n_2407),
.B1(n_2096),
.B2(n_2153),
.Y(n_3024)
);

INVxp67_ASAP7_75t_SL g3025 ( 
.A(n_2795),
.Y(n_3025)
);

AOI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2677),
.A2(n_2150),
.B1(n_2341),
.B2(n_2299),
.Y(n_3026)
);

INVx6_ASAP7_75t_L g3027 ( 
.A(n_2750),
.Y(n_3027)
);

BUFx3_ASAP7_75t_L g3028 ( 
.A(n_2720),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2685),
.Y(n_3029)
);

INVx6_ASAP7_75t_L g3030 ( 
.A(n_2720),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2696),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2523),
.B(n_2368),
.Y(n_3032)
);

BUFx8_ASAP7_75t_SL g3033 ( 
.A(n_2687),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2712),
.Y(n_3034)
);

OAI22xp33_ASAP7_75t_L g3035 ( 
.A1(n_2787),
.A2(n_2046),
.B1(n_2113),
.B2(n_2072),
.Y(n_3035)
);

BUFx10_ASAP7_75t_L g3036 ( 
.A(n_2734),
.Y(n_3036)
);

INVx6_ASAP7_75t_L g3037 ( 
.A(n_2655),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2714),
.Y(n_3038)
);

OAI21xp33_ASAP7_75t_L g3039 ( 
.A1(n_2636),
.A2(n_2180),
.B(n_2290),
.Y(n_3039)
);

AOI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_2636),
.A2(n_2682),
.B1(n_2747),
.B2(n_2756),
.Y(n_3040)
);

AOI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2795),
.A2(n_2057),
.B1(n_2390),
.B2(n_2388),
.Y(n_3041)
);

OAI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2800),
.A2(n_2094),
.B1(n_2234),
.B2(n_2134),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2600),
.B(n_2072),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2800),
.A2(n_2071),
.B1(n_2331),
.B2(n_2316),
.Y(n_3044)
);

BUFx2_ASAP7_75t_SL g3045 ( 
.A(n_2523),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2503),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2794),
.Y(n_3047)
);

INVx3_ASAP7_75t_L g3048 ( 
.A(n_2691),
.Y(n_3048)
);

NAND2x1p5_ASAP7_75t_L g3049 ( 
.A(n_2525),
.B(n_2251),
.Y(n_3049)
);

INVx6_ASAP7_75t_L g3050 ( 
.A(n_2655),
.Y(n_3050)
);

BUFx4_ASAP7_75t_R g3051 ( 
.A(n_2626),
.Y(n_3051)
);

INVx6_ASAP7_75t_L g3052 ( 
.A(n_2710),
.Y(n_3052)
);

INVx3_ASAP7_75t_L g3053 ( 
.A(n_2530),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2751),
.Y(n_3054)
);

OAI22xp33_ASAP7_75t_R g3055 ( 
.A1(n_2626),
.A2(n_300),
.B1(n_297),
.B2(n_299),
.Y(n_3055)
);

OAI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2525),
.A2(n_2124),
.B1(n_2246),
.B2(n_2113),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_2606),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_SL g3058 ( 
.A1(n_2576),
.A2(n_1744),
.B(n_1957),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_2716),
.A2(n_2453),
.B1(n_2246),
.B2(n_2261),
.Y(n_3059)
);

AOI22xp33_ASAP7_75t_L g3060 ( 
.A1(n_2772),
.A2(n_2261),
.B1(n_2266),
.B2(n_2124),
.Y(n_3060)
);

HB1xp67_ASAP7_75t_L g3061 ( 
.A(n_2791),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2751),
.Y(n_3062)
);

CKINVDCx5p33_ASAP7_75t_R g3063 ( 
.A(n_2487),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2584),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2778),
.A2(n_2277),
.B1(n_2311),
.B2(n_2266),
.Y(n_3065)
);

BUFx2_ASAP7_75t_L g3066 ( 
.A(n_2599),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2590),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2611),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2628),
.A2(n_2311),
.B1(n_2324),
.B2(n_2277),
.Y(n_3069)
);

CKINVDCx20_ASAP7_75t_R g3070 ( 
.A(n_2532),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2807),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2612),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2807),
.Y(n_3073)
);

AOI22xp33_ASAP7_75t_L g3074 ( 
.A1(n_2628),
.A2(n_2324),
.B1(n_2345),
.B2(n_2344),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2767),
.A2(n_2353),
.B1(n_2346),
.B2(n_2178),
.Y(n_3075)
);

BUFx10_ASAP7_75t_L g3076 ( 
.A(n_2701),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_2775),
.A2(n_2158),
.B1(n_1845),
.B2(n_2362),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_SL g3078 ( 
.A1(n_2786),
.A2(n_1942),
.B1(n_2381),
.B2(n_2367),
.Y(n_3078)
);

INVx6_ASAP7_75t_L g3079 ( 
.A(n_2710),
.Y(n_3079)
);

INVx4_ASAP7_75t_L g3080 ( 
.A(n_2525),
.Y(n_3080)
);

INVx6_ASAP7_75t_L g3081 ( 
.A(n_2530),
.Y(n_3081)
);

INVx2_ASAP7_75t_SL g3082 ( 
.A(n_2791),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_SL g3083 ( 
.A1(n_2528),
.A2(n_2381),
.B1(n_2367),
.B2(n_1999),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_SL g3084 ( 
.A1(n_2528),
.A2(n_1784),
.B1(n_2436),
.B2(n_2239),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2807),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_SL g3086 ( 
.A1(n_2528),
.A2(n_2436),
.B1(n_2239),
.B2(n_2338),
.Y(n_3086)
);

HB1xp67_ASAP7_75t_L g3087 ( 
.A(n_2801),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2541),
.A2(n_2122),
.B1(n_2098),
.B2(n_2241),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2841),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_3055),
.A2(n_2815),
.B1(n_2789),
.B2(n_2500),
.Y(n_3090)
);

INVx3_ASAP7_75t_L g3091 ( 
.A(n_3003),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2859),
.B(n_2821),
.Y(n_3092)
);

AOI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_2939),
.A2(n_2994),
.B1(n_2845),
.B2(n_2902),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2878),
.B(n_2615),
.Y(n_3094)
);

INVx4_ASAP7_75t_SL g3095 ( 
.A(n_3081),
.Y(n_3095)
);

INVx2_ASAP7_75t_SL g3096 ( 
.A(n_2914),
.Y(n_3096)
);

CKINVDCx5p33_ASAP7_75t_R g3097 ( 
.A(n_3051),
.Y(n_3097)
);

OAI21xp5_ASAP7_75t_SL g3098 ( 
.A1(n_2845),
.A2(n_2585),
.B(n_2550),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2826),
.Y(n_3099)
);

AOI22xp33_ASAP7_75t_L g3100 ( 
.A1(n_2834),
.A2(n_2815),
.B1(n_2789),
.B2(n_2500),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_2902),
.A2(n_2500),
.B1(n_2476),
.B2(n_2810),
.Y(n_3101)
);

AOI222xp33_ASAP7_75t_L g3102 ( 
.A1(n_2823),
.A2(n_2556),
.B1(n_2586),
.B2(n_2551),
.C1(n_2524),
.C2(n_2777),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_2919),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2846),
.A2(n_2585),
.B1(n_2568),
.B2(n_2541),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_2852),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2938),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2860),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2934),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2827),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2875),
.Y(n_3110)
);

HB1xp67_ASAP7_75t_L g3111 ( 
.A(n_3002),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2832),
.Y(n_3112)
);

OAI22xp5_ASAP7_75t_L g3113 ( 
.A1(n_2846),
.A2(n_2568),
.B1(n_2541),
.B2(n_2764),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2839),
.A2(n_2500),
.B1(n_2476),
.B2(n_2810),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_2884),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_L g3116 ( 
.A1(n_2828),
.A2(n_2568),
.B1(n_2597),
.B2(n_2781),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_3000),
.Y(n_3117)
);

INVx5_ASAP7_75t_SL g3118 ( 
.A(n_2983),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_2990),
.B(n_2818),
.Y(n_3119)
);

AOI22xp33_ASAP7_75t_L g3120 ( 
.A1(n_2873),
.A2(n_2510),
.B1(n_2520),
.B2(n_2517),
.Y(n_3120)
);

AOI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_3004),
.A2(n_2692),
.B1(n_2713),
.B2(n_2693),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_3074),
.A2(n_2729),
.B1(n_2650),
.B2(n_2759),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_3054),
.B(n_2818),
.Y(n_3123)
);

BUFx6f_ASAP7_75t_L g3124 ( 
.A(n_2824),
.Y(n_3124)
);

OAI22xp5_ASAP7_75t_L g3125 ( 
.A1(n_2861),
.A2(n_2796),
.B1(n_2765),
.B2(n_2804),
.Y(n_3125)
);

BUFx2_ASAP7_75t_L g3126 ( 
.A(n_2983),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2836),
.Y(n_3127)
);

OAI221xp5_ASAP7_75t_L g3128 ( 
.A1(n_3018),
.A2(n_2863),
.B1(n_2966),
.B2(n_2924),
.C(n_2946),
.Y(n_3128)
);

INVx4_ASAP7_75t_SL g3129 ( 
.A(n_3081),
.Y(n_3129)
);

OAI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_2868),
.A2(n_2796),
.B1(n_2765),
.B2(n_2727),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_SL g3131 ( 
.A1(n_2857),
.A2(n_2544),
.B1(n_2491),
.B2(n_2484),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_SL g3132 ( 
.A1(n_2943),
.A2(n_2544),
.B1(n_2491),
.B2(n_2484),
.Y(n_3132)
);

BUFx3_ASAP7_75t_L g3133 ( 
.A(n_2824),
.Y(n_3133)
);

AOI22xp33_ASAP7_75t_L g3134 ( 
.A1(n_3019),
.A2(n_2650),
.B1(n_2594),
.B2(n_2571),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_3062),
.A2(n_2556),
.B1(n_2804),
.B2(n_2586),
.Y(n_3135)
);

NOR2x1_ASAP7_75t_L g3136 ( 
.A(n_2868),
.B(n_2538),
.Y(n_3136)
);

AOI22xp33_ASAP7_75t_L g3137 ( 
.A1(n_2979),
.A2(n_2706),
.B1(n_2690),
.B2(n_2639),
.Y(n_3137)
);

HB1xp67_ASAP7_75t_L g3138 ( 
.A(n_3011),
.Y(n_3138)
);

CKINVDCx20_ASAP7_75t_R g3139 ( 
.A(n_2830),
.Y(n_3139)
);

INVx4_ASAP7_75t_L g3140 ( 
.A(n_2824),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2881),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2979),
.A2(n_2718),
.B1(n_2651),
.B2(n_2614),
.Y(n_3142)
);

OAI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_2844),
.A2(n_2501),
.B1(n_2466),
.B2(n_2508),
.Y(n_3143)
);

OAI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_2987),
.A2(n_2509),
.B1(n_2508),
.B2(n_2727),
.Y(n_3144)
);

OAI22xp5_ASAP7_75t_L g3145 ( 
.A1(n_2987),
.A2(n_2509),
.B1(n_2620),
.B2(n_2618),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2998),
.A2(n_2627),
.B1(n_2637),
.B2(n_2622),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_3069),
.A2(n_2651),
.B1(n_2496),
.B2(n_2742),
.Y(n_3147)
);

AOI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_3035),
.A2(n_2742),
.B1(n_2719),
.B2(n_2608),
.Y(n_3148)
);

OAI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_2998),
.A2(n_2501),
.B1(n_2466),
.B2(n_2544),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2885),
.Y(n_3150)
);

BUFx3_ASAP7_75t_L g3151 ( 
.A(n_2869),
.Y(n_3151)
);

OAI21xp33_ASAP7_75t_L g3152 ( 
.A1(n_3039),
.A2(n_2215),
.B(n_2181),
.Y(n_3152)
);

HB1xp67_ASAP7_75t_L g3153 ( 
.A(n_2943),
.Y(n_3153)
);

OAI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_2909),
.A2(n_2719),
.B1(n_2608),
.B2(n_2496),
.Y(n_3154)
);

BUFx2_ASAP7_75t_L g3155 ( 
.A(n_2983),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_2984),
.Y(n_3156)
);

BUFx4f_ASAP7_75t_SL g3157 ( 
.A(n_2833),
.Y(n_3157)
);

BUFx12f_ASAP7_75t_L g3158 ( 
.A(n_3036),
.Y(n_3158)
);

INVx4_ASAP7_75t_L g3159 ( 
.A(n_2869),
.Y(n_3159)
);

INVx4_ASAP7_75t_L g3160 ( 
.A(n_2869),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_SL g3161 ( 
.A1(n_2913),
.A2(n_2644),
.B(n_2566),
.Y(n_3161)
);

AOI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_2956),
.A2(n_2577),
.B1(n_2623),
.B2(n_2581),
.Y(n_3162)
);

AND2x4_ASAP7_75t_SL g3163 ( 
.A(n_3036),
.B(n_2538),
.Y(n_3163)
);

AOI222xp33_ASAP7_75t_L g3164 ( 
.A1(n_3015),
.A2(n_2551),
.B1(n_2524),
.B2(n_2587),
.C1(n_2519),
.C2(n_2761),
.Y(n_3164)
);

AOI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_2896),
.A2(n_2577),
.B1(n_2629),
.B2(n_2761),
.Y(n_3165)
);

AOI22xp33_ASAP7_75t_SL g3166 ( 
.A1(n_2856),
.A2(n_2537),
.B1(n_2502),
.B2(n_2755),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2895),
.A2(n_2968),
.B(n_3058),
.Y(n_3167)
);

INVx4_ASAP7_75t_L g3168 ( 
.A(n_2893),
.Y(n_3168)
);

CKINVDCx5p33_ASAP7_75t_R g3169 ( 
.A(n_3001),
.Y(n_3169)
);

OAI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_2905),
.A2(n_2560),
.B1(n_2566),
.B2(n_2644),
.Y(n_3170)
);

INVx2_ASAP7_75t_SL g3171 ( 
.A(n_2893),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_3040),
.A2(n_2625),
.B1(n_2654),
.B2(n_2580),
.Y(n_3172)
);

BUFx4f_ASAP7_75t_L g3173 ( 
.A(n_2893),
.Y(n_3173)
);

CKINVDCx16_ASAP7_75t_R g3174 ( 
.A(n_2928),
.Y(n_3174)
);

AOI22xp33_ASAP7_75t_L g3175 ( 
.A1(n_2831),
.A2(n_2625),
.B1(n_2654),
.B2(n_2580),
.Y(n_3175)
);

AOI22xp33_ASAP7_75t_SL g3176 ( 
.A1(n_2840),
.A2(n_2899),
.B1(n_2907),
.B2(n_3045),
.Y(n_3176)
);

OAI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_3025),
.A2(n_2560),
.B1(n_2766),
.B2(n_2548),
.Y(n_3177)
);

HB1xp67_ASAP7_75t_L g3178 ( 
.A(n_2988),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2886),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2838),
.Y(n_3180)
);

AOI22xp33_ASAP7_75t_L g3181 ( 
.A1(n_2975),
.A2(n_2665),
.B1(n_2624),
.B2(n_2531),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2848),
.Y(n_3182)
);

NAND3xp33_ASAP7_75t_L g3183 ( 
.A(n_2985),
.B(n_3039),
.C(n_2891),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_3012),
.B(n_2601),
.Y(n_3184)
);

OAI21xp5_ASAP7_75t_SL g3185 ( 
.A1(n_3061),
.A2(n_2624),
.B(n_2548),
.Y(n_3185)
);

AOI22xp33_ASAP7_75t_SL g3186 ( 
.A1(n_2840),
.A2(n_2899),
.B1(n_2895),
.B2(n_2971),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_3023),
.A2(n_2665),
.B1(n_2531),
.B2(n_2609),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2853),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2855),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_L g3190 ( 
.A1(n_2940),
.A2(n_2609),
.B1(n_2805),
.B2(n_2724),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2953),
.B(n_2960),
.Y(n_3191)
);

OAI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_3042),
.A2(n_2766),
.B1(n_2569),
.B2(n_2572),
.Y(n_3192)
);

AOI22xp33_ASAP7_75t_SL g3193 ( 
.A1(n_2971),
.A2(n_2769),
.B1(n_2807),
.B2(n_2540),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_2985),
.A2(n_2724),
.B1(n_2785),
.B2(n_2709),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_3026),
.A2(n_2785),
.B1(n_2803),
.B2(n_2709),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_2871),
.A2(n_2543),
.B1(n_2807),
.B2(n_2564),
.Y(n_3196)
);

CKINVDCx20_ASAP7_75t_R g3197 ( 
.A(n_2847),
.Y(n_3197)
);

OR2x2_ASAP7_75t_SL g3198 ( 
.A(n_3027),
.B(n_2784),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_3047),
.B(n_2808),
.Y(n_3199)
);

OAI21xp5_ASAP7_75t_SL g3200 ( 
.A1(n_2910),
.A2(n_2572),
.B(n_2569),
.Y(n_3200)
);

CKINVDCx11_ASAP7_75t_R g3201 ( 
.A(n_2825),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3010),
.B(n_2817),
.Y(n_3202)
);

INVx3_ASAP7_75t_L g3203 ( 
.A(n_3003),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2889),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_3005),
.B(n_2813),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_2872),
.A2(n_2534),
.B1(n_2784),
.B2(n_2737),
.Y(n_3206)
);

OAI222xp33_ASAP7_75t_L g3207 ( 
.A1(n_3056),
.A2(n_2540),
.B1(n_2737),
.B2(n_2645),
.C1(n_2726),
.C2(n_2602),
.Y(n_3207)
);

OAI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_3042),
.A2(n_2783),
.B1(n_2707),
.B2(n_2763),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_2951),
.A2(n_2803),
.B1(n_2642),
.B2(n_2645),
.Y(n_3209)
);

INVx3_ASAP7_75t_L g3210 ( 
.A(n_3080),
.Y(n_3210)
);

BUFx6f_ASAP7_75t_L g3211 ( 
.A(n_3005),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_2835),
.Y(n_3212)
);

CKINVDCx5p33_ASAP7_75t_R g3213 ( 
.A(n_2927),
.Y(n_3213)
);

AOI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_3008),
.A2(n_2888),
.B1(n_3024),
.B2(n_3022),
.Y(n_3214)
);

HB1xp67_ASAP7_75t_L g3215 ( 
.A(n_2890),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2858),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_2897),
.A2(n_2662),
.B1(n_2679),
.B2(n_2653),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2862),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3005),
.B(n_299),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2901),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_2965),
.B(n_300),
.Y(n_3221)
);

BUFx4f_ASAP7_75t_SL g3222 ( 
.A(n_2843),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_2999),
.Y(n_3223)
);

AOI22xp33_ASAP7_75t_L g3224 ( 
.A1(n_2908),
.A2(n_2662),
.B1(n_2679),
.B2(n_2653),
.Y(n_3224)
);

OR2x2_ASAP7_75t_L g3225 ( 
.A(n_2915),
.B(n_2916),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2874),
.B(n_2602),
.Y(n_3226)
);

OAI21xp5_ASAP7_75t_SL g3227 ( 
.A1(n_3082),
.A2(n_2790),
.B(n_2673),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2922),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2876),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3078),
.A2(n_2783),
.B1(n_2707),
.B2(n_2763),
.Y(n_3230)
);

OAI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_3044),
.A2(n_2721),
.B1(n_2773),
.B2(n_2686),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_SL g3232 ( 
.A1(n_3027),
.A2(n_2739),
.B1(n_2748),
.B2(n_2730),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2877),
.B(n_2632),
.Y(n_3233)
);

AOI22xp33_ASAP7_75t_L g3234 ( 
.A1(n_2936),
.A2(n_2738),
.B1(n_2798),
.B2(n_2735),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2879),
.B(n_2632),
.Y(n_3235)
);

OAI222xp33_ASAP7_75t_L g3236 ( 
.A1(n_3056),
.A2(n_2737),
.B1(n_2680),
.B2(n_2728),
.C1(n_2673),
.C2(n_2744),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_3044),
.A2(n_2773),
.B1(n_2721),
.B2(n_2686),
.Y(n_3237)
);

OAI22xp5_ASAP7_75t_L g3238 ( 
.A1(n_3041),
.A2(n_3083),
.B1(n_3060),
.B2(n_3065),
.Y(n_3238)
);

AOI22xp33_ASAP7_75t_L g3239 ( 
.A1(n_2996),
.A2(n_2738),
.B1(n_2798),
.B2(n_2735),
.Y(n_3239)
);

AOI22xp33_ASAP7_75t_L g3240 ( 
.A1(n_3075),
.A2(n_2799),
.B1(n_2575),
.B2(n_2758),
.Y(n_3240)
);

AOI22xp33_ASAP7_75t_L g3241 ( 
.A1(n_2854),
.A2(n_2799),
.B1(n_2575),
.B2(n_2426),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2925),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2882),
.B(n_2680),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2883),
.Y(n_3244)
);

BUFx12f_ASAP7_75t_L g3245 ( 
.A(n_2906),
.Y(n_3245)
);

AO22x1_ASAP7_75t_L g3246 ( 
.A1(n_2920),
.A2(n_2640),
.B1(n_2702),
.B2(n_2588),
.Y(n_3246)
);

AOI22xp33_ASAP7_75t_L g3247 ( 
.A1(n_2849),
.A2(n_2338),
.B1(n_2728),
.B2(n_2726),
.Y(n_3247)
);

AOI22xp33_ASAP7_75t_L g3248 ( 
.A1(n_2866),
.A2(n_2744),
.B1(n_2752),
.B2(n_2740),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2944),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_SL g3250 ( 
.A1(n_2829),
.A2(n_2921),
.B1(n_3050),
.B2(n_3037),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_2921),
.B(n_2740),
.Y(n_3251)
);

BUFx3_ASAP7_75t_L g3252 ( 
.A(n_2941),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_2941),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3046),
.B(n_301),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_2837),
.A2(n_2752),
.B1(n_2434),
.B2(n_2239),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_2904),
.A2(n_2917),
.B1(n_3059),
.B2(n_2864),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2892),
.Y(n_3257)
);

AOI22xp33_ASAP7_75t_L g3258 ( 
.A1(n_3041),
.A2(n_2434),
.B1(n_2239),
.B2(n_2275),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_2867),
.A2(n_2275),
.B1(n_2439),
.B2(n_2436),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_SL g3260 ( 
.A1(n_3037),
.A2(n_2640),
.B1(n_2702),
.B2(n_2588),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_2952),
.A2(n_2790),
.B1(n_2408),
.B2(n_2640),
.Y(n_3261)
);

NOR2xp33_ASAP7_75t_L g3262 ( 
.A(n_2887),
.B(n_302),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2945),
.Y(n_3263)
);

CKINVDCx5p33_ASAP7_75t_R g3264 ( 
.A(n_2842),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2923),
.B(n_2247),
.Y(n_3265)
);

OAI21xp5_ASAP7_75t_SL g3266 ( 
.A1(n_2963),
.A2(n_2782),
.B(n_2776),
.Y(n_3266)
);

OAI21xp5_ASAP7_75t_SL g3267 ( 
.A1(n_2926),
.A2(n_2782),
.B(n_2776),
.Y(n_3267)
);

INVx2_ASAP7_75t_SL g3268 ( 
.A(n_2880),
.Y(n_3268)
);

OAI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_2970),
.A2(n_2408),
.B1(n_2702),
.B2(n_2588),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2930),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_3077),
.A2(n_2275),
.B1(n_2439),
.B2(n_2161),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_L g3272 ( 
.A1(n_2967),
.A2(n_2275),
.B1(n_2161),
.B2(n_2171),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_2880),
.A2(n_2267),
.B1(n_2254),
.B2(n_2171),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_SL g3274 ( 
.A1(n_3050),
.A2(n_2749),
.B1(n_2368),
.B2(n_2415),
.Y(n_3274)
);

AOI22xp33_ASAP7_75t_L g3275 ( 
.A1(n_3066),
.A2(n_2166),
.B1(n_2415),
.B2(n_2368),
.Y(n_3275)
);

AOI22xp33_ASAP7_75t_L g3276 ( 
.A1(n_3087),
.A2(n_2166),
.B1(n_2415),
.B2(n_2310),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2931),
.Y(n_3277)
);

OAI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3058),
.A2(n_2315),
.B1(n_2337),
.B2(n_2286),
.Y(n_3278)
);

OAI21xp5_ASAP7_75t_SL g3279 ( 
.A1(n_2950),
.A2(n_2073),
.B(n_2060),
.Y(n_3279)
);

INVx1_ASAP7_75t_SL g3280 ( 
.A(n_3007),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_2948),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_2865),
.B(n_302),
.Y(n_3282)
);

AOI22xp33_ASAP7_75t_L g3283 ( 
.A1(n_3102),
.A2(n_2973),
.B1(n_2976),
.B2(n_2972),
.Y(n_3283)
);

OAI221xp5_ASAP7_75t_L g3284 ( 
.A1(n_3128),
.A2(n_2970),
.B1(n_2850),
.B2(n_2937),
.C(n_3043),
.Y(n_3284)
);

OAI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3090),
.A2(n_3053),
.B1(n_3048),
.B2(n_3070),
.Y(n_3285)
);

OAI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_3137),
.A2(n_3053),
.B1(n_3048),
.B2(n_3017),
.Y(n_3286)
);

NAND3xp33_ASAP7_75t_L g3287 ( 
.A(n_3183),
.B(n_2981),
.C(n_2980),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_SL g3288 ( 
.A1(n_3130),
.A2(n_3144),
.B1(n_3125),
.B2(n_3149),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_3102),
.A2(n_2982),
.B1(n_3009),
.B2(n_2991),
.Y(n_3289)
);

AOI22xp33_ASAP7_75t_L g3290 ( 
.A1(n_3164),
.A2(n_3029),
.B1(n_3031),
.B2(n_3021),
.Y(n_3290)
);

AOI21xp33_ASAP7_75t_L g3291 ( 
.A1(n_3164),
.A2(n_3013),
.B(n_3007),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_3238),
.A2(n_3038),
.B1(n_3034),
.B2(n_3064),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_L g3293 ( 
.A1(n_3238),
.A2(n_3068),
.B1(n_3072),
.B2(n_3067),
.Y(n_3293)
);

HB1xp67_ASAP7_75t_L g3294 ( 
.A(n_3103),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3099),
.Y(n_3295)
);

OAI21xp5_ASAP7_75t_SL g3296 ( 
.A1(n_3161),
.A2(n_3185),
.B(n_3166),
.Y(n_3296)
);

AOI222xp33_ASAP7_75t_SL g3297 ( 
.A1(n_3125),
.A2(n_2933),
.B1(n_2955),
.B2(n_2920),
.C1(n_2997),
.C2(n_3015),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3092),
.A2(n_3052),
.B1(n_3079),
.B2(n_2968),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3138),
.B(n_3013),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3109),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3215),
.B(n_3020),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_3134),
.A2(n_3020),
.B1(n_2964),
.B2(n_3080),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_3154),
.A2(n_3028),
.B1(n_3014),
.B2(n_2894),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_SL g3304 ( 
.A1(n_3144),
.A2(n_3079),
.B1(n_3052),
.B2(n_3088),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3119),
.B(n_2942),
.Y(n_3305)
);

OAI21xp33_ASAP7_75t_L g3306 ( 
.A1(n_3167),
.A2(n_2215),
.B(n_2181),
.Y(n_3306)
);

AOI22xp33_ASAP7_75t_L g3307 ( 
.A1(n_3154),
.A2(n_2894),
.B1(n_3030),
.B2(n_3017),
.Y(n_3307)
);

INVx4_ASAP7_75t_L g3308 ( 
.A(n_3095),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3106),
.B(n_2894),
.Y(n_3309)
);

OAI21xp5_ASAP7_75t_SL g3310 ( 
.A1(n_3136),
.A2(n_2903),
.B(n_2851),
.Y(n_3310)
);

AOI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_3214),
.A2(n_2961),
.B1(n_2918),
.B2(n_2929),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3114),
.A2(n_2894),
.B1(n_3030),
.B2(n_2947),
.Y(n_3312)
);

AOI22xp33_ASAP7_75t_L g3313 ( 
.A1(n_3149),
.A2(n_2894),
.B1(n_2947),
.B2(n_2870),
.Y(n_3313)
);

AOI22xp33_ASAP7_75t_L g3314 ( 
.A1(n_3100),
.A2(n_2912),
.B1(n_2954),
.B2(n_2935),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_3101),
.A2(n_3088),
.B1(n_3084),
.B2(n_2957),
.Y(n_3315)
);

AOI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3148),
.A2(n_2929),
.B1(n_2918),
.B2(n_2959),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_3094),
.A2(n_2949),
.B1(n_2974),
.B2(n_2958),
.Y(n_3317)
);

AOI22xp33_ASAP7_75t_L g3318 ( 
.A1(n_3256),
.A2(n_2986),
.B1(n_3073),
.B2(n_3071),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_3142),
.A2(n_3085),
.B1(n_2977),
.B2(n_2898),
.Y(n_3319)
);

OAI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3093),
.A2(n_3086),
.B1(n_2993),
.B2(n_2992),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3147),
.A2(n_3016),
.B1(n_2900),
.B2(n_2989),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3131),
.A2(n_3049),
.B1(n_2959),
.B2(n_2962),
.Y(n_3322)
);

AOI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_3146),
.A2(n_2900),
.B1(n_2989),
.B2(n_2825),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3123),
.B(n_3076),
.Y(n_3324)
);

AOI222xp33_ASAP7_75t_L g3325 ( 
.A1(n_3173),
.A2(n_2955),
.B1(n_2995),
.B2(n_2962),
.C1(n_3063),
.C2(n_3057),
.Y(n_3325)
);

AOI22xp33_ASAP7_75t_SL g3326 ( 
.A1(n_3177),
.A2(n_3076),
.B1(n_3006),
.B2(n_2932),
.Y(n_3326)
);

AOI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_3146),
.A2(n_2210),
.B1(n_3032),
.B2(n_2359),
.Y(n_3327)
);

AOI22xp33_ASAP7_75t_L g3328 ( 
.A1(n_3165),
.A2(n_2359),
.B1(n_3006),
.B2(n_2258),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3117),
.B(n_3006),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3156),
.B(n_304),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3108),
.B(n_304),
.Y(n_3331)
);

OAI22xp5_ASAP7_75t_L g3332 ( 
.A1(n_3198),
.A2(n_2749),
.B1(n_2060),
.B2(n_2114),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3112),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_3177),
.A2(n_2258),
.B1(n_2264),
.B2(n_2240),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_SL g3335 ( 
.A1(n_3104),
.A2(n_3113),
.B1(n_3170),
.B2(n_3178),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_SL g3336 ( 
.A1(n_3104),
.A2(n_2978),
.B1(n_2911),
.B2(n_2969),
.Y(n_3336)
);

NAND3xp33_ASAP7_75t_L g3337 ( 
.A(n_3153),
.B(n_2749),
.C(n_1953),
.Y(n_3337)
);

OAI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_3140),
.A2(n_2822),
.B1(n_2816),
.B2(n_2477),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3186),
.A2(n_2264),
.B1(n_2258),
.B2(n_2373),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3225),
.Y(n_3340)
);

AOI211xp5_ASAP7_75t_L g3341 ( 
.A1(n_3098),
.A2(n_2422),
.B(n_2444),
.C(n_2433),
.Y(n_3341)
);

NAND3xp33_ASAP7_75t_L g3342 ( 
.A(n_3240),
.B(n_1953),
.C(n_2454),
.Y(n_3342)
);

AOI22xp33_ASAP7_75t_L g3343 ( 
.A1(n_3111),
.A2(n_2264),
.B1(n_2464),
.B2(n_2456),
.Y(n_3343)
);

AOI22xp33_ASAP7_75t_L g3344 ( 
.A1(n_3145),
.A2(n_2114),
.B1(n_2073),
.B2(n_2816),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_3145),
.A2(n_2822),
.B1(n_2477),
.B2(n_2506),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3184),
.B(n_305),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3135),
.A2(n_2822),
.B1(n_2477),
.B2(n_2506),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3127),
.Y(n_3348)
);

AOI22xp33_ASAP7_75t_L g3349 ( 
.A1(n_3241),
.A2(n_2506),
.B1(n_2507),
.B2(n_2471),
.Y(n_3349)
);

NAND3xp33_ASAP7_75t_L g3350 ( 
.A(n_3162),
.B(n_3250),
.C(n_3190),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3221),
.A2(n_2507),
.B1(n_2513),
.B2(n_2471),
.Y(n_3351)
);

NAND3xp33_ASAP7_75t_SL g3352 ( 
.A(n_3097),
.B(n_3033),
.C(n_2978),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3122),
.A2(n_2507),
.B1(n_2513),
.B2(n_2471),
.Y(n_3353)
);

AOI221xp5_ASAP7_75t_L g3354 ( 
.A1(n_3254),
.A2(n_1704),
.B1(n_1703),
.B2(n_308),
.C(n_309),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_SL g3355 ( 
.A1(n_3139),
.A2(n_2522),
.B1(n_2546),
.B2(n_2513),
.Y(n_3355)
);

AOI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3121),
.A2(n_1704),
.B1(n_1703),
.B2(n_2522),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3192),
.A2(n_2546),
.B1(n_2552),
.B2(n_2522),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_SL g3358 ( 
.A1(n_3192),
.A2(n_3159),
.B1(n_3160),
.B2(n_3140),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3180),
.B(n_305),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_3116),
.A2(n_2552),
.B1(n_2561),
.B2(n_2546),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_3120),
.A2(n_2561),
.B1(n_2589),
.B2(n_2552),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_3219),
.A2(n_2589),
.B1(n_2613),
.B2(n_2561),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3182),
.B(n_306),
.Y(n_3363)
);

OAI221xp5_ASAP7_75t_L g3364 ( 
.A1(n_3234),
.A2(n_2797),
.B1(n_2732),
.B2(n_2723),
.C(n_2699),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_3258),
.A2(n_2613),
.B1(n_2621),
.B2(n_2589),
.Y(n_3365)
);

OAI222xp33_ASAP7_75t_L g3366 ( 
.A1(n_3176),
.A2(n_3159),
.B1(n_3160),
.B2(n_3168),
.C1(n_3193),
.C2(n_3132),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_3282),
.A2(n_2621),
.B1(n_2635),
.B2(n_2613),
.Y(n_3367)
);

OAI222xp33_ASAP7_75t_L g3368 ( 
.A1(n_3168),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.C1(n_312),
.C2(n_313),
.Y(n_3368)
);

AOI22xp33_ASAP7_75t_L g3369 ( 
.A1(n_3202),
.A2(n_3231),
.B1(n_3237),
.B2(n_3217),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_3187),
.A2(n_2635),
.B1(n_2643),
.B2(n_2621),
.Y(n_3370)
);

OAI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_3181),
.A2(n_2643),
.B1(n_2674),
.B2(n_2635),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_3199),
.B(n_3188),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3189),
.B(n_312),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_SL g3374 ( 
.A1(n_3173),
.A2(n_2674),
.B1(n_2695),
.B2(n_2643),
.Y(n_3374)
);

AOI22xp5_ASAP7_75t_L g3375 ( 
.A1(n_3196),
.A2(n_3239),
.B1(n_3206),
.B2(n_3248),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3231),
.A2(n_3237),
.B1(n_3278),
.B2(n_3251),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_3158),
.A2(n_2695),
.B1(n_2699),
.B2(n_2674),
.Y(n_3377)
);

OAI21xp5_ASAP7_75t_SL g3378 ( 
.A1(n_3163),
.A2(n_2699),
.B(n_2695),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3262),
.A2(n_2732),
.B1(n_2797),
.B2(n_2723),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_3257),
.A2(n_2732),
.B1(n_2797),
.B2(n_2723),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_3091),
.Y(n_3381)
);

OAI221xp5_ASAP7_75t_SL g3382 ( 
.A1(n_3200),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.C(n_317),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3216),
.B(n_314),
.Y(n_3383)
);

OAI222xp33_ASAP7_75t_L g3384 ( 
.A1(n_3230),
.A2(n_3143),
.B1(n_3172),
.B2(n_3091),
.C1(n_3210),
.C2(n_3203),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3175),
.A2(n_318),
.B1(n_315),
.B2(n_316),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3218),
.B(n_318),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_3280),
.Y(n_3387)
);

AOI22xp33_ASAP7_75t_L g3388 ( 
.A1(n_3270),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3229),
.B(n_321),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_3244),
.B(n_322),
.Y(n_3390)
);

AOI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3224),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_3277),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_3278),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_3393)
);

OAI22xp5_ASAP7_75t_L g3394 ( 
.A1(n_3209),
.A2(n_328),
.B1(n_329),
.B2(n_334),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_SL g3395 ( 
.A1(n_3230),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3205),
.B(n_335),
.Y(n_3396)
);

OAI21xp33_ASAP7_75t_SL g3397 ( 
.A1(n_3203),
.A2(n_3210),
.B(n_3194),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3245),
.A2(n_3191),
.B1(n_3152),
.B2(n_3124),
.Y(n_3398)
);

AOI22xp33_ASAP7_75t_L g3399 ( 
.A1(n_3124),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_3124),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3247),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3126),
.B(n_340),
.Y(n_3402)
);

AOI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3226),
.A2(n_342),
.B1(n_343),
.B2(n_346),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3372),
.B(n_3280),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3340),
.B(n_3089),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3294),
.B(n_3107),
.Y(n_3406)
);

OAI221xp5_ASAP7_75t_SL g3407 ( 
.A1(n_3296),
.A2(n_3227),
.B1(n_3266),
.B2(n_3133),
.C(n_3151),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3283),
.B(n_3110),
.Y(n_3408)
);

NAND4xp25_ASAP7_75t_L g3409 ( 
.A(n_3288),
.B(n_3255),
.C(n_3195),
.D(n_3232),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_3352),
.B(n_3174),
.Y(n_3410)
);

OAI221xp5_ASAP7_75t_SL g3411 ( 
.A1(n_3292),
.A2(n_3171),
.B1(n_3267),
.B2(n_3252),
.C(n_3253),
.Y(n_3411)
);

NOR3xp33_ASAP7_75t_L g3412 ( 
.A(n_3382),
.B(n_3246),
.C(n_3201),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_SL g3413 ( 
.A1(n_3308),
.A2(n_3261),
.B(n_3269),
.Y(n_3413)
);

AOI221xp5_ASAP7_75t_L g3414 ( 
.A1(n_3292),
.A2(n_3233),
.B1(n_3243),
.B2(n_3235),
.C(n_3268),
.Y(n_3414)
);

AOI221xp5_ASAP7_75t_L g3415 ( 
.A1(n_3293),
.A2(n_3265),
.B1(n_3207),
.B2(n_3236),
.C(n_3169),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3283),
.B(n_3141),
.Y(n_3416)
);

INVxp67_ASAP7_75t_L g3417 ( 
.A(n_3387),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3305),
.B(n_3155),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3289),
.B(n_3150),
.Y(n_3419)
);

AND2x2_ASAP7_75t_L g3420 ( 
.A(n_3329),
.B(n_3179),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3289),
.B(n_3293),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3324),
.B(n_3204),
.Y(n_3422)
);

OR2x2_ASAP7_75t_L g3423 ( 
.A(n_3299),
.B(n_3220),
.Y(n_3423)
);

NAND3xp33_ASAP7_75t_L g3424 ( 
.A(n_3287),
.B(n_3208),
.C(n_3211),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3295),
.B(n_3228),
.Y(n_3425)
);

NAND3xp33_ASAP7_75t_L g3426 ( 
.A(n_3350),
.B(n_3208),
.C(n_3211),
.Y(n_3426)
);

NAND3xp33_ASAP7_75t_L g3427 ( 
.A(n_3304),
.B(n_3284),
.C(n_3398),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3300),
.B(n_3242),
.Y(n_3428)
);

OAI221xp5_ASAP7_75t_SL g3429 ( 
.A1(n_3290),
.A2(n_3298),
.B1(n_3323),
.B2(n_3358),
.C(n_3321),
.Y(n_3429)
);

OAI221xp5_ASAP7_75t_SL g3430 ( 
.A1(n_3290),
.A2(n_3096),
.B1(n_3279),
.B2(n_3271),
.C(n_3259),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3333),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3348),
.B(n_3249),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3301),
.B(n_3263),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3316),
.B(n_3105),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3369),
.B(n_3281),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3318),
.B(n_3211),
.Y(n_3436)
);

OAI221xp5_ASAP7_75t_SL g3437 ( 
.A1(n_3298),
.A2(n_3276),
.B1(n_3260),
.B2(n_3274),
.C(n_3275),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3317),
.B(n_3118),
.Y(n_3438)
);

OAI221xp5_ASAP7_75t_L g3439 ( 
.A1(n_3336),
.A2(n_3115),
.B1(n_3273),
.B2(n_3272),
.C(n_3223),
.Y(n_3439)
);

NAND4xp25_ASAP7_75t_L g3440 ( 
.A(n_3335),
.B(n_3157),
.C(n_347),
.D(n_348),
.Y(n_3440)
);

AOI21xp33_ASAP7_75t_L g3441 ( 
.A1(n_3320),
.A2(n_3213),
.B(n_3212),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3383),
.B(n_3118),
.Y(n_3442)
);

OAI22xp5_ASAP7_75t_L g3443 ( 
.A1(n_3326),
.A2(n_3222),
.B1(n_3118),
.B2(n_3197),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3396),
.B(n_3381),
.Y(n_3444)
);

OAI221xp5_ASAP7_75t_L g3445 ( 
.A1(n_3303),
.A2(n_3264),
.B1(n_3129),
.B2(n_3095),
.C(n_352),
.Y(n_3445)
);

AND2x2_ASAP7_75t_L g3446 ( 
.A(n_3381),
.B(n_3095),
.Y(n_3446)
);

AND2x2_ASAP7_75t_SL g3447 ( 
.A(n_3308),
.B(n_3129),
.Y(n_3447)
);

NAND4xp25_ASAP7_75t_L g3448 ( 
.A(n_3307),
.B(n_343),
.C(n_349),
.D(n_350),
.Y(n_3448)
);

OAI21xp5_ASAP7_75t_SL g3449 ( 
.A1(n_3366),
.A2(n_3325),
.B(n_3322),
.Y(n_3449)
);

OAI21xp5_ASAP7_75t_SL g3450 ( 
.A1(n_3310),
.A2(n_3129),
.B(n_350),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3386),
.B(n_353),
.Y(n_3451)
);

AOI221xp5_ASAP7_75t_L g3452 ( 
.A1(n_3368),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.C(n_358),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3330),
.B(n_355),
.Y(n_3453)
);

NAND3xp33_ASAP7_75t_L g3454 ( 
.A(n_3398),
.B(n_356),
.C(n_358),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3389),
.B(n_359),
.Y(n_3455)
);

NAND3xp33_ASAP7_75t_L g3456 ( 
.A(n_3395),
.B(n_3297),
.C(n_3341),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3346),
.B(n_359),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3390),
.B(n_360),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3376),
.B(n_360),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3309),
.B(n_361),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3313),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_3461)
);

AND2x2_ASAP7_75t_L g3462 ( 
.A(n_3375),
.B(n_362),
.Y(n_3462)
);

OAI21xp5_ASAP7_75t_SL g3463 ( 
.A1(n_3384),
.A2(n_363),
.B(n_364),
.Y(n_3463)
);

OAI22xp5_ASAP7_75t_SL g3464 ( 
.A1(n_3314),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_3464)
);

AO21x2_ASAP7_75t_L g3465 ( 
.A1(n_3426),
.A2(n_3291),
.B(n_3331),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3431),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3404),
.B(n_3357),
.Y(n_3467)
);

NAND3xp33_ASAP7_75t_L g3468 ( 
.A(n_3449),
.B(n_3397),
.C(n_3337),
.Y(n_3468)
);

NOR3xp33_ASAP7_75t_L g3469 ( 
.A(n_3429),
.B(n_3285),
.C(n_3306),
.Y(n_3469)
);

INVx3_ASAP7_75t_L g3470 ( 
.A(n_3447),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3408),
.B(n_3302),
.Y(n_3471)
);

AO21x2_ASAP7_75t_L g3472 ( 
.A1(n_3424),
.A2(n_3363),
.B(n_3359),
.Y(n_3472)
);

NAND4xp75_ASAP7_75t_L g3473 ( 
.A(n_3447),
.B(n_3311),
.C(n_3402),
.D(n_3391),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3420),
.B(n_3422),
.Y(n_3474)
);

AOI22xp33_ASAP7_75t_L g3475 ( 
.A1(n_3440),
.A2(n_3394),
.B1(n_3385),
.B2(n_3401),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3416),
.B(n_3373),
.Y(n_3476)
);

AOI211xp5_ASAP7_75t_L g3477 ( 
.A1(n_3429),
.A2(n_3355),
.B(n_3378),
.C(n_3338),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3417),
.B(n_3345),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3419),
.B(n_3344),
.Y(n_3479)
);

NAND4xp25_ASAP7_75t_L g3480 ( 
.A(n_3407),
.B(n_3319),
.C(n_3312),
.D(n_3400),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3412),
.A2(n_3401),
.B1(n_3403),
.B2(n_3393),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3418),
.B(n_3349),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3412),
.A2(n_3403),
.B1(n_3393),
.B2(n_3392),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3421),
.B(n_3347),
.Y(n_3484)
);

NOR3xp33_ASAP7_75t_L g3485 ( 
.A(n_3407),
.B(n_3354),
.C(n_3286),
.Y(n_3485)
);

NOR2x1_ASAP7_75t_L g3486 ( 
.A(n_3450),
.B(n_3342),
.Y(n_3486)
);

AOI22xp33_ASAP7_75t_L g3487 ( 
.A1(n_3462),
.A2(n_3392),
.B1(n_3388),
.B2(n_3400),
.Y(n_3487)
);

AO21x2_ASAP7_75t_L g3488 ( 
.A1(n_3435),
.A2(n_3454),
.B(n_3436),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3444),
.B(n_3334),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3417),
.B(n_3315),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3423),
.B(n_3367),
.Y(n_3491)
);

NAND3xp33_ASAP7_75t_L g3492 ( 
.A(n_3430),
.B(n_3388),
.C(n_3399),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3425),
.Y(n_3493)
);

AO21x2_ASAP7_75t_L g3494 ( 
.A1(n_3463),
.A2(n_3356),
.B(n_3364),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3433),
.B(n_3327),
.Y(n_3495)
);

NOR3xp33_ASAP7_75t_SL g3496 ( 
.A(n_3443),
.B(n_3371),
.C(n_3332),
.Y(n_3496)
);

OR2x2_ASAP7_75t_L g3497 ( 
.A(n_3406),
.B(n_3370),
.Y(n_3497)
);

NAND4xp75_ASAP7_75t_L g3498 ( 
.A(n_3410),
.B(n_3379),
.C(n_3339),
.D(n_3353),
.Y(n_3498)
);

NOR2x1_ASAP7_75t_L g3499 ( 
.A(n_3413),
.B(n_3374),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_L g3500 ( 
.A1(n_3409),
.A2(n_3399),
.B1(n_3379),
.B2(n_3351),
.Y(n_3500)
);

AOI211xp5_ASAP7_75t_L g3501 ( 
.A1(n_3430),
.A2(n_3377),
.B(n_3361),
.C(n_3360),
.Y(n_3501)
);

OR2x2_ASAP7_75t_L g3502 ( 
.A(n_3405),
.B(n_3380),
.Y(n_3502)
);

INVxp67_ASAP7_75t_SL g3503 ( 
.A(n_3428),
.Y(n_3503)
);

OR2x2_ASAP7_75t_L g3504 ( 
.A(n_3432),
.B(n_3380),
.Y(n_3504)
);

NOR4xp75_ASAP7_75t_L g3505 ( 
.A(n_3445),
.B(n_366),
.C(n_368),
.D(n_370),
.Y(n_3505)
);

AOI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3415),
.A2(n_3343),
.B1(n_3362),
.B2(n_3328),
.Y(n_3506)
);

OA211x2_ASAP7_75t_L g3507 ( 
.A1(n_3427),
.A2(n_3456),
.B(n_3414),
.C(n_3434),
.Y(n_3507)
);

NAND3xp33_ASAP7_75t_L g3508 ( 
.A(n_3411),
.B(n_3365),
.C(n_3377),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3460),
.Y(n_3509)
);

BUFx3_ASAP7_75t_L g3510 ( 
.A(n_3446),
.Y(n_3510)
);

AOI22xp5_ASAP7_75t_L g3511 ( 
.A1(n_3459),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.Y(n_3511)
);

NOR3xp33_ASAP7_75t_SL g3512 ( 
.A(n_3468),
.B(n_3437),
.C(n_3411),
.Y(n_3512)
);

HB1xp67_ASAP7_75t_L g3513 ( 
.A(n_3503),
.Y(n_3513)
);

NAND3xp33_ASAP7_75t_L g3514 ( 
.A(n_3469),
.B(n_3448),
.C(n_3437),
.Y(n_3514)
);

NOR3xp33_ASAP7_75t_L g3515 ( 
.A(n_3492),
.B(n_3464),
.C(n_3452),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3474),
.B(n_3438),
.Y(n_3516)
);

NAND3xp33_ASAP7_75t_L g3517 ( 
.A(n_3486),
.B(n_3485),
.C(n_3496),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3474),
.B(n_3442),
.Y(n_3518)
);

OR2x2_ASAP7_75t_L g3519 ( 
.A(n_3493),
.B(n_3457),
.Y(n_3519)
);

INVx1_ASAP7_75t_SL g3520 ( 
.A(n_3510),
.Y(n_3520)
);

XOR2x2_ASAP7_75t_L g3521 ( 
.A(n_3499),
.B(n_3473),
.Y(n_3521)
);

OR2x2_ASAP7_75t_L g3522 ( 
.A(n_3493),
.B(n_3502),
.Y(n_3522)
);

XOR2x2_ASAP7_75t_L g3523 ( 
.A(n_3505),
.B(n_3439),
.Y(n_3523)
);

NAND3xp33_ASAP7_75t_L g3524 ( 
.A(n_3496),
.B(n_3477),
.C(n_3481),
.Y(n_3524)
);

NOR3xp33_ASAP7_75t_L g3525 ( 
.A(n_3480),
.B(n_3441),
.C(n_3461),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3504),
.Y(n_3526)
);

INVx3_ASAP7_75t_L g3527 ( 
.A(n_3470),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3466),
.Y(n_3528)
);

INVx1_ASAP7_75t_SL g3529 ( 
.A(n_3510),
.Y(n_3529)
);

XNOR2xp5_ASAP7_75t_L g3530 ( 
.A(n_3507),
.B(n_3453),
.Y(n_3530)
);

AOI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3483),
.A2(n_3481),
.B1(n_3484),
.B2(n_3487),
.Y(n_3531)
);

OR2x2_ASAP7_75t_L g3532 ( 
.A(n_3497),
.B(n_3451),
.Y(n_3532)
);

AOI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3483),
.A2(n_3458),
.B1(n_3455),
.B2(n_374),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_3478),
.B(n_371),
.Y(n_3534)
);

INVx1_ASAP7_75t_SL g3535 ( 
.A(n_3478),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3491),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3467),
.B(n_373),
.Y(n_3537)
);

AND2x4_ASAP7_75t_L g3538 ( 
.A(n_3470),
.B(n_374),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3467),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3482),
.B(n_376),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3471),
.B(n_376),
.Y(n_3541)
);

OR2x2_ASAP7_75t_L g3542 ( 
.A(n_3509),
.B(n_377),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3495),
.Y(n_3543)
);

XOR2x2_ASAP7_75t_L g3544 ( 
.A(n_3498),
.B(n_377),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3490),
.Y(n_3545)
);

INVx2_ASAP7_75t_SL g3546 ( 
.A(n_3470),
.Y(n_3546)
);

XNOR2xp5_ASAP7_75t_L g3547 ( 
.A(n_3509),
.B(n_378),
.Y(n_3547)
);

NAND4xp75_ASAP7_75t_L g3548 ( 
.A(n_3506),
.B(n_3479),
.C(n_3495),
.D(n_3511),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3489),
.B(n_378),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3476),
.B(n_379),
.Y(n_3550)
);

XNOR2x2_ASAP7_75t_L g3551 ( 
.A(n_3508),
.B(n_381),
.Y(n_3551)
);

XOR2x2_ASAP7_75t_L g3552 ( 
.A(n_3501),
.B(n_381),
.Y(n_3552)
);

XOR2x2_ASAP7_75t_L g3553 ( 
.A(n_3500),
.B(n_382),
.Y(n_3553)
);

INVxp67_ASAP7_75t_L g3554 ( 
.A(n_3517),
.Y(n_3554)
);

XOR2xp5_ASAP7_75t_L g3555 ( 
.A(n_3530),
.B(n_3500),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3513),
.Y(n_3556)
);

XOR2x2_ASAP7_75t_L g3557 ( 
.A(n_3524),
.B(n_3487),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3524),
.B(n_3472),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3543),
.B(n_3488),
.Y(n_3559)
);

AOI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_3514),
.A2(n_3465),
.B1(n_3472),
.B2(n_3494),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3526),
.B(n_3488),
.Y(n_3561)
);

XNOR2x1_ASAP7_75t_L g3562 ( 
.A(n_3521),
.B(n_382),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3522),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3529),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3528),
.Y(n_3565)
);

AO22x1_ASAP7_75t_L g3566 ( 
.A1(n_3529),
.A2(n_3465),
.B1(n_3494),
.B2(n_3475),
.Y(n_3566)
);

XNOR2x1_ASAP7_75t_L g3567 ( 
.A(n_3552),
.B(n_383),
.Y(n_3567)
);

INVx2_ASAP7_75t_SL g3568 ( 
.A(n_3520),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3539),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3519),
.Y(n_3570)
);

XOR2x2_ASAP7_75t_L g3571 ( 
.A(n_3517),
.B(n_3475),
.Y(n_3571)
);

XOR2x2_ASAP7_75t_L g3572 ( 
.A(n_3553),
.B(n_3523),
.Y(n_3572)
);

XNOR2x2_ASAP7_75t_L g3573 ( 
.A(n_3551),
.B(n_384),
.Y(n_3573)
);

OA22x2_ASAP7_75t_L g3574 ( 
.A1(n_3531),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_3535),
.B(n_385),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3536),
.Y(n_3576)
);

XNOR2x1_ASAP7_75t_L g3577 ( 
.A(n_3548),
.B(n_387),
.Y(n_3577)
);

INVxp67_ASAP7_75t_L g3578 ( 
.A(n_3537),
.Y(n_3578)
);

XOR2x2_ASAP7_75t_L g3579 ( 
.A(n_3531),
.B(n_390),
.Y(n_3579)
);

XNOR2xp5_ASAP7_75t_L g3580 ( 
.A(n_3512),
.B(n_390),
.Y(n_3580)
);

INVx1_ASAP7_75t_SL g3581 ( 
.A(n_3568),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3564),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3555),
.B(n_3514),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3556),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3556),
.Y(n_3585)
);

AND2x4_ASAP7_75t_L g3586 ( 
.A(n_3564),
.B(n_3527),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3576),
.Y(n_3587)
);

HB1xp67_ASAP7_75t_L g3588 ( 
.A(n_3565),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3563),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3554),
.A2(n_3525),
.B1(n_3515),
.B2(n_3535),
.Y(n_3590)
);

XOR2x2_ASAP7_75t_L g3591 ( 
.A(n_3572),
.B(n_3544),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3569),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3570),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3554),
.A2(n_3545),
.B1(n_3533),
.B2(n_3540),
.Y(n_3594)
);

OA22x2_ASAP7_75t_L g3595 ( 
.A1(n_3560),
.A2(n_3533),
.B1(n_3547),
.B2(n_3546),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3570),
.Y(n_3596)
);

AOI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3571),
.A2(n_3557),
.B1(n_3558),
.B2(n_3579),
.Y(n_3597)
);

OA22x2_ASAP7_75t_L g3598 ( 
.A1(n_3560),
.A2(n_3527),
.B1(n_3538),
.B2(n_3549),
.Y(n_3598)
);

OA22x2_ASAP7_75t_L g3599 ( 
.A1(n_3580),
.A2(n_3538),
.B1(n_3541),
.B2(n_3550),
.Y(n_3599)
);

XNOR2xp5_ASAP7_75t_L g3600 ( 
.A(n_3562),
.B(n_3534),
.Y(n_3600)
);

OA22x2_ASAP7_75t_L g3601 ( 
.A1(n_3578),
.A2(n_3518),
.B1(n_3516),
.B2(n_3532),
.Y(n_3601)
);

XNOR2x1_ASAP7_75t_L g3602 ( 
.A(n_3577),
.B(n_3542),
.Y(n_3602)
);

INVx3_ASAP7_75t_L g3603 ( 
.A(n_3573),
.Y(n_3603)
);

INVx1_ASAP7_75t_SL g3604 ( 
.A(n_3575),
.Y(n_3604)
);

INVx2_ASAP7_75t_SL g3605 ( 
.A(n_3574),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3561),
.Y(n_3606)
);

OAI22x1_ASAP7_75t_L g3607 ( 
.A1(n_3558),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_3607)
);

AO22x1_ASAP7_75t_L g3608 ( 
.A1(n_3566),
.A2(n_392),
.B1(n_393),
.B2(n_395),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3584),
.Y(n_3609)
);

INVx1_ASAP7_75t_SL g3610 ( 
.A(n_3581),
.Y(n_3610)
);

HB1xp67_ASAP7_75t_L g3611 ( 
.A(n_3582),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3596),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3588),
.Y(n_3613)
);

OA22x2_ASAP7_75t_L g3614 ( 
.A1(n_3597),
.A2(n_3578),
.B1(n_3559),
.B2(n_3567),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3589),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3587),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3592),
.Y(n_3617)
);

HB1xp67_ASAP7_75t_L g3618 ( 
.A(n_3585),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3605),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3593),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3590),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3604),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3586),
.Y(n_3623)
);

INVx8_ASAP7_75t_L g3624 ( 
.A(n_3603),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3608),
.Y(n_3625)
);

OAI322xp33_ASAP7_75t_L g3626 ( 
.A1(n_3583),
.A2(n_3574),
.A3(n_396),
.B1(n_398),
.B2(n_399),
.C1(n_400),
.C2(n_401),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3606),
.Y(n_3627)
);

INVx5_ASAP7_75t_L g3628 ( 
.A(n_3603),
.Y(n_3628)
);

INVxp67_ASAP7_75t_L g3629 ( 
.A(n_3607),
.Y(n_3629)
);

HB1xp67_ASAP7_75t_SL g3630 ( 
.A(n_3619),
.Y(n_3630)
);

OAI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3628),
.A2(n_3601),
.B1(n_3595),
.B2(n_3598),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3610),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3624),
.Y(n_3633)
);

OAI322xp33_ASAP7_75t_L g3634 ( 
.A1(n_3614),
.A2(n_3599),
.A3(n_3594),
.B1(n_3602),
.B2(n_3600),
.C1(n_3606),
.C2(n_3591),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3624),
.Y(n_3635)
);

AOI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3628),
.A2(n_3608),
.B1(n_3586),
.B2(n_400),
.Y(n_3636)
);

OAI222xp33_ASAP7_75t_L g3637 ( 
.A1(n_3628),
.A2(n_395),
.B1(n_396),
.B2(n_401),
.C1(n_403),
.C2(n_404),
.Y(n_3637)
);

INVx1_ASAP7_75t_SL g3638 ( 
.A(n_3622),
.Y(n_3638)
);

AOI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_3621),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_3639)
);

AOI22xp5_ASAP7_75t_L g3640 ( 
.A1(n_3629),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.Y(n_3640)
);

AO22x2_ASAP7_75t_L g3641 ( 
.A1(n_3625),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_3641)
);

AOI22xp5_ASAP7_75t_SL g3642 ( 
.A1(n_3613),
.A2(n_3609),
.B1(n_3615),
.B2(n_3623),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_3609),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3627),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.Y(n_3644)
);

OA22x2_ASAP7_75t_L g3645 ( 
.A1(n_3627),
.A2(n_410),
.B1(n_413),
.B2(n_414),
.Y(n_3645)
);

NAND4xp25_ASAP7_75t_L g3646 ( 
.A(n_3616),
.B(n_416),
.C(n_417),
.D(n_418),
.Y(n_3646)
);

AOI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_3631),
.A2(n_3611),
.B1(n_3617),
.B2(n_3612),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3632),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3641),
.Y(n_3649)
);

O2A1O1Ixp33_ASAP7_75t_SL g3650 ( 
.A1(n_3633),
.A2(n_3618),
.B(n_3620),
.C(n_3626),
.Y(n_3650)
);

AOI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3635),
.A2(n_3630),
.B1(n_3638),
.B2(n_3636),
.Y(n_3651)
);

AOI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3640),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_3652)
);

AOI22xp33_ASAP7_75t_L g3653 ( 
.A1(n_3634),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_3653)
);

AOI22xp5_ASAP7_75t_L g3654 ( 
.A1(n_3641),
.A2(n_420),
.B1(n_422),
.B2(n_423),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3645),
.Y(n_3655)
);

A2O1A1Ixp33_ASAP7_75t_L g3656 ( 
.A1(n_3642),
.A2(n_422),
.B(n_425),
.C(n_426),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3643),
.Y(n_3657)
);

INVxp33_ASAP7_75t_L g3658 ( 
.A(n_3646),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3639),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3644),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_SL g3661 ( 
.A1(n_3637),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_3661)
);

AOI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_3653),
.A2(n_427),
.B1(n_428),
.B2(n_430),
.Y(n_3662)
);

NOR2x1_ASAP7_75t_L g3663 ( 
.A(n_3655),
.B(n_430),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3648),
.Y(n_3664)
);

AOI22xp5_ASAP7_75t_L g3665 ( 
.A1(n_3651),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.Y(n_3665)
);

INVxp67_ASAP7_75t_L g3666 ( 
.A(n_3649),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3657),
.Y(n_3667)
);

AO22x2_ASAP7_75t_L g3668 ( 
.A1(n_3659),
.A2(n_431),
.B1(n_433),
.B2(n_434),
.Y(n_3668)
);

AOI31xp33_ASAP7_75t_L g3669 ( 
.A1(n_3658),
.A2(n_435),
.A3(n_436),
.B(n_437),
.Y(n_3669)
);

AOI221xp5_ASAP7_75t_L g3670 ( 
.A1(n_3650),
.A2(n_3660),
.B1(n_3656),
.B2(n_3647),
.C(n_3661),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3654),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3652),
.B(n_435),
.Y(n_3672)
);

AOI22xp5_ASAP7_75t_L g3673 ( 
.A1(n_3653),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3670),
.B(n_438),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3663),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3668),
.Y(n_3676)
);

AOI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_3671),
.A2(n_439),
.B1(n_441),
.B2(n_443),
.Y(n_3677)
);

AOI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3665),
.A2(n_439),
.B1(n_441),
.B2(n_444),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3667),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3664),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3669),
.Y(n_3681)
);

INVxp67_ASAP7_75t_SL g3682 ( 
.A(n_3666),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3672),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3662),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3673),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3663),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3679),
.Y(n_3687)
);

AND4x1_ASAP7_75t_L g3688 ( 
.A(n_3677),
.B(n_445),
.C(n_446),
.D(n_447),
.Y(n_3688)
);

AO22x1_ASAP7_75t_L g3689 ( 
.A1(n_3676),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_3689)
);

AOI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3681),
.A2(n_448),
.B1(n_449),
.B2(n_452),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3683),
.Y(n_3691)
);

AO22x2_ASAP7_75t_L g3692 ( 
.A1(n_3674),
.A2(n_449),
.B1(n_453),
.B2(n_454),
.Y(n_3692)
);

OAI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3684),
.A2(n_453),
.B1(n_525),
.B2(n_527),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3689),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3692),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3690),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3691),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3687),
.Y(n_3698)
);

INVxp67_ASAP7_75t_L g3699 ( 
.A(n_3697),
.Y(n_3699)
);

AO22x2_ASAP7_75t_L g3700 ( 
.A1(n_3695),
.A2(n_3682),
.B1(n_3680),
.B2(n_3685),
.Y(n_3700)
);

OAI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_3694),
.A2(n_3682),
.B1(n_3686),
.B2(n_3675),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3698),
.Y(n_3702)
);

AOI22xp5_ASAP7_75t_L g3703 ( 
.A1(n_3696),
.A2(n_3693),
.B1(n_3678),
.B2(n_3688),
.Y(n_3703)
);

XOR2xp5_ASAP7_75t_L g3704 ( 
.A(n_3703),
.B(n_3698),
.Y(n_3704)
);

INVxp67_ASAP7_75t_SL g3705 ( 
.A(n_3699),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3700),
.Y(n_3706)
);

AOI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3705),
.A2(n_3701),
.B1(n_3702),
.B2(n_531),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_3707),
.Y(n_3708)
);

AOI22x1_ASAP7_75t_L g3709 ( 
.A1(n_3708),
.A2(n_3704),
.B1(n_3706),
.B2(n_532),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3709),
.Y(n_3710)
);

AOI221xp5_ASAP7_75t_L g3711 ( 
.A1(n_3710),
.A2(n_3708),
.B1(n_529),
.B2(n_533),
.C(n_535),
.Y(n_3711)
);

AOI211xp5_ASAP7_75t_L g3712 ( 
.A1(n_3711),
.A2(n_528),
.B(n_536),
.C(n_537),
.Y(n_3712)
);


endmodule