module fake_jpeg_22311_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_55),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_24),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_53),
.B(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_18),
.B1(n_24),
.B2(n_32),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_60),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_62),
.Y(n_101)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_18),
.B1(n_32),
.B2(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_67),
.Y(n_108)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_72),
.Y(n_109)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_79),
.Y(n_116)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_33),
.B1(n_23),
.B2(n_30),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_84),
.B(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_91),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_33),
.B1(n_23),
.B2(n_30),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_66),
.B1(n_39),
.B2(n_46),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_25),
.B1(n_29),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_29),
.B1(n_21),
.B2(n_36),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_17),
.B1(n_26),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_96),
.A2(n_34),
.B1(n_22),
.B2(n_26),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_28),
.B1(n_17),
.B2(n_26),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_1),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_17),
.B(n_22),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_111),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_28),
.B1(n_21),
.B2(n_31),
.Y(n_107)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_31),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_132),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_97),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_136),
.B(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_35),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_27),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_73),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_137),
.C(n_87),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_49),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_47),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_83),
.B1(n_103),
.B2(n_112),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_85),
.B1(n_27),
.B2(n_75),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_67),
.C(n_54),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_106),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_54),
.CI(n_47),
.CON(n_140),
.SN(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_146),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_144),
.A2(n_118),
.B(n_129),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_157),
.B1(n_160),
.B2(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_75),
.B1(n_95),
.B2(n_92),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_153),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_110),
.B1(n_93),
.B2(n_104),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_129),
.B1(n_139),
.B2(n_114),
.Y(n_190)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_115),
.Y(n_151)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_87),
.B1(n_93),
.B2(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_78),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_163),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_87),
.B1(n_90),
.B2(n_79),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_112),
.A3(n_100),
.B1(n_94),
.B2(n_81),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_77),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_123),
.B(n_1),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_1),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_2),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_3),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_138),
.C(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_195),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_120),
.B(n_140),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_184),
.B(n_192),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_162),
.B1(n_158),
.B2(n_157),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_140),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_135),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_150),
.C(n_172),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_193),
.B(n_143),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_197),
.B1(n_7),
.B2(n_8),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_116),
.B(n_118),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_115),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_116),
.B(n_5),
.C(n_6),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_149),
.A2(n_130),
.B(n_95),
.C(n_114),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_199),
.B(n_113),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_130),
.B1(n_113),
.B2(n_7),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_201),
.B(n_220),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_215),
.B1(n_218),
.B2(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_162),
.B1(n_160),
.B2(n_171),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_224),
.B1(n_186),
.B2(n_196),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_163),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_209),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_206),
.A2(n_211),
.B(n_221),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_182),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_219),
.C(n_189),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_153),
.C(n_150),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_172),
.C(n_146),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_168),
.B1(n_148),
.B2(n_142),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_151),
.C(n_156),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_218)
);

XOR2x2_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_6),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_16),
.B(n_10),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_9),
.B(n_10),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_195),
.B(n_191),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_237),
.B1(n_203),
.B2(n_186),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_238),
.B1(n_221),
.B2(n_215),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_233),
.C(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_241),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_175),
.B1(n_190),
.B2(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_212),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_196),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_208),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_213),
.C(n_209),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_249),
.C(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_208),
.C(n_204),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_216),
.C(n_202),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_231),
.B(n_219),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_255),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_224),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_205),
.C(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_230),
.C(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_198),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_253),
.C(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_226),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_239),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_243),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_222),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_174),
.Y(n_278)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_273),
.B(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_245),
.C(n_244),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_242),
.B(n_256),
.C(n_226),
.D(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_232),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_270),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_262),
.B1(n_236),
.B2(n_218),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_196),
.B1(n_267),
.B2(n_260),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_286),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_273),
.B(n_272),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_274),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_199),
.B(n_176),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_282),
.B1(n_276),
.B2(n_280),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_12),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_292),
.B(n_293),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_287),
.Y(n_292)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_293),
.B(n_188),
.C(n_15),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_14),
.C(n_15),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_294),
.B1(n_14),
.B2(n_16),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_14),
.Y(n_299)
);


endmodule