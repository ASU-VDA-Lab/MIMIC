module real_jpeg_16064_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_523),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_0),
.B(n_524),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_1),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_1),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_1),
.B(n_96),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_2),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_3),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_3),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_4),
.B(n_96),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_4),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_4),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_4),
.B(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_4),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_4),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_4),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_5),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_6),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_246),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_7),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_7),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_7),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_8),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_8),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_8),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_8),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_8),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_8),
.A2(n_9),
.B1(n_279),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_9),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_9),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_9),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_9),
.B(n_490),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_10),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_11),
.B(n_63),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_11),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_11),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_11),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_11),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_11),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_11),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_11),
.B(n_449),
.Y(n_448)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_12),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_12),
.Y(n_312)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_13),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_13),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_13),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_13),
.B(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_15),
.B(n_34),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_15),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_15),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_15),
.B(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_15),
.B(n_416),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_15),
.B(n_500),
.Y(n_499)
);

BUFx4f_ASAP7_75t_L g125 ( 
.A(n_16),
.Y(n_125)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_16),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g454 ( 
.A(n_16),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_16),
.Y(n_488)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_17),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_17),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_166),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_165),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_103),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_23),
.B(n_103),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.C(n_68),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_25),
.A2(n_26),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_42),
.C(n_48),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.C(n_37),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_28),
.A2(n_29),
.B1(n_37),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_31),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_33),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_33),
.Y(n_152)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_37),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_37),
.B(n_198),
.C(n_202),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_37),
.B(n_202),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_39),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_42),
.B(n_197),
.C(n_203),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_42),
.A2(n_43),
.B1(n_203),
.B2(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_43),
.B(n_164),
.Y(n_207)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_45),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_46),
.Y(n_338)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_53),
.B(n_154),
.C(n_163),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_64),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_55),
.A2(n_56),
.B1(n_121),
.B2(n_122),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_55),
.A2(n_56),
.B1(n_298),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_121),
.C(n_126),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_56),
.B(n_298),
.C(n_300),
.Y(n_297)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_58),
.Y(n_341)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_59),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_64),
.A2(n_78),
.B1(n_142),
.B2(n_143),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_64),
.B(n_143),
.C(n_286),
.Y(n_343)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_79),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_78),
.C(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_74),
.A2(n_79),
.B1(n_225),
.B2(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_77),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_79),
.B(n_147),
.C(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_101),
.B2(n_102),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_111),
.C(n_116),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_87),
.B(n_239),
.C(n_248),
.Y(n_238)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_89),
.A2(n_248),
.B1(n_249),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_89),
.Y(n_370)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_90),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_128),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_104),
.B(n_107),
.Y(n_173)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_120),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_110),
.B(n_120),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_116),
.A2(n_147),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_119),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_122),
.B1(n_160),
.B2(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_156),
.C(n_160),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_122),
.B(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_122),
.B(n_350),
.Y(n_413)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_127),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_148),
.C(n_153),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_145),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_133),
.B(n_145),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.C(n_142),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_195)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_137),
.Y(n_301)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_137),
.Y(n_472)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AO22x1_ASAP7_75t_SL g206 ( 
.A1(n_154),
.A2(n_155),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_185),
.C(n_189),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_160),
.A2(n_161),
.B1(n_189),
.B2(n_190),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_160),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_161),
.B(n_420),
.Y(n_456)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_162),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_162),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_251),
.B(n_520),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_209),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_171),
.A2(n_521),
.B(n_522),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_172),
.B(n_174),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_179),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_177),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_196),
.C(n_206),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_181),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_194),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_182),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_184),
.B(n_194),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_186),
.B(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_189),
.A2(n_190),
.B1(n_293),
.B2(n_294),
.Y(n_317)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_190),
.B(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_191),
.Y(n_309)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_206),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);

OR2x6_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_210),
.B(n_212),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_219),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_213),
.B(n_216),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_219),
.B(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_232),
.C(n_237),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_220),
.A2(n_221),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.C(n_229),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_222),
.B(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_224),
.A2(n_229),
.B1(n_230),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_224),
.Y(n_378)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_390)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_239),
.A2(n_240),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_241),
.A2(n_245),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_241),
.Y(n_349)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_242),
.Y(n_422)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_244),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_245),
.Y(n_350)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_247),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_250),
.Y(n_418)
);

NAND2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_403),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_380),
.B(n_396),
.C(n_397),
.D(n_402),
.Y(n_252)
);

OAI21x1_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_356),
.B(n_379),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_327),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_SL g519 ( 
.A(n_255),
.B(n_327),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_288),
.C(n_313),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_256),
.B(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_268),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_257),
.B(n_269),
.C(n_285),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.C(n_263),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_258),
.B(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_411)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_285),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_275),
.B(n_278),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_278),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_288),
.A2(n_289),
.B1(n_313),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_302),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_296),
.B2(n_297),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_291),
.B(n_297),
.C(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_307),
.C(n_310),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_313),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.C(n_318),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_314),
.B(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_317),
.B(n_318),
.Y(n_409)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.C(n_325),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_319),
.B(n_325),
.Y(n_461)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_322),
.B(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_345),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_346),
.C(n_355),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_344),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_339),
.B1(n_340),
.B2(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_336),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_340),
.B(n_343),
.C(n_372),
.Y(n_371)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_342),
.Y(n_372)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_360),
.C(n_361),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_355),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_353),
.C(n_354),
.Y(n_365)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

NOR2x1_ASAP7_75t_L g518 ( 
.A(n_356),
.B(n_519),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_358),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_362),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_382),
.C(n_383),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_375),
.B2(n_376),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_371),
.B1(n_373),
.B2(n_374),
.Y(n_366)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_371),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_371),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_386),
.C(n_387),
.Y(n_385)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_376),
.Y(n_383)
);

NAND4xp25_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_397),
.C(n_404),
.D(n_518),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_384),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_392),
.B1(n_394),
.B2(n_395),
.Y(n_388)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_390),
.Y(n_391)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_394),
.C(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_400),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_426),
.B(n_517),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_423),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_406),
.B(n_423),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.C(n_412),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_407),
.A2(n_408),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_410),
.B(n_412),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.C(n_419),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_413),
.A2(n_414),
.B1(n_415),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_419),
.B(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_511),
.B(n_516),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_465),
.B(n_510),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_457),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_429),
.B(n_457),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_446),
.C(n_455),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_430),
.A2(n_431),
.B1(n_476),
.B2(n_478),
.Y(n_475)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_441),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_439),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_439),
.C(n_441),
.Y(n_459)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_446),
.A2(n_455),
.B1(n_456),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_447),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_468)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_454),
.Y(n_501)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_462),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_459),
.B(n_460),
.C(n_462),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_479),
.B(n_509),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_475),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_467),
.B(n_475),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.C(n_473),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_492),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_469),
.A2(n_470),
.B1(n_473),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_473),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_476),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_480),
.A2(n_494),
.B(n_508),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_491),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_481),
.B(n_491),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_489),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_489),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_498),
.B(n_507),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_497),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_496),
.B(n_497),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_512),
.B(n_513),
.Y(n_516)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);


endmodule