module fake_aes_2255_n_710 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_710);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_710;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_703;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_478;
wire n_442;
wire n_331;
wire n_485;
wire n_482;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_31), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_50), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_13), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_12), .Y(n_81) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_10), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_41), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_61), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_58), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_49), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_8), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_32), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_29), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_39), .Y(n_90) );
OR2x2_ASAP7_75t_L g91 ( .A(n_63), .B(n_34), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_59), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_56), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_68), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_47), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_22), .Y(n_97) );
INVx2_ASAP7_75t_SL g98 ( .A(n_60), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_53), .Y(n_99) );
BUFx10_ASAP7_75t_L g100 ( .A(n_3), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_55), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_36), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_48), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_66), .Y(n_107) );
INVx4_ASAP7_75t_R g108 ( .A(n_44), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_11), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_30), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_76), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_3), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_25), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_37), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_14), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_46), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_62), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_24), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
INVxp33_ASAP7_75t_L g124 ( .A(n_6), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_7), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_98), .B(n_0), .Y(n_127) );
AND2x6_ASAP7_75t_L g128 ( .A(n_97), .B(n_28), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_125), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_124), .A2(n_1), .B1(n_4), .B2(n_5), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_98), .B(n_5), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_104), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_125), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_104), .Y(n_138) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_113), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_113), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
AOI22xp5_ASAP7_75t_SL g143 ( .A1(n_122), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_97), .B(n_45), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_80), .B(n_15), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_83), .B(n_16), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_92), .A2(n_16), .B1(n_17), .B2(n_19), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_117), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
INVx6_ASAP7_75t_L g153 ( .A(n_120), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_90), .Y(n_155) );
BUFx8_ASAP7_75t_L g156 ( .A(n_91), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_120), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_89), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_95), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_82), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_87), .B(n_123), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_105), .B(n_17), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_106), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_109), .B(n_20), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_107), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_82), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_82), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_163), .A2(n_116), .B1(n_100), .B2(n_93), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_161), .B(n_101), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_137), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_142), .B(n_103), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_163), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_142), .B(n_121), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_163), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_165), .B(n_119), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_131), .Y(n_177) );
CKINVDCx11_ASAP7_75t_R g178 ( .A(n_132), .Y(n_178) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_155), .B(n_119), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_152), .B(n_78), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_152), .B(n_118), .Y(n_183) );
INVx6_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
NAND2xp33_ASAP7_75t_SL g185 ( .A(n_147), .B(n_92), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_155), .Y(n_186) );
OR2x2_ASAP7_75t_L g187 ( .A(n_141), .B(n_78), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_158), .B(n_86), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_165), .Y(n_190) );
NOR2x1p5_ASAP7_75t_L g191 ( .A(n_161), .B(n_86), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_165), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_156), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_161), .B(n_88), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_161), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_147), .B(n_158), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_127), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_159), .B(n_88), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_159), .B(n_100), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
NOR3xp33_ASAP7_75t_L g204 ( .A(n_129), .B(n_114), .C(n_110), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_134), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_162), .B(n_100), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_156), .B(n_111), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_128), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_128), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_128), .Y(n_212) );
OR2x6_ASAP7_75t_L g213 ( .A(n_139), .B(n_136), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_128), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_162), .B(n_111), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_137), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_128), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_137), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_128), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_164), .B(n_99), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_144), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_144), .Y(n_223) );
NOR2x1p5_ASAP7_75t_L g224 ( .A(n_146), .B(n_99), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_137), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_144), .A2(n_94), .B1(n_112), .B2(n_102), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_164), .B(n_94), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx4_ASAP7_75t_SL g229 ( .A(n_144), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_166), .B(n_112), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_151), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_203), .B(n_156), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_198), .B(n_166), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_205), .B(n_144), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_192), .A2(n_144), .B(n_151), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_192), .A2(n_126), .B(n_135), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_185), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_177), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_172), .B(n_144), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_193), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_180), .B(n_126), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_177), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_196), .B(n_143), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_173), .A2(n_130), .B1(n_135), .B2(n_138), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_196), .B(n_130), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_195), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_203), .B(n_149), .Y(n_248) );
NAND2x1_ASAP7_75t_L g249 ( .A(n_184), .B(n_108), .Y(n_249) );
BUFx2_ASAP7_75t_SL g250 ( .A(n_170), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_170), .A2(n_149), .B1(n_102), .B2(n_138), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_195), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_202), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_203), .B(n_157), .Y(n_254) );
INVx2_ASAP7_75t_SL g255 ( .A(n_187), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_202), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_207), .A2(n_168), .B1(n_160), .B2(n_140), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_181), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_189), .B(n_168), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_210), .B(n_157), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_207), .B(n_168), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_206), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_210), .B(n_157), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_182), .Y(n_265) );
OR2x6_ASAP7_75t_L g266 ( .A(n_213), .B(n_153), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_220), .B(n_160), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_210), .B(n_157), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_191), .B(n_160), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_227), .B(n_140), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_182), .Y(n_271) );
AO22x1_ASAP7_75t_L g272 ( .A1(n_186), .A2(n_140), .B1(n_167), .B2(n_154), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_200), .B(n_167), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_194), .B(n_153), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_215), .B(n_167), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_214), .B(n_167), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_231), .A2(n_153), .B1(n_167), .B2(n_154), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_214), .B(n_157), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_188), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_176), .B(n_153), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_224), .B(n_154), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_169), .B(n_154), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_187), .B(n_154), .Y(n_284) );
NOR2x1p5_ASAP7_75t_L g285 ( .A(n_193), .B(n_21), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_211), .Y(n_286) );
O2A1O1Ixp5_ASAP7_75t_L g287 ( .A1(n_214), .A2(n_23), .B(n_26), .C(n_33), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_201), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_175), .B(n_35), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_197), .B(n_38), .Y(n_290) );
NAND2xp33_ASAP7_75t_SL g291 ( .A(n_226), .B(n_40), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_185), .Y(n_292) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_219), .B(n_42), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_190), .B(n_52), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_184), .A2(n_54), .B1(n_57), .B2(n_64), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_SL g296 ( .A1(n_174), .A2(n_65), .B(n_67), .C(n_69), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_190), .B(n_70), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_206), .Y(n_298) );
NAND2xp33_ASAP7_75t_L g299 ( .A(n_221), .B(n_72), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_184), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_239), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_234), .B(n_190), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_286), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_253), .B(n_208), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_250), .A2(n_178), .B1(n_204), .B2(n_184), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_244), .A2(n_178), .B1(n_213), .B2(n_183), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_235), .A2(n_219), .B(n_223), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_246), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_293), .B(n_219), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_256), .B(n_179), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_238), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_255), .B(n_222), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_239), .Y(n_314) );
OAI22x1_ASAP7_75t_L g315 ( .A1(n_251), .A2(n_186), .B1(n_213), .B2(n_222), .Y(n_315) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_293), .B(n_223), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_248), .A2(n_213), .B1(n_232), .B2(n_206), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_236), .A2(n_223), .B(n_221), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_266), .B(n_229), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_286), .B(n_221), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_269), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_266), .B(n_201), .Y(n_322) );
NOR2xp33_ASAP7_75t_SL g323 ( .A(n_292), .B(n_217), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_266), .A2(n_217), .B1(n_211), .B2(n_212), .Y(n_324) );
NOR2xp33_ASAP7_75t_SL g325 ( .A(n_300), .B(n_212), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_245), .A2(n_230), .B1(n_228), .B2(n_209), .C(n_232), .Y(n_326) );
NOR2xp33_ASAP7_75t_R g327 ( .A(n_291), .B(n_221), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_263), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_286), .B(n_221), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_242), .A2(n_232), .B(n_218), .C(n_199), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_240), .A2(n_229), .B(n_199), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_269), .B(n_233), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_245), .B(n_229), .Y(n_334) );
OAI21xp33_ASAP7_75t_L g335 ( .A1(n_247), .A2(n_229), .B(n_216), .Y(n_335) );
INVxp33_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_286), .B(n_171), .Y(n_337) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_287), .A2(n_216), .B(n_218), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_257), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_243), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_243), .B(n_77), .Y(n_341) );
OAI21xp33_ASAP7_75t_SL g342 ( .A1(n_262), .A2(n_225), .B(n_171), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_258), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_233), .B(n_225), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_258), .B(n_171), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_285), .Y(n_346) );
NOR3xp33_ASAP7_75t_SL g347 ( .A(n_274), .B(n_171), .C(n_280), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_294), .A2(n_171), .B(n_297), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_265), .A2(n_252), .B1(n_282), .B2(n_279), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_265), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_254), .A2(n_278), .B(n_264), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_271), .B(n_288), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_SL g353 ( .A1(n_310), .A2(n_296), .B(n_290), .C(n_289), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_309), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_298), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_333), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_308), .A2(n_268), .B(n_278), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_348), .A2(n_268), .B(n_254), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_311), .A2(n_283), .B(n_259), .C(n_281), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_SL g361 ( .A1(n_310), .A2(n_296), .B(n_275), .C(n_273), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_331), .A2(n_260), .B(n_264), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_237), .B(n_260), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_318), .A2(n_276), .B(n_249), .Y(n_364) );
AO31x2_ASAP7_75t_L g365 ( .A1(n_349), .A2(n_280), .A3(n_267), .B(n_270), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g366 ( .A1(n_316), .A2(n_263), .B1(n_298), .B2(n_274), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_352), .A2(n_277), .B(n_295), .C(n_299), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_301), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_317), .B(n_295), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_306), .A2(n_272), .B1(n_315), .B2(n_305), .Y(n_370) );
NAND3xp33_ASAP7_75t_SL g371 ( .A(n_312), .B(n_317), .C(n_332), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_337), .A2(n_341), .B(n_338), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_304), .B(n_339), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_302), .A2(n_334), .B(n_325), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_314), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_322), .B(n_350), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_330), .B(n_332), .C(n_344), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_320), .A2(n_329), .B(n_344), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_328), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_346), .B(n_321), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_307), .A2(n_326), .B1(n_336), .B2(n_319), .C(n_328), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_319), .A2(n_324), .B1(n_345), .B2(n_347), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_303), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_342), .A2(n_347), .B(n_335), .C(n_323), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_377), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_372), .A2(n_337), .B(n_320), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_353), .A2(n_338), .B(n_329), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_370), .A2(n_303), .B1(n_338), .B2(n_327), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_373), .A2(n_303), .B(n_327), .C(n_378), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_373), .B(n_303), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_356), .A2(n_371), .B1(n_355), .B2(n_354), .Y(n_394) );
BUFx8_ASAP7_75t_L g395 ( .A(n_375), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_374), .A2(n_359), .B(n_379), .Y(n_396) );
AO21x2_ASAP7_75t_L g397 ( .A1(n_378), .A2(n_385), .B(n_367), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_384), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_384), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_367), .A2(n_385), .B(n_369), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_380), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_357), .B(n_365), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_380), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_365), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_365), .B(n_382), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_363), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_360), .B(n_383), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_358), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_381), .A2(n_361), .B1(n_353), .B2(n_366), .C(n_364), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_381), .B(n_361), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_385), .B(n_367), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_402), .B(n_406), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_395), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_402), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_388), .A2(n_392), .B(n_409), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_390), .B(n_406), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_404), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_394), .A2(n_406), .B1(n_395), .B2(n_409), .Y(n_424) );
AOI21x1_ASAP7_75t_L g425 ( .A1(n_388), .A2(n_389), .B(n_412), .Y(n_425) );
AO21x2_ASAP7_75t_L g426 ( .A1(n_392), .A2(n_389), .B(n_410), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_386), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g428 ( .A1(n_394), .A2(n_412), .B(n_411), .C(n_401), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_404), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_408), .A2(n_405), .B1(n_407), .B2(n_393), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_407), .A2(n_393), .B(n_410), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_408), .B(n_405), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_408), .A2(n_401), .B1(n_405), .B2(n_403), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_391), .B(n_405), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_405), .B(n_400), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_403), .B(n_398), .Y(n_439) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_411), .A2(n_399), .B(n_398), .C(n_404), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_395), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_395), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_396), .A2(n_397), .B(n_413), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_397), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_396), .A2(n_397), .B(n_413), .Y(n_446) );
OAI211xp5_ASAP7_75t_SL g447 ( .A1(n_399), .A2(n_395), .B(n_397), .C(n_413), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_387), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_436), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_423), .Y(n_451) );
NAND2x1_ASAP7_75t_L g452 ( .A(n_415), .B(n_387), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_397), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_442), .Y(n_454) );
OAI221xp5_ASAP7_75t_SL g455 ( .A1(n_424), .A2(n_403), .B1(n_413), .B2(n_399), .C(n_400), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_414), .B(n_413), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_421), .B(n_400), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_414), .B(n_400), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_416), .B(n_400), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_416), .B(n_400), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_417), .B(n_399), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_436), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_445), .B(n_387), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_417), .B(n_387), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_445), .B(n_387), .Y(n_466) );
NOR2x1_ASAP7_75t_L g467 ( .A(n_415), .B(n_387), .Y(n_467) );
AOI21xp5_ASAP7_75t_SL g468 ( .A1(n_442), .A2(n_435), .B(n_431), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_435), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_419), .A2(n_425), .B(n_440), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_421), .B(n_420), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_423), .Y(n_476) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_415), .B(n_441), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
BUFx2_ASAP7_75t_SL g479 ( .A(n_442), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_418), .B(n_427), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_430), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_415), .B(n_441), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_427), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_434), .B(n_443), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_443), .B(n_432), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_420), .B(n_433), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_444), .B(n_446), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_439), .B(n_432), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_433), .B(n_437), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_438), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_441), .B(n_428), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_444), .B(n_446), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_444), .B(n_446), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_439), .B(n_446), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_438), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_480), .B(n_428), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_473), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_492), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_473), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_458), .B(n_446), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_458), .B(n_444), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_477), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_458), .B(n_444), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_484), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_494), .B(n_419), .C(n_447), .D(n_431), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_454), .B(n_447), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_492), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_453), .B(n_426), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_453), .B(n_426), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_456), .B(n_426), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_462), .B(n_426), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_456), .B(n_449), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_484), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_497), .B(n_449), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_479), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_451), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_451), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_489), .B(n_449), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_497), .B(n_425), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_490), .B(n_448), .Y(n_526) );
INVx3_ASAP7_75t_R g527 ( .A(n_479), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_475), .Y(n_528) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_496), .B(n_422), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_480), .Y(n_530) );
NOR2xp33_ASAP7_75t_R g531 ( .A(n_483), .B(n_448), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_454), .B(n_440), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_490), .B(n_422), .Y(n_533) );
BUFx4f_ASAP7_75t_SL g534 ( .A(n_454), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_469), .A2(n_422), .B1(n_491), .B2(n_463), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_452), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_491), .B(n_422), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_491), .B(n_422), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_462), .B(n_422), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_474), .B(n_485), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_464), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_464), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_471), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_450), .B(n_487), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_477), .B(n_481), .C(n_471), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_475), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_481), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_499), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_491), .B(n_466), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_466), .B(n_450), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_466), .B(n_465), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_489), .B(n_495), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_487), .B(n_474), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_499), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_465), .B(n_493), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_493), .B(n_461), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_534), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_524), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_544), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_553), .B(n_495), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_503), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_553), .B(n_496), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_521), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_553), .B(n_457), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_553), .B(n_457), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_505), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_524), .Y(n_571) );
AOI211xp5_ASAP7_75t_SL g572 ( .A1(n_512), .A2(n_468), .B(n_455), .C(n_489), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_505), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_531), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_552), .B(n_495), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_532), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_510), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_519), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_545), .B(n_459), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_530), .B(n_461), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_552), .B(n_463), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_506), .B(n_463), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_545), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_519), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_530), .B(n_459), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_554), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_554), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_539), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_539), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_542), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_542), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_551), .B(n_460), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_551), .B(n_460), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_546), .B(n_498), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_541), .B(n_498), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_506), .B(n_469), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_558), .B(n_486), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_501), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_549), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_543), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_501), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_529), .B(n_508), .Y(n_606) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_546), .B(n_468), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_507), .B(n_463), .Y(n_608) );
AND2x2_ASAP7_75t_SL g609 ( .A(n_527), .B(n_476), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_507), .B(n_467), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_543), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_509), .B(n_467), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_586), .B(n_509), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_562), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_594), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g616 ( .A(n_565), .B(n_508), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_595), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_590), .B(n_502), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_606), .B(n_529), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_604), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_560), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_611), .Y(n_622) );
AOI21xp33_ASAP7_75t_SL g623 ( .A1(n_609), .A2(n_527), .B(n_517), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_591), .B(n_558), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_592), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_593), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_609), .A2(n_455), .B1(n_498), .B2(n_535), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_579), .B(n_526), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_565), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_576), .B(n_526), .Y(n_630) );
OR4x1_ASAP7_75t_L g631 ( .A(n_574), .B(n_548), .C(n_452), .D(n_556), .Y(n_631) );
AOI322xp5_ASAP7_75t_SL g632 ( .A1(n_575), .A2(n_550), .A3(n_525), .B1(n_515), .B2(n_516), .C1(n_514), .C2(n_520), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_607), .A2(n_599), .B1(n_610), .B2(n_612), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_576), .B(n_514), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_584), .B(n_550), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_574), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_563), .A2(n_511), .B(n_515), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_577), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_584), .B(n_533), .Y(n_639) );
AOI32xp33_ASAP7_75t_L g640 ( .A1(n_572), .A2(n_525), .A3(n_516), .B1(n_520), .B2(n_533), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_596), .B(n_518), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_567), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_577), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_603), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_568), .A2(n_569), .B1(n_600), .B2(n_597), .Y(n_645) );
AOI311xp33_ASAP7_75t_L g646 ( .A1(n_601), .A2(n_548), .A3(n_559), .B(n_557), .C(n_556), .Y(n_646) );
NAND2x1_ASAP7_75t_L g647 ( .A(n_606), .B(n_536), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_568), .A2(n_517), .B1(n_540), .B2(n_549), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_569), .A2(n_511), .B1(n_536), .B2(n_540), .Y(n_649) );
AOI211x1_ASAP7_75t_L g650 ( .A1(n_637), .A2(n_598), .B(n_563), .C(n_612), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_629), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_640), .B(n_598), .C(n_600), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_632), .A2(n_582), .B1(n_589), .B2(n_583), .C(n_588), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_621), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_615), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
NAND3x1_ASAP7_75t_L g657 ( .A(n_633), .B(n_610), .C(n_608), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_642), .B(n_608), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g659 ( .A1(n_634), .A2(n_585), .A3(n_518), .B1(n_580), .B2(n_581), .C1(n_564), .C2(n_566), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_646), .B(n_603), .C(n_582), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_617), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_628), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_636), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_613), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_639), .B(n_585), .Y(n_666) );
OAI32xp33_ASAP7_75t_L g667 ( .A1(n_645), .A2(n_596), .A3(n_597), .B1(n_573), .B2(n_578), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_627), .A2(n_606), .B1(n_536), .B2(n_573), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_616), .B(n_578), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_620), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_645), .A2(n_570), .B1(n_561), .B2(n_571), .C(n_555), .Y(n_671) );
INVxp67_ASAP7_75t_SL g672 ( .A(n_649), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_651), .Y(n_673) );
AOI321xp33_ASAP7_75t_L g674 ( .A1(n_653), .A2(n_627), .A3(n_648), .B1(n_623), .B2(n_618), .C(n_619), .Y(n_674) );
AOI222xp33_ASAP7_75t_L g675 ( .A1(n_652), .A2(n_648), .B1(n_625), .B2(n_626), .C1(n_622), .C2(n_619), .Y(n_675) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_672), .A2(n_630), .A3(n_624), .B1(n_635), .B2(n_638), .C1(n_643), .C2(n_644), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_660), .A2(n_537), .B1(n_538), .B2(n_561), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_661), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_659), .B(n_571), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_668), .A2(n_647), .A3(n_537), .B1(n_538), .B2(n_631), .C1(n_557), .C2(n_555), .Y(n_680) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_668), .A2(n_513), .A3(n_504), .B1(n_605), .B2(n_602), .C1(n_587), .C2(n_486), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_657), .A2(n_513), .B(n_504), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_671), .B(n_605), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_671), .B(n_602), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_654), .A2(n_536), .B(n_472), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_650), .A2(n_587), .B1(n_536), .B2(n_547), .C(n_528), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_677), .A2(n_667), .B1(n_656), .B2(n_663), .C(n_661), .Y(n_687) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_677), .A2(n_656), .B1(n_665), .B2(n_658), .C1(n_655), .C2(n_670), .Y(n_688) );
NAND3xp33_ASAP7_75t_SL g689 ( .A(n_674), .B(n_662), .C(n_666), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_685), .B(n_664), .C(n_669), .Y(n_690) );
A2O1A1O1Ixp25_ASAP7_75t_L g691 ( .A1(n_679), .A2(n_669), .B(n_472), .C(n_470), .D(n_522), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_676), .B(n_472), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_678), .A2(n_547), .B1(n_528), .B2(n_523), .C(n_522), .Y(n_693) );
INVxp67_ASAP7_75t_L g694 ( .A(n_673), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_689), .A2(n_680), .B(n_681), .C(n_682), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_694), .Y(n_696) );
NOR4xp25_ASAP7_75t_L g697 ( .A(n_692), .B(n_684), .C(n_683), .D(n_675), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_688), .A2(n_686), .B(n_470), .C(n_523), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_698), .A2(n_690), .B1(n_687), .B2(n_693), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_696), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_695), .B(n_691), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_700), .B(n_697), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_701), .Y(n_703) );
XNOR2x1_ASAP7_75t_L g704 ( .A(n_703), .B(n_699), .Y(n_704) );
AO22x2_ASAP7_75t_L g705 ( .A1(n_702), .A2(n_470), .B1(n_475), .B2(n_476), .Y(n_705) );
AOI22x1_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_702), .B1(n_470), .B2(n_476), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_706), .B(n_704), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_472), .B(n_478), .Y(n_708) );
OA21x2_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_478), .B(n_482), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_709), .A2(n_478), .B1(n_482), .B2(n_488), .Y(n_710) );
endmodule