module fake_jpeg_24556_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_31),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_31),
.B1(n_21),
.B2(n_22),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_48),
.B1(n_62),
.B2(n_68),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_52),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_57),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_20),
.B(n_25),
.C(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_66),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_27),
.B1(n_25),
.B2(n_29),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_6),
.C(n_7),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_26),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_26),
.B1(n_4),
.B2(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_86),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_95),
.B1(n_99),
.B2(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_3),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_3),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_6),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_7),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_116),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_94),
.C(n_87),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_85),
.C(n_101),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_93),
.B1(n_92),
.B2(n_78),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_117),
.B1(n_121),
.B2(n_125),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_52),
.A3(n_67),
.B1(n_55),
.B2(n_56),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_67),
.B1(n_59),
.B2(n_58),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_67),
.B(n_8),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_59),
.B1(n_12),
.B2(n_10),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_7),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_9),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_77),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_8),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_97),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_79),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_9),
.B1(n_15),
.B2(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_139),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_85),
.C(n_72),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_146),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_79),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_76),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_107),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_113),
.B1(n_117),
.B2(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_120),
.B(n_124),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_141),
.B(n_137),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_127),
.B(n_115),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_156),
.B(n_109),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_127),
.B(n_115),
.C(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_132),
.B(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_123),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_103),
.B1(n_126),
.B2(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_118),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_132),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_167),
.A2(n_175),
.B(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_134),
.C(n_138),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_173),
.C(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_179),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_133),
.B(n_146),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_180),
.B(n_155),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_133),
.C(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_162),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_182),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_156),
.B1(n_161),
.B2(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

AOI321xp33_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_163),
.A3(n_175),
.B1(n_150),
.B2(n_154),
.C(n_159),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_152),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_176),
.C(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_157),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_200),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_169),
.B(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_206),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_195),
.B1(n_192),
.B2(n_169),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_203),
.B1(n_186),
.B2(n_159),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_151),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_208),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_182),
.B(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_205),
.C(n_183),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_183),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_194),
.C(n_181),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_211),
.B(n_166),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_217),
.B1(n_194),
.B2(n_106),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_142),
.Y(n_219)
);


endmodule