module fake_jpeg_18605_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_0),
.CON(n_42),
.SN(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_44),
.Y(n_66)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_46),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_1),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_33),
.B1(n_22),
.B2(n_23),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_57),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_22),
.B(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_73),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_28),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_47),
.B1(n_19),
.B2(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_94),
.B1(n_71),
.B2(n_35),
.Y(n_128)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_87),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_19),
.B1(n_30),
.B2(n_47),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_86),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_91),
.B(n_17),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_34),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_32),
.B1(n_25),
.B2(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_52),
.B1(n_66),
.B2(n_54),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_52),
.B1(n_72),
.B2(n_65),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_68),
.B(n_28),
.Y(n_119)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_R g103 ( 
.A(n_67),
.B(n_24),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_17),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_15),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_67),
.B(n_70),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_105),
.B(n_77),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_124),
.B1(n_89),
.B2(n_2),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_49),
.B1(n_53),
.B2(n_48),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_113),
.B1(n_123),
.B2(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_49),
.B1(n_53),
.B2(n_60),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_78),
.B1(n_104),
.B2(n_99),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_49),
.B1(n_58),
.B2(n_51),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_79),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_100),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_118),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_49),
.B1(n_74),
.B2(n_71),
.Y(n_123)
);

OAI22x1_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_68),
.B1(n_34),
.B2(n_35),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_35),
.B1(n_17),
.B2(n_3),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_99),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_76),
.A2(n_1),
.B(n_2),
.Y(n_133)
);

AO22x2_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_78),
.B1(n_101),
.B2(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_138),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_143),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_100),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_146),
.B(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_154),
.B1(n_129),
.B2(n_113),
.Y(n_168)
);

XOR2x2_ASAP7_75t_SL g143 ( 
.A(n_124),
.B(n_92),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_R g172 ( 
.A(n_144),
.B(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_107),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_155),
.Y(n_175)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_95),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_108),
.A2(n_1),
.B(n_4),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_121),
.B1(n_109),
.B2(n_133),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_144),
.B1(n_146),
.B2(n_137),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_176),
.B1(n_136),
.B2(n_138),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_126),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_121),
.C(n_125),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_164),
.C(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_190),
.C(n_196),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_164),
.B(n_181),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_194),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_158),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_137),
.C(n_146),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_145),
.B1(n_136),
.B2(n_143),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_130),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_123),
.C(n_110),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_178),
.C(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_201),
.B(n_214),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_180),
.B1(n_173),
.B2(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_210),
.B1(n_189),
.B2(n_185),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_167),
.C(n_171),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_211),
.C(n_184),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_165),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_163),
.C(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

OAI322xp33_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_172),
.A3(n_176),
.B1(n_170),
.B2(n_166),
.C1(n_162),
.C2(n_153),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_170),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_190),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_192),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_222),
.B(n_215),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_193),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_211),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_138),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_200),
.B1(n_166),
.B2(n_138),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_205),
.B1(n_203),
.B2(n_8),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_5),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_229),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_216),
.A2(n_203),
.B1(n_14),
.B2(n_11),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_14),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_231),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_219),
.A2(n_221),
.B1(n_220),
.B2(n_217),
.Y(n_231)
);

AOI21x1_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_8),
.B(n_9),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_238),
.C(n_229),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_5),
.B(n_6),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_10),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_5),
.B(n_6),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_10),
.B(n_227),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.C(n_242),
.Y(n_243)
);

INVxp33_ASAP7_75t_SL g241 ( 
.A(n_233),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_237),
.B(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_235),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_231),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_244),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_247),
.Y(n_250)
);


endmodule