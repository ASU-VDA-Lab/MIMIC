module fake_jpeg_31667_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_62),
.Y(n_69)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_54),
.B1(n_56),
.B2(n_44),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_76),
.B1(n_78),
.B2(n_3),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_71),
.B(n_73),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_24),
.B(n_28),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_54),
.C(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_48),
.B1(n_47),
.B2(n_51),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_75),
.A2(n_61),
.B1(n_21),
.B2(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_20),
.B1(n_41),
.B2(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_82),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_19),
.A3(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_15),
.B1(n_34),
.B2(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_4),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_9),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_102),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_103),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_31),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_101),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_42),
.C(n_30),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_87),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_27),
.C(n_25),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_116)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_23),
.C(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_111),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_9),
.B(n_10),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_98),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_124),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_109),
.B(n_102),
.C(n_100),
.D(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_112),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_112),
.B1(n_123),
.B2(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_118),
.Y(n_130)
);

AOI211xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_117),
.B(n_126),
.C(n_119),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_113),
.C(n_106),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_104),
.Y(n_133)
);


endmodule