module real_aes_8770_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_385;
wire n_214;
wire n_275;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_314;
wire n_252;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_516;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g452 ( .A(n_0), .Y(n_452) );
INVx1_ASAP7_75t_L g545 ( .A(n_1), .Y(n_545) );
INVx1_ASAP7_75t_L g159 ( .A(n_2), .Y(n_159) );
AOI222xp33_ASAP7_75t_L g458 ( .A1(n_3), .A2(n_459), .B1(n_743), .B2(n_744), .C1(n_753), .C2(n_755), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_4), .A2(n_39), .B1(n_184), .B2(n_491), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g191 ( .A1(n_5), .A2(n_175), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_6), .B(n_173), .Y(n_557) );
AND2x6_ASAP7_75t_L g152 ( .A(n_7), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_8), .A2(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g110 ( .A(n_9), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_9), .B(n_40), .Y(n_453) );
INVx1_ASAP7_75t_L g197 ( .A(n_10), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_11), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_13), .B(n_165), .Y(n_500) );
INVx1_ASAP7_75t_L g268 ( .A(n_14), .Y(n_268) );
INVx1_ASAP7_75t_L g539 ( .A(n_15), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_16), .B(n_140), .Y(n_528) );
AO32x2_ASAP7_75t_L g512 ( .A1(n_17), .A2(n_139), .A3(n_173), .B1(n_493), .B2(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_18), .B(n_184), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_19), .B(n_180), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_20), .B(n_140), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_21), .A2(n_50), .B1(n_184), .B2(n_491), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_22), .B(n_175), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_23), .A2(n_100), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_23), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g492 ( .A1(n_24), .A2(n_77), .B1(n_165), .B2(n_184), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_25), .B(n_184), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_26), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_27), .A2(n_266), .B(n_267), .C(n_269), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_28), .B(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_30), .B(n_170), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_31), .B(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_32), .A2(n_90), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_32), .Y(n_130) );
INVx1_ASAP7_75t_L g212 ( .A(n_33), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_34), .B(n_170), .Y(n_484) );
INVx2_ASAP7_75t_L g150 ( .A(n_35), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_36), .B(n_184), .Y(n_561) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_37), .A2(n_70), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_37), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_37), .B(n_170), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_38), .A2(n_152), .B(n_155), .C(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_40), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g210 ( .A(n_41), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_42), .B(n_163), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_43), .B(n_184), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_44), .A2(n_88), .B1(n_232), .B2(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_45), .B(n_184), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_46), .B(n_184), .Y(n_540) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_47), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_48), .B(n_544), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_49), .B(n_175), .Y(n_256) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_51), .A2(n_62), .B1(n_165), .B2(n_184), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_52), .A2(n_748), .B1(n_749), .B2(n_752), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_52), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_53), .A2(n_155), .B1(n_165), .B2(n_208), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_54), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_55), .B(n_184), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_56), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_57), .B(n_184), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_58), .A2(n_183), .B(n_195), .C(n_196), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_59), .Y(n_245) );
INVx1_ASAP7_75t_L g193 ( .A(n_60), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_61), .A2(n_105), .B1(n_117), .B2(n_759), .Y(n_104) );
INVx1_ASAP7_75t_L g153 ( .A(n_63), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_64), .B(n_184), .Y(n_546) );
INVx1_ASAP7_75t_L g143 ( .A(n_65), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_66), .Y(n_122) );
AO32x2_ASAP7_75t_L g488 ( .A1(n_67), .A2(n_173), .A3(n_248), .B1(n_489), .B2(n_493), .Y(n_488) );
INVx1_ASAP7_75t_L g564 ( .A(n_68), .Y(n_564) );
INVx1_ASAP7_75t_L g479 ( .A(n_69), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_70), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_71), .A2(n_180), .B(n_181), .C(n_183), .Y(n_179) );
INVxp67_ASAP7_75t_L g182 ( .A(n_72), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_73), .B(n_165), .Y(n_480) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_75), .Y(n_215) );
INVx1_ASAP7_75t_L g238 ( .A(n_76), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_78), .A2(n_152), .B(n_155), .C(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_79), .B(n_491), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_80), .B(n_165), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_81), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_81), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_82), .B(n_160), .Y(n_228) );
INVx2_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_84), .B(n_180), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_85), .B(n_165), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_86), .A2(n_152), .B(n_155), .C(n_158), .Y(n_154) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g449 ( .A(n_87), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g462 ( .A(n_87), .B(n_451), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_89), .A2(n_103), .B1(n_165), .B2(n_166), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_90), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_91), .B(n_170), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_92), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_93), .A2(n_152), .B(n_155), .C(n_251), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_94), .Y(n_258) );
INVx1_ASAP7_75t_L g178 ( .A(n_95), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_96), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_97), .B(n_160), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_98), .B(n_165), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_99), .B(n_173), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_100), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_101), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_102), .A2(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g759 ( .A(n_107), .Y(n_759) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g466 ( .A(n_113), .B(n_451), .Y(n_466) );
NOR2x2_ASAP7_75t_L g757 ( .A(n_113), .B(n_450), .Y(n_757) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_457), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g758 ( .A(n_121), .Y(n_758) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_446), .B(n_454), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_128), .B1(n_444), .B2(n_445), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_125), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_128), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
INVx1_ASAP7_75t_L g463 ( .A(n_132), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_132), .A2(n_464), .B1(n_468), .B2(n_754), .Y(n_753) );
NAND2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_360), .Y(n_132) );
NOR5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_283), .C(n_315), .D(n_330), .E(n_347), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_199), .B(n_220), .C(n_271), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_171), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_136), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_136), .B(n_335), .Y(n_398) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_137), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_137), .B(n_217), .Y(n_284) );
AND2x2_ASAP7_75t_L g325 ( .A(n_137), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_137), .B(n_294), .Y(n_329) );
OR2x2_ASAP7_75t_L g366 ( .A(n_137), .B(n_205), .Y(n_366) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g204 ( .A(n_138), .B(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g274 ( .A(n_138), .Y(n_274) );
OR2x2_ASAP7_75t_L g437 ( .A(n_138), .B(n_277), .Y(n_437) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_167), .Y(n_138) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_139), .A2(n_206), .B(n_214), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_139), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g233 ( .A(n_139), .Y(n_233) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_141), .B(n_142), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_154), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g206 ( .A1(n_147), .A2(n_185), .B1(n_207), .B2(n_213), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_147), .A2(n_238), .B(n_239), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AND2x4_ASAP7_75t_L g175 ( .A(n_148), .B(n_152), .Y(n_175) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g544 ( .A(n_149), .Y(n_544) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx3_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
INVx4_ASAP7_75t_SL g185 ( .A(n_152), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_152), .A2(n_478), .B(n_481), .Y(n_477) );
BUFx3_ASAP7_75t_L g493 ( .A(n_152), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_152), .A2(n_498), .B(n_502), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_152), .A2(n_538), .B(n_542), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_152), .A2(n_551), .B(n_554), .Y(n_550) );
INVx5_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
BUFx3_ASAP7_75t_L g232 ( .A(n_156), .Y(n_232) );
INVx1_ASAP7_75t_L g491 ( .A(n_156), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .C(n_164), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_SL g478 ( .A1(n_160), .A2(n_183), .B(n_479), .C(n_480), .Y(n_478) );
INVx2_ASAP7_75t_L g515 ( .A(n_160), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_160), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_160), .A2(n_561), .B(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_161), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_161), .B(n_197), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_161), .A2(n_163), .B1(n_490), .B2(n_492), .Y(n_489) );
INVx2_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
INVx4_ASAP7_75t_L g254 ( .A(n_163), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_163), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_163), .A2(n_515), .B1(n_531), .B2(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_164), .A2(n_539), .B(n_540), .C(n_541), .Y(n_538) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_169), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_169), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g248 ( .A(n_170), .Y(n_248) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_170), .A2(n_261), .B(n_270), .Y(n_260) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_170), .A2(n_477), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_170), .A2(n_497), .B(n_505), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_171), .A2(n_340), .B1(n_341), .B2(n_344), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_171), .B(n_274), .Y(n_423) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_189), .Y(n_171) );
AND2x2_ASAP7_75t_L g219 ( .A(n_172), .B(n_205), .Y(n_219) );
AND2x2_ASAP7_75t_L g276 ( .A(n_172), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g281 ( .A(n_172), .Y(n_281) );
INVx3_ASAP7_75t_L g294 ( .A(n_172), .Y(n_294) );
OR2x2_ASAP7_75t_L g314 ( .A(n_172), .B(n_277), .Y(n_314) );
AND2x2_ASAP7_75t_L g333 ( .A(n_172), .B(n_190), .Y(n_333) );
BUFx2_ASAP7_75t_L g365 ( .A(n_172), .Y(n_365) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_186), .Y(n_172) );
INVx4_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_173), .A2(n_550), .B(n_557), .Y(n_549) );
BUFx2_ASAP7_75t_L g262 ( .A(n_175), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_185), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_177), .A2(n_185), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_177), .A2(n_185), .B(n_264), .C(n_265), .Y(n_263) );
INVx1_ASAP7_75t_L g501 ( .A(n_180), .Y(n_501) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_184), .Y(n_255) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_187), .A2(n_191), .B(n_198), .Y(n_190) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_SL g234 ( .A(n_188), .B(n_235), .Y(n_234) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_188), .B(n_493), .C(n_530), .Y(n_529) );
AO21x1_ASAP7_75t_L g619 ( .A1(n_188), .A2(n_530), .B(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g280 ( .A(n_189), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g203 ( .A(n_190), .Y(n_203) );
INVx2_ASAP7_75t_L g218 ( .A(n_190), .Y(n_218) );
OR2x2_ASAP7_75t_L g296 ( .A(n_190), .B(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_L g326 ( .A(n_190), .B(n_205), .Y(n_326) );
AND2x2_ASAP7_75t_L g343 ( .A(n_190), .B(n_274), .Y(n_343) );
AND2x2_ASAP7_75t_L g383 ( .A(n_190), .B(n_294), .Y(n_383) );
AND2x2_ASAP7_75t_SL g419 ( .A(n_190), .B(n_219), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_195), .A2(n_503), .B(n_504), .Y(n_502) );
O2A1O1Ixp5_ASAP7_75t_L g563 ( .A1(n_195), .A2(n_543), .B(n_564), .C(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp33_ASAP7_75t_SL g200 ( .A(n_201), .B(n_216), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_202), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g357 ( .A1(n_203), .A2(n_219), .B(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_203), .B(n_205), .Y(n_413) );
AND2x2_ASAP7_75t_L g349 ( .A(n_204), .B(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g277 ( .A(n_205), .Y(n_277) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_205), .Y(n_375) );
OAI22xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_208) );
INVx2_ASAP7_75t_L g211 ( .A(n_209), .Y(n_211) );
INVx4_ASAP7_75t_L g266 ( .A(n_209), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_216), .B(n_274), .Y(n_442) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_217), .A2(n_385), .B1(n_386), .B2(n_391), .Y(n_384) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x2_ASAP7_75t_L g275 ( .A(n_218), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g313 ( .A(n_218), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g350 ( .A(n_218), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_219), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g404 ( .A(n_219), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_246), .Y(n_221) );
INVx4_ASAP7_75t_L g290 ( .A(n_222), .Y(n_290) );
AND2x2_ASAP7_75t_L g368 ( .A(n_222), .B(n_335), .Y(n_368) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
INVx3_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
AND2x2_ASAP7_75t_L g301 ( .A(n_223), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g305 ( .A(n_223), .Y(n_305) );
INVx2_ASAP7_75t_L g319 ( .A(n_223), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_223), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g376 ( .A(n_223), .B(n_371), .Y(n_376) );
AND2x2_ASAP7_75t_L g441 ( .A(n_223), .B(n_411), .Y(n_441) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_234), .Y(n_223) );
AOI21xp5_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_226), .B(n_233), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_230), .A2(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g269 ( .A(n_232), .Y(n_269) );
INVx1_ASAP7_75t_L g243 ( .A(n_233), .Y(n_243) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_233), .A2(n_537), .B(n_547), .Y(n_536) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_233), .A2(n_559), .B(n_566), .Y(n_558) );
AND2x2_ASAP7_75t_L g282 ( .A(n_236), .B(n_260), .Y(n_282) );
INVx2_ASAP7_75t_L g302 ( .A(n_236), .Y(n_302) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_243), .B(n_244), .Y(n_236) );
INVx1_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
AND2x2_ASAP7_75t_L g353 ( .A(n_246), .B(n_301), .Y(n_353) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_259), .Y(n_246) );
INVx2_ASAP7_75t_L g292 ( .A(n_247), .Y(n_292) );
INVx1_ASAP7_75t_L g300 ( .A(n_247), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_247), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_247), .B(n_302), .Y(n_356) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_257), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_256), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_255), .Y(n_251) );
AND2x2_ASAP7_75t_L g335 ( .A(n_259), .B(n_292), .Y(n_335) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
AND2x2_ASAP7_75t_L g371 ( .A(n_260), .B(n_302), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_266), .B(n_268), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_266), .A2(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g541 ( .A(n_266), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_278), .B(n_282), .Y(n_271) );
INVx1_ASAP7_75t_SL g316 ( .A(n_272), .Y(n_316) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_273), .B(n_280), .Y(n_373) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g322 ( .A(n_274), .B(n_277), .Y(n_322) );
AND2x2_ASAP7_75t_L g351 ( .A(n_274), .B(n_295), .Y(n_351) );
OR2x2_ASAP7_75t_L g354 ( .A(n_274), .B(n_314), .Y(n_354) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_275), .A2(n_367), .B1(n_419), .B2(n_420), .C1(n_422), .C2(n_424), .Y(n_418) );
BUFx2_ASAP7_75t_L g332 ( .A(n_277), .Y(n_332) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g321 ( .A(n_280), .B(n_322), .Y(n_321) );
INVx3_ASAP7_75t_SL g338 ( .A(n_280), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_280), .B(n_332), .Y(n_392) );
AND2x2_ASAP7_75t_L g327 ( .A(n_282), .B(n_287), .Y(n_327) );
INVx1_ASAP7_75t_L g346 ( .A(n_282), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_285), .B1(n_289), .B2(n_293), .C(n_297), .Y(n_283) );
OR2x2_ASAP7_75t_L g355 ( .A(n_285), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g340 ( .A(n_287), .B(n_310), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_287), .B(n_300), .Y(n_380) );
AND2x2_ASAP7_75t_L g385 ( .A(n_287), .B(n_335), .Y(n_385) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_287), .Y(n_395) );
NAND2x1_ASAP7_75t_SL g406 ( .A(n_287), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g291 ( .A(n_288), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_288), .B(n_306), .Y(n_337) );
INVx1_ASAP7_75t_L g403 ( .A(n_288), .Y(n_403) );
INVx1_ASAP7_75t_L g378 ( .A(n_289), .Y(n_378) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g390 ( .A(n_290), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g402 ( .A(n_290), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g407 ( .A(n_291), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_291), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g310 ( .A(n_292), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_292), .B(n_302), .Y(n_323) );
INVx1_ASAP7_75t_L g389 ( .A(n_292), .Y(n_389) );
INVx1_ASAP7_75t_L g410 ( .A(n_293), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_303), .B(n_312), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g443 ( .A(n_299), .B(n_376), .Y(n_443) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g411 ( .A(n_300), .B(n_371), .Y(n_411) );
AOI32xp33_ASAP7_75t_L g324 ( .A1(n_301), .A2(n_307), .A3(n_325), .B1(n_327), .B2(n_328), .Y(n_324) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_301), .A2(n_333), .A3(n_416), .B1(n_427), .B2(n_428), .C1(n_429), .C2(n_431), .Y(n_426) );
INVx2_ASAP7_75t_L g306 ( .A(n_302), .Y(n_306) );
INVx1_ASAP7_75t_L g416 ( .A(n_302), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B1(n_308), .B2(n_309), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_304), .B(n_310), .Y(n_359) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_305), .B(n_371), .Y(n_421) );
INVx1_ASAP7_75t_L g308 ( .A(n_306), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_306), .B(n_335), .Y(n_425) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_314), .B(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_317), .B1(n_320), .B2(n_323), .C(n_324), .Y(n_315) );
OR2x2_ASAP7_75t_L g336 ( .A(n_317), .B(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g345 ( .A(n_317), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g370 ( .A(n_318), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g374 ( .A(n_328), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_336), .B2(n_338), .C(n_339), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_332), .A2(n_363), .B1(n_367), .B2(n_368), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_333), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_333), .Y(n_438) );
INVx1_ASAP7_75t_L g432 ( .A(n_335), .Y(n_432) );
INVx1_ASAP7_75t_SL g367 ( .A(n_336), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_338), .B(n_366), .Y(n_428) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_343), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g409 ( .A(n_343), .Y(n_409) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
OAI221xp5_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_352), .B1(n_354), .B2(n_355), .C(n_357), .Y(n_347) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_349), .A2(n_367), .B1(n_413), .B2(n_414), .Y(n_412) );
CKINVDCx14_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_354), .A2(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR3xp33_ASAP7_75t_SL g360 ( .A(n_361), .B(n_393), .C(n_417), .Y(n_360) );
NAND4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_369), .C(n_377), .D(n_384), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g440 ( .A(n_365), .Y(n_440) );
INVx3_ASAP7_75t_SL g434 ( .A(n_366), .Y(n_434) );
OR2x2_ASAP7_75t_L g439 ( .A(n_366), .B(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B1(n_374), .B2(n_376), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_371), .B(n_389), .Y(n_430) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_379), .B(n_381), .Y(n_377) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_396), .B(n_399), .C(n_412), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g427 ( .A(n_398), .Y(n_427) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_404), .B1(n_405), .B2(n_408), .C1(n_410), .C2(n_411), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND4xp25_ASAP7_75t_SL g436 ( .A(n_409), .B(n_437), .C(n_438), .D(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_426), .C(n_435), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_435) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g456 ( .A(n_449), .Y(n_456) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g457 ( .A1(n_454), .A2(n_458), .B(n_758), .Y(n_457) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_464), .B2(n_467), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g754 ( .A(n_461), .Y(n_754) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_664), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_613), .C(n_655), .Y(n_469) );
AOI211xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_522), .B(n_567), .C(n_589), .Y(n_470) );
OAI211xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_485), .B(n_506), .C(n_517), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_473), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g676 ( .A(n_473), .B(n_593), .Y(n_676) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g578 ( .A(n_474), .B(n_509), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_474), .B(n_496), .Y(n_695) );
INVx1_ASAP7_75t_L g713 ( .A(n_474), .Y(n_713) );
AND2x2_ASAP7_75t_L g722 ( .A(n_474), .B(n_610), .Y(n_722) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g605 ( .A(n_475), .B(n_496), .Y(n_605) );
AND2x2_ASAP7_75t_L g663 ( .A(n_475), .B(n_610), .Y(n_663) );
INVx1_ASAP7_75t_L g707 ( .A(n_475), .Y(n_707) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g584 ( .A(n_476), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g592 ( .A(n_476), .Y(n_592) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_476), .Y(n_632) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_494), .Y(n_486) );
AND2x2_ASAP7_75t_L g571 ( .A(n_487), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g604 ( .A(n_487), .Y(n_604) );
OR2x2_ASAP7_75t_L g730 ( .A(n_487), .B(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_487), .B(n_496), .Y(n_734) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g509 ( .A(n_488), .Y(n_509) );
INVx1_ASAP7_75t_L g520 ( .A(n_488), .Y(n_520) );
AND2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_511), .Y(n_593) );
AND2x2_ASAP7_75t_L g633 ( .A(n_488), .B(n_512), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_493), .A2(n_560), .B(n_563), .Y(n_559) );
INVxp67_ASAP7_75t_L g675 ( .A(n_494), .Y(n_675) );
AND2x4_ASAP7_75t_L g700 ( .A(n_494), .B(n_593), .Y(n_700) );
BUFx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_495), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g510 ( .A(n_496), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g579 ( .A(n_496), .B(n_512), .Y(n_579) );
INVx1_ASAP7_75t_L g585 ( .A(n_496), .Y(n_585) );
INVx2_ASAP7_75t_L g611 ( .A(n_496), .Y(n_611) );
AND2x2_ASAP7_75t_L g627 ( .A(n_496), .B(n_628), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_507), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g582 ( .A(n_509), .Y(n_582) );
AND2x2_ASAP7_75t_L g690 ( .A(n_509), .B(n_511), .Y(n_690) );
AND2x2_ASAP7_75t_L g607 ( .A(n_510), .B(n_592), .Y(n_607) );
AND2x2_ASAP7_75t_L g706 ( .A(n_510), .B(n_707), .Y(n_706) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_511), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g731 ( .A(n_511), .B(n_592), .Y(n_731) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g521 ( .A(n_512), .Y(n_521) );
AND2x2_ASAP7_75t_L g610 ( .A(n_512), .B(n_611), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_515), .A2(n_543), .B(n_545), .C(n_546), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_515), .A2(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
AND2x2_ASAP7_75t_L g656 ( .A(n_519), .B(n_591), .Y(n_656) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_520), .B(n_592), .Y(n_641) );
INVx2_ASAP7_75t_L g640 ( .A(n_521), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_521), .A2(n_584), .B1(n_645), .B2(n_647), .C1(n_648), .C2(n_651), .Y(n_644) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_533), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g569 ( .A(n_526), .Y(n_569) );
OR2x2_ASAP7_75t_L g680 ( .A(n_526), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g602 ( .A(n_527), .Y(n_602) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_527), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g659 ( .A(n_527), .B(n_573), .Y(n_659) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g620 ( .A(n_528), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_533), .A2(n_623), .B1(n_662), .B2(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_548), .Y(n_533) );
INVx3_ASAP7_75t_L g595 ( .A(n_534), .Y(n_595) );
OR2x2_ASAP7_75t_L g728 ( .A(n_534), .B(n_604), .Y(n_728) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g617 ( .A(n_535), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g625 ( .A(n_535), .B(n_573), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_535), .B(n_549), .Y(n_681) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g572 ( .A(n_536), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g576 ( .A(n_536), .B(n_549), .Y(n_576) );
AND2x2_ASAP7_75t_L g652 ( .A(n_536), .B(n_599), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_536), .B(n_558), .Y(n_692) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_548), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g608 ( .A(n_548), .B(n_569), .Y(n_608) );
AND2x2_ASAP7_75t_L g612 ( .A(n_548), .B(n_602), .Y(n_612) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_558), .Y(n_548) );
INVx3_ASAP7_75t_L g573 ( .A(n_549), .Y(n_573) );
AND2x2_ASAP7_75t_L g598 ( .A(n_549), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g733 ( .A(n_549), .B(n_716), .Y(n_733) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_558), .Y(n_587) );
INVx2_ASAP7_75t_L g599 ( .A(n_558), .Y(n_599) );
AND2x2_ASAP7_75t_L g643 ( .A(n_558), .B(n_619), .Y(n_643) );
INVx1_ASAP7_75t_L g686 ( .A(n_558), .Y(n_686) );
OR2x2_ASAP7_75t_L g717 ( .A(n_558), .B(n_619), .Y(n_717) );
AND2x2_ASAP7_75t_L g737 ( .A(n_558), .B(n_573), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_574), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g575 ( .A(n_569), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_569), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g694 ( .A(n_571), .Y(n_694) );
INVx2_ASAP7_75t_SL g588 ( .A(n_572), .Y(n_588) );
AND2x2_ASAP7_75t_L g708 ( .A(n_572), .B(n_602), .Y(n_708) );
INVx2_ASAP7_75t_L g654 ( .A(n_573), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_573), .B(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B1(n_580), .B2(n_586), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_576), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g742 ( .A(n_576), .Y(n_742) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g667 ( .A(n_578), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_578), .B(n_610), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_579), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g683 ( .A(n_579), .B(n_632), .Y(n_683) );
INVx2_ASAP7_75t_L g739 ( .A(n_579), .Y(n_739) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_L g609 ( .A(n_582), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_582), .B(n_627), .Y(n_660) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_584), .B(n_604), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g721 ( .A(n_587), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_SL g671 ( .A1(n_588), .A2(n_672), .B(n_674), .C(n_677), .Y(n_671) );
OR2x2_ASAP7_75t_L g698 ( .A(n_588), .B(n_602), .Y(n_698) );
OAI221xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_594), .B1(n_596), .B2(n_603), .C(n_606), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_591), .B(n_640), .Y(n_647) );
AND2x2_ASAP7_75t_L g689 ( .A(n_591), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g725 ( .A(n_591), .Y(n_725) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_592), .Y(n_616) );
INVx1_ASAP7_75t_L g629 ( .A(n_592), .Y(n_629) );
NOR2xp67_ASAP7_75t_L g649 ( .A(n_595), .B(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g703 ( .A(n_595), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_595), .B(n_643), .Y(n_719) );
INVx2_ASAP7_75t_L g705 ( .A(n_596), .Y(n_705) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g646 ( .A(n_598), .B(n_617), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_598), .A2(n_614), .B(n_656), .C(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g624 ( .A(n_599), .B(n_619), .Y(n_624) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_603), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OR2x2_ASAP7_75t_L g672 ( .A(n_604), .B(n_673), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_609), .B2(n_612), .Y(n_606) );
INVx1_ASAP7_75t_L g726 ( .A(n_608), .Y(n_726) );
INVx1_ASAP7_75t_L g673 ( .A(n_610), .Y(n_673) );
INVx1_ASAP7_75t_L g724 ( .A(n_612), .Y(n_724) );
AOI211xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_617), .B(n_621), .C(n_644), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g636 ( .A(n_616), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g687 ( .A(n_617), .Y(n_687) );
AND2x2_ASAP7_75t_L g736 ( .A(n_617), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_626), .B(n_634), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx2_ASAP7_75t_L g650 ( .A(n_624), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_624), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g642 ( .A(n_625), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g718 ( .A(n_625), .Y(n_718) );
OAI32xp33_ASAP7_75t_L g729 ( .A1(n_625), .A2(n_677), .A3(n_684), .B1(n_725), .B2(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_SL g626 ( .A(n_627), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_SL g697 ( .A(n_627), .Y(n_697) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g637 ( .A(n_633), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B(n_642), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g709 ( .A1(n_636), .A2(n_684), .B1(n_710), .B2(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_640), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g677 ( .A(n_643), .Y(n_677) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g670 ( .A(n_654), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_663), .A2(n_705), .B1(n_706), .B2(n_708), .C(n_709), .Y(n_704) );
NAND5xp2_ASAP7_75t_L g664 ( .A(n_665), .B(n_688), .C(n_704), .D(n_714), .E(n_732), .Y(n_664) );
AOI211xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_668), .B(n_671), .C(n_678), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g735 ( .A(n_672), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_684), .Y(n_678) );
INVx1_ASAP7_75t_SL g711 ( .A(n_681), .Y(n_711) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI322xp33_ASAP7_75t_L g693 ( .A1(n_684), .A2(n_694), .A3(n_695), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_699), .Y(n_693) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g696 ( .A(n_686), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_686), .B(n_711), .Y(n_710) );
AOI211xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_691), .B(n_693), .C(n_701), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_697), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g740 ( .A(n_707), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_722), .B1(n_723), .B2(n_727), .C(n_729), .Y(n_714) );
OAI211xp5_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_718), .B(n_719), .C(n_720), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g741 ( .A(n_717), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B1(n_735), .B2(n_736), .C(n_738), .Y(n_732) );
AOI21xp33_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_740), .B(n_741), .Y(n_738) );
CKINVDCx16_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
CKINVDCx16_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx3_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
endmodule