module fake_ariane_3053_n_140 (n_8, n_56, n_60, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_47, n_18, n_32, n_28, n_37, n_58, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_59, n_31, n_42, n_57, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_61, n_35, n_10, n_54, n_25, n_140);

input n_8;
input n_56;
input n_60;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_58;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_59;
input n_31;
input n_42;
input n_57;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_61;
input n_35;
input n_10;
input n_54;
input n_25;

output n_140;

wire n_83;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_120;
wire n_106;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_100;
wire n_132;
wire n_62;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_128;
wire n_105;
wire n_82;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_94;
wire n_101;
wire n_134;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_108;
wire n_102;
wire n_125;
wire n_81;
wire n_87;
wire n_136;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_63;
wire n_99;
wire n_127;

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_29),
.B(n_1),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_45),
.B1(n_35),
.B2(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_36),
.B1(n_53),
.B2(n_33),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_13),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_28),
.A2(n_5),
.B1(n_56),
.B2(n_32),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_3),
.A2(n_43),
.B1(n_59),
.B2(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_38),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_46),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_15),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_42),
.A2(n_10),
.B1(n_20),
.B2(n_44),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_0),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_6),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_9),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_92),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_12),
.B(n_16),
.Y(n_105)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_23),
.C(n_24),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_37),
.B1(n_48),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_78),
.B1(n_68),
.B2(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_97),
.B(n_108),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_87),
.B(n_79),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_76),
.B(n_83),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_72),
.B1(n_64),
.B2(n_65),
.C(n_63),
.Y(n_114)
);

AO31x2_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_86),
.A3(n_91),
.B(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_80),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_109),
.B(n_104),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_110),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_96),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_128),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_123),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_131),
.Y(n_134)
);

NAND4xp25_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_106),
.C(n_107),
.D(n_112),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_120),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_88),
.B1(n_86),
.B2(n_113),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_137),
.B(n_105),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_80),
.B(n_82),
.C(n_67),
.Y(n_140)
);


endmodule