module fake_netlist_1_9358_n_656 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_656);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_656;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g76 ( .A(n_62), .Y(n_76) );
INVxp33_ASAP7_75t_L g77 ( .A(n_67), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_46), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_71), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_66), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_7), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_52), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_40), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_45), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_17), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_29), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_61), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_50), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_35), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_58), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_0), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_38), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_68), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_74), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_56), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_23), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_37), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_69), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_3), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_72), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_8), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_6), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_49), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_10), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_60), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_32), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_20), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_33), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_22), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_15), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_7), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_81), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_102), .B(n_0), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_102), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_92), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_76), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_111), .B(n_1), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_78), .B(n_34), .Y(n_132) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_78), .A2(n_31), .B(n_70), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_77), .B(n_1), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_85), .B(n_2), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_98), .B(n_4), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_98), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_109), .B(n_4), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_107), .B(n_5), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_99), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_107), .A2(n_5), .B1(n_8), .B2(n_9), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_86), .A2(n_41), .B(n_64), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_97), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
INVx6_ASAP7_75t_L g150 ( .A(n_117), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_88), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_93), .B(n_11), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_101), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_106), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_104), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_105), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_110), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_112), .B(n_13), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_119), .Y(n_160) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_120), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_79), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_162), .B(n_95), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_139), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_162), .B(n_95), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_124), .B(n_79), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_150), .B(n_83), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_134), .A2(n_96), .B1(n_90), .B2(n_115), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_150), .B(n_103), .Y(n_172) );
NAND2xp33_ASAP7_75t_L g173 ( .A(n_132), .B(n_89), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_156), .B(n_103), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_150), .B(n_108), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
AO22x2_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_121), .B1(n_16), .B2(n_14), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_136), .B(n_118), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_150), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_137), .B(n_118), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_143), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_137), .B(n_113), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_161), .B(n_113), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_147), .B(n_148), .Y(n_188) );
INVx1_ASAP7_75t_SL g189 ( .A(n_134), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_139), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_147), .B(n_116), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_140), .A2(n_116), .B1(n_108), .B2(n_94), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_152), .B(n_94), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_148), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_157), .B(n_123), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_145), .B(n_84), .Y(n_198) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_140), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_140), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_138), .B(n_87), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_127), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_157), .B(n_87), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_138), .B(n_84), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_152), .A2(n_83), .B1(n_16), .B2(n_19), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_159), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_159), .A2(n_18), .B1(n_21), .B2(n_25), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_125), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
INVxp33_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_145), .B(n_27), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_127), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_125), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_132), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_181), .A2(n_155), .B1(n_154), .B2(n_153), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_196), .B(n_153), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_195), .B(n_154), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_209), .B(n_151), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_189), .A2(n_144), .B1(n_155), .B2(n_149), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_211), .Y(n_224) );
AND2x6_ASAP7_75t_SL g225 ( .A(n_166), .B(n_122), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_183), .B(n_122), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_194), .B(n_126), .Y(n_227) );
INVx1_ASAP7_75t_SL g228 ( .A(n_187), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_183), .B(n_126), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_203), .Y(n_230) );
NAND3xp33_ASAP7_75t_L g231 ( .A(n_193), .B(n_127), .C(n_129), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_199), .Y(n_232) );
NAND2xp33_ASAP7_75t_L g233 ( .A(n_203), .B(n_132), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_192), .B(n_130), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_192), .B(n_130), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_204), .B(n_128), .Y(n_236) );
INVxp67_ASAP7_75t_SL g237 ( .A(n_199), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_181), .A2(n_149), .B1(n_128), .B2(n_142), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_204), .B(n_135), .Y(n_239) );
NOR2xp33_ASAP7_75t_SL g240 ( .A(n_178), .B(n_132), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_181), .A2(n_149), .B1(n_132), .B2(n_160), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_174), .B(n_135), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_186), .B(n_142), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g244 ( .A1(n_177), .A2(n_133), .B1(n_146), .B2(n_160), .Y(n_244) );
NAND2xp33_ASAP7_75t_L g245 ( .A(n_203), .B(n_149), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_181), .A2(n_149), .B1(n_160), .B2(n_129), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_169), .B(n_160), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_166), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_215), .B(n_146), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_169), .B(n_160), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_178), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_172), .B(n_129), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_172), .B(n_129), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_201), .B(n_129), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_181), .A2(n_127), .B1(n_36), .B2(n_39), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_216), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_180), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_213), .B(n_127), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_213), .B(n_28), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_215), .B(n_42), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_201), .B(n_43), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_194), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g265 ( .A(n_180), .B(n_44), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_164), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_173), .A2(n_47), .B(n_48), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_217), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_165), .B(n_51), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_184), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_177), .B(n_57), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_193), .B(n_59), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_218), .B(n_63), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_185), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_165), .B(n_75), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_167), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_198), .B(n_188), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_SL g278 ( .A1(n_240), .A2(n_188), .B(n_179), .C(n_210), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_264), .B(n_184), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_264), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_274), .Y(n_281) );
AOI21xp33_ASAP7_75t_L g282 ( .A1(n_272), .A2(n_214), .B(n_210), .Y(n_282) );
AOI21xp33_ASAP7_75t_L g283 ( .A1(n_263), .A2(n_163), .B(n_191), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_220), .B(n_206), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_274), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_228), .B(n_171), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g287 ( .A1(n_249), .A2(n_206), .B(n_175), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_233), .A2(n_200), .B(n_218), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_271), .A2(n_205), .B1(n_179), .B2(n_170), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_SL g290 ( .A1(n_250), .A2(n_168), .B(n_182), .C(n_176), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_277), .A2(n_208), .B(n_202), .C(n_177), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_L g292 ( .A1(n_271), .A2(n_208), .B(n_202), .C(n_190), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_271), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_276), .A2(n_197), .B(n_176), .C(n_190), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_232), .B(n_197), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_252), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_244), .B(n_197), .C(n_164), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
CKINVDCx14_ASAP7_75t_R g301 ( .A(n_252), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_227), .Y(n_302) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_263), .B(n_197), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_259), .Y(n_304) );
NAND2xp33_ASAP7_75t_SL g305 ( .A(n_261), .B(n_207), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_230), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_263), .B(n_207), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_232), .B(n_212), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_233), .A2(n_212), .B(n_230), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_222), .A2(n_255), .B1(n_259), .B2(n_231), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_SL g311 ( .A1(n_250), .A2(n_275), .B(n_269), .C(n_273), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_222), .B(n_225), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_242), .A2(n_222), .B(n_235), .C(n_229), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_221), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_247), .A2(n_245), .B(n_254), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_226), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_224), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_255), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_223), .B(n_234), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_245), .A2(n_253), .B(n_248), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_268), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_237), .B(n_236), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_239), .A2(n_243), .B(n_251), .C(n_255), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_318), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_317), .B(n_219), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_299), .A2(n_267), .B(n_265), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_289), .A2(n_238), .B1(n_265), .B2(n_241), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_313), .B(n_246), .Y(n_329) );
OAI21x1_ASAP7_75t_SL g330 ( .A1(n_289), .A2(n_270), .B(n_256), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g331 ( .A1(n_293), .A2(n_262), .B1(n_273), .B2(n_257), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_311), .A2(n_262), .B(n_266), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_315), .B(n_257), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_316), .A2(n_266), .B(n_260), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_SL g335 ( .A1(n_278), .A2(n_260), .B(n_282), .C(n_296), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_290), .A2(n_288), .B(n_309), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_322), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_279), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_321), .A2(n_307), .B(n_283), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
AO32x2_ASAP7_75t_L g343 ( .A1(n_291), .A2(n_292), .A3(n_295), .B1(n_282), .B2(n_310), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_304), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_SL g345 ( .A1(n_283), .A2(n_307), .B(n_324), .C(n_320), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_284), .B(n_303), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_323), .A2(n_287), .B(n_297), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_286), .A2(n_312), .B1(n_319), .B2(n_298), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_279), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_305), .A2(n_314), .B(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_308), .A2(n_294), .B(n_280), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_281), .B(n_285), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_SL g354 ( .A1(n_294), .A2(n_308), .B(n_300), .C(n_306), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_326), .A2(n_301), .B(n_300), .Y(n_355) );
INVx4_ASAP7_75t_SL g356 ( .A(n_338), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_325), .B(n_314), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_338), .Y(n_358) );
AO31x2_ASAP7_75t_L g359 ( .A1(n_336), .A2(n_314), .A3(n_328), .B(n_329), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_333), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_333), .B(n_344), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_339), .B(n_346), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_345), .A2(n_335), .B(n_332), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_339), .B(n_346), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_341), .B(n_350), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_331), .A2(n_334), .B(n_330), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_344), .B(n_337), .Y(n_368) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_327), .A2(n_330), .B(n_347), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_340), .B(n_349), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_342), .A2(n_352), .B(n_351), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_354), .A2(n_342), .B(n_351), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_348), .A2(n_340), .B1(n_349), .B2(n_353), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_343), .A2(n_313), .B(n_271), .C(n_291), .Y(n_374) );
CKINVDCx11_ASAP7_75t_R g375 ( .A(n_343), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_343), .B(n_317), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_343), .A2(n_341), .B(n_327), .Y(n_377) );
AO21x2_ASAP7_75t_L g378 ( .A1(n_343), .A2(n_341), .B(n_299), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_344), .B(n_271), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_360), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g382 ( .A1(n_374), .A2(n_379), .B(n_367), .C(n_376), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_362), .B(n_376), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_364), .A2(n_366), .B(n_371), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_361), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_378), .A2(n_366), .B(n_372), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_365), .B1(n_373), .B2(n_355), .C(n_368), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_361), .B(n_379), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_377), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_377), .Y(n_393) );
OA21x2_ASAP7_75t_L g394 ( .A1(n_371), .A2(n_357), .B(n_377), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_377), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_357), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
INVx3_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_370), .B(n_368), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_356), .B(n_370), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_378), .B(n_369), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_378), .B(n_369), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_359), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_359), .A2(n_369), .B(n_375), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_369), .B(n_359), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_356), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_358), .Y(n_408) );
OA21x2_ASAP7_75t_L g409 ( .A1(n_359), .A2(n_380), .B(n_358), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_356), .B(n_362), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_356), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_367), .A2(n_364), .B(n_374), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_367), .A2(n_364), .B(n_374), .Y(n_413) );
INVx5_ASAP7_75t_SL g414 ( .A(n_400), .Y(n_414) );
AO21x2_ASAP7_75t_L g415 ( .A1(n_406), .A2(n_401), .B(n_389), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_393), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_405), .Y(n_417) );
INVx2_ASAP7_75t_SL g418 ( .A(n_411), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_393), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_405), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_381), .B(n_386), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_392), .B(n_383), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_392), .B(n_383), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_392), .B(n_383), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_384), .B(n_408), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_395), .B(n_403), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_384), .B(n_408), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_386), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_391), .B(n_388), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_403), .B(n_400), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_406), .A2(n_401), .B(n_389), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
INVxp33_ASAP7_75t_L g434 ( .A(n_410), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_409), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_391), .B(n_410), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_399), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_403), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_411), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_390), .B(n_399), .C(n_382), .D(n_387), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_402), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_387), .B(n_402), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_409), .B(n_402), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_394), .B(n_404), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_390), .A2(n_410), .B1(n_398), .B2(n_396), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_394), .B(n_404), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_404), .B(n_382), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_398), .A2(n_396), .B1(n_397), .B2(n_400), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_409), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_389), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_400), .B(n_398), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_398), .B(n_397), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_423), .B(n_409), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_419), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_423), .B(n_404), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_419), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_423), .B(n_404), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_424), .B(n_409), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_421), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_424), .B(n_389), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
AND2x4_ASAP7_75t_SL g470 ( .A(n_456), .B(n_400), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_424), .B(n_389), .Y(n_471) );
AND2x4_ASAP7_75t_SL g472 ( .A(n_456), .B(n_407), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_433), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_425), .B(n_412), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_425), .B(n_412), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_425), .B(n_412), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_444), .B(n_412), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_442), .B(n_412), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_442), .B(n_413), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_413), .Y(n_482) );
NOR4xp25_ASAP7_75t_SL g483 ( .A(n_454), .B(n_411), .C(n_407), .D(n_413), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_436), .B(n_398), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_436), .B(n_407), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_422), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_443), .B(n_413), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_416), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_431), .B(n_413), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_443), .B(n_385), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_418), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_443), .B(n_385), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_420), .Y(n_493) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_421), .B(n_385), .C(n_455), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_427), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_430), .B(n_385), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_430), .B(n_385), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_422), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_444), .B(n_385), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_418), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_426), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_417), .B(n_428), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_426), .B(n_428), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_418), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_437), .B(n_445), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_427), .B(n_431), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_427), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_440), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_435), .B(n_445), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_414), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_439), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_431), .B(n_451), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_440), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_471), .B(n_447), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_501), .B(n_434), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_503), .B(n_449), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_467), .A2(n_452), .B1(n_441), .B2(n_454), .C(n_451), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_472), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_471), .B(n_447), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_503), .B(n_435), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_495), .B(n_447), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_472), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_495), .B(n_451), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_463), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_512), .B(n_452), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_512), .B(n_452), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_458), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_486), .B(n_457), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_461), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_505), .B(n_446), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_463), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_491), .B(n_440), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_469), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_506), .B(n_431), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_491), .Y(n_539) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_510), .B(n_441), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_505), .B(n_446), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_506), .B(n_450), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_486), .B(n_457), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_461), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_476), .B(n_448), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_448), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_477), .B(n_448), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_477), .B(n_450), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_474), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_462), .B(n_450), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_459), .B(n_432), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_498), .B(n_453), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_498), .B(n_438), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_459), .B(n_415), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_462), .B(n_415), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_464), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_502), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_489), .B(n_456), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_507), .B(n_438), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_489), .B(n_456), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_518), .B(n_502), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_560), .B(n_465), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_558), .B(n_487), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_558), .B(n_487), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_514), .B(n_465), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_523), .B(n_466), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_529), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_532), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_520), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_532), .Y(n_573) );
AOI21xp33_ASAP7_75t_SL g574 ( .A1(n_524), .A2(n_510), .B(n_513), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_520), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_540), .A2(n_466), .B1(n_414), .B2(n_475), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_524), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_542), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_535), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_561), .B(n_500), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_561), .B(n_500), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_539), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_534), .B(n_510), .Y(n_583) );
NOR2xp33_ASAP7_75t_SL g584 ( .A(n_534), .B(n_513), .Y(n_584) );
OAI32xp33_ASAP7_75t_L g585 ( .A1(n_554), .A2(n_509), .A3(n_508), .B1(n_504), .B2(n_475), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_535), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_523), .B(n_470), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_516), .A2(n_482), .B1(n_480), .B2(n_479), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_521), .B(n_542), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_536), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_514), .B(n_482), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_536), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_537), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_525), .B(n_509), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_519), .B(n_480), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_517), .A2(n_479), .B1(n_490), .B2(n_492), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_537), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_519), .B(n_492), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_589), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_594), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_576), .A2(n_534), .B1(n_563), .B2(n_561), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_576), .A2(n_534), .B1(n_563), .B2(n_554), .Y(n_604) );
AOI322xp5_ASAP7_75t_L g605 ( .A1(n_596), .A2(n_525), .A3(n_527), .B1(n_528), .B2(n_515), .C1(n_553), .C2(n_547), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_574), .A2(n_557), .B1(n_414), .B2(n_468), .Y(n_606) );
XOR2x2_ASAP7_75t_L g607 ( .A(n_587), .B(n_538), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_584), .A2(n_563), .B1(n_470), .B2(n_414), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_575), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_582), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_588), .B(n_528), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_579), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_566), .B(n_527), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_570), .B(n_556), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_564), .A2(n_546), .B1(n_547), .B2(n_549), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_584), .A2(n_557), .B1(n_562), .B2(n_555), .C(n_559), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_586), .Y(n_617) );
OAI22xp33_ASAP7_75t_SL g618 ( .A1(n_577), .A2(n_499), .B1(n_478), .B2(n_468), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g619 ( .A(n_583), .B(n_414), .Y(n_619) );
AO22x1_ASAP7_75t_L g620 ( .A1(n_580), .A2(n_538), .B1(n_543), .B2(n_553), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_566), .B(n_549), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_620), .A2(n_585), .B(n_580), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_605), .B(n_567), .Y(n_623) );
O2A1O1Ixp5_ASAP7_75t_SL g624 ( .A1(n_610), .A2(n_599), .B(n_590), .C(n_597), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_602), .A2(n_581), .B(n_598), .Y(n_625) );
OAI31xp33_ASAP7_75t_L g626 ( .A1(n_618), .A2(n_581), .A3(n_567), .B(n_569), .Y(n_626) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_604), .A2(n_595), .B(n_591), .C(n_568), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_614), .A2(n_565), .B1(n_578), .B2(n_573), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_611), .B(n_571), .Y(n_629) );
AOI221xp5_ASAP7_75t_SL g630 ( .A1(n_616), .A2(n_544), .B1(n_530), .B2(n_546), .C(n_548), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_608), .B(n_478), .C(n_494), .D(n_489), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_615), .A2(n_548), .B(n_593), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_600), .A2(n_543), .B1(n_592), .B2(n_490), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_601), .B(n_552), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_SL g635 ( .A1(n_626), .A2(n_606), .B(n_483), .C(n_603), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_623), .A2(n_606), .B(n_617), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_622), .A2(n_619), .B(n_613), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_630), .A2(n_625), .B1(n_632), .B2(n_627), .C(n_631), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_624), .B(n_612), .C(n_609), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_628), .A2(n_607), .B1(n_619), .B2(n_621), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_633), .A2(n_551), .B1(n_541), .B2(n_533), .C(n_526), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_640), .B(n_629), .Y(n_642) );
AO22x2_ASAP7_75t_L g643 ( .A1(n_637), .A2(n_634), .B1(n_522), .B2(n_485), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_635), .B(n_455), .C(n_484), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_638), .A2(n_496), .B1(n_497), .B2(n_507), .C(n_531), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_642), .B(n_639), .Y(n_646) );
NOR4xp75_ASAP7_75t_L g647 ( .A(n_645), .B(n_641), .C(n_636), .D(n_499), .Y(n_647) );
NAND3xp33_ASAP7_75t_SL g648 ( .A(n_644), .B(n_455), .C(n_550), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_647), .B(n_550), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_646), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_643), .B1(n_648), .B2(n_545), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_651), .A2(n_649), .B(n_545), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_649), .B1(n_415), .B2(n_432), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_531), .B(n_511), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_654), .B(n_415), .Y(n_655) );
AOI22xp5_ASAP7_75t_SL g656 ( .A1(n_655), .A2(n_511), .B1(n_493), .B2(n_488), .Y(n_656) );
endmodule