module fake_netlist_5_1304_n_747 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_747);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_747;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_509;
wire n_568;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_685;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_32),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_68),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_4),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_54),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_90),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_53),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_55),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_51),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_102),
.Y(n_172)
);

INVxp33_ASAP7_75t_SL g173 ( 
.A(n_94),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_89),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_60),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_112),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_4),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_91),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_47),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_9),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_95),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_25),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_16),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_59),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_70),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_46),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_0),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_21),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_141),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_49),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_23),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_15),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_20),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_33),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_12),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_151),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

AOI22x1_ASAP7_75t_SL g221 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_162),
.B(n_3),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_5),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_5),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_194),
.B(n_6),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_195),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_162),
.B(n_209),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_175),
.B(n_19),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_167),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_157),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_183),
.Y(n_259)
);

AOI21x1_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_188),
.B(n_184),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_185),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_196),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

BUFx6f_ASAP7_75t_SL g269 ( 
.A(n_241),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_198),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_229),
.B(n_199),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_234),
.B(n_161),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_237),
.B(n_166),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_202),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_219),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_237),
.B(n_171),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_222),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_255),
.Y(n_292)
);

BUFx6f_ASAP7_75t_SL g293 ( 
.A(n_213),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_217),
.B(n_172),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_216),
.B(n_174),
.Y(n_296)
);

AND3x2_ASAP7_75t_L g297 ( 
.A(n_215),
.B(n_14),
.C(n_15),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_219),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_231),
.B(n_178),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_215),
.A2(n_170),
.B1(n_204),
.B2(n_210),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_182),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_259),
.B(n_263),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_275),
.B(n_223),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_275),
.B(n_231),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_243),
.B1(n_228),
.B2(n_251),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_246),
.B(n_245),
.C(n_214),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_221),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_275),
.B(n_242),
.Y(n_313)
);

OR2x6_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_225),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_214),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

OAI22x1_ASAP7_75t_L g317 ( 
.A1(n_277),
.A2(n_238),
.B1(n_239),
.B2(n_242),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_279),
.B(n_186),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_279),
.B(n_189),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_220),
.C(n_200),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_261),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_264),
.B(n_268),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_193),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

OR2x6_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_239),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

O2A1O1Ixp5_ASAP7_75t_L g328 ( 
.A1(n_260),
.A2(n_245),
.B(n_218),
.C(n_224),
.Y(n_328)
);

OR2x2_ASAP7_75t_SL g329 ( 
.A(n_297),
.B(n_218),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_227),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_279),
.B(n_201),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_276),
.A2(n_227),
.B1(n_232),
.B2(n_230),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_268),
.B(n_224),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_279),
.B(n_212),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_271),
.B(n_230),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_232),
.B1(n_227),
.B2(n_246),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_257),
.B(n_236),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_257),
.B(n_232),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_283),
.B(n_236),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_22),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_296),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_283),
.B(n_219),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_271),
.B(n_233),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_233),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_283),
.B(n_233),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_274),
.A2(n_233),
.B(n_17),
.C(n_18),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_286),
.B(n_233),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_16),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_278),
.B(n_17),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g352 ( 
.A(n_270),
.B(n_18),
.Y(n_352)
);

OR2x6_ASAP7_75t_L g353 ( 
.A(n_292),
.B(n_24),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_273),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_269),
.B(n_26),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_260),
.B(n_27),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_269),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_272),
.B(n_28),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_273),
.A2(n_280),
.B(n_282),
.C(n_281),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_285),
.B(n_29),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_272),
.B(n_30),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_291),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_280),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_303),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_287),
.B(n_294),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_368),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_262),
.B(n_287),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_305),
.B(n_294),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_312),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_343),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_304),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_337),
.A2(n_323),
.B(n_366),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_284),
.B(n_298),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_323),
.A2(n_262),
.B(n_303),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_324),
.Y(n_382)
);

AOI21x1_ASAP7_75t_L g383 ( 
.A1(n_356),
.A2(n_333),
.B(n_315),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_307),
.A2(n_293),
.B1(n_290),
.B2(n_289),
.Y(n_384)
);

A2O1A1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_350),
.A2(n_290),
.B(n_289),
.C(n_298),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_304),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_308),
.A2(n_293),
.B1(n_290),
.B2(n_289),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_311),
.A2(n_298),
.B(n_284),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_318),
.B(n_293),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_365),
.A2(n_262),
.B(n_303),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_363),
.Y(n_392)
);

AOI22x1_ASAP7_75t_L g393 ( 
.A1(n_317),
.A2(n_298),
.B1(n_284),
.B2(n_304),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_346),
.Y(n_394)
);

BUFx12f_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_L g397 ( 
.A1(n_367),
.A2(n_359),
.B(n_320),
.C(n_313),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_315),
.A2(n_262),
.B(n_303),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_339),
.B(n_31),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_34),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_322),
.B(n_284),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_349),
.Y(n_403)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_309),
.B(n_35),
.C(n_36),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_333),
.A2(n_262),
.B(n_303),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_335),
.A2(n_262),
.B(n_38),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_362),
.B(n_37),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_335),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_345),
.A2(n_39),
.B(n_40),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_336),
.B(n_41),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_345),
.A2(n_42),
.B(n_43),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_326),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_359),
.A2(n_52),
.B(n_56),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_310),
.B(n_57),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_353),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_319),
.B(n_64),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_321),
.B(n_65),
.Y(n_418)
);

AND3x2_ASAP7_75t_L g419 ( 
.A(n_357),
.B(n_66),
.C(n_67),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_325),
.A2(n_69),
.B(n_71),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_340),
.B(n_72),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_341),
.B(n_73),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_342),
.A2(n_74),
.B(n_75),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_76),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_331),
.B(n_77),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_361),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_347),
.A2(n_78),
.B(n_79),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_SL g431 ( 
.A1(n_351),
.A2(n_80),
.B(n_81),
.C(n_84),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_360),
.A2(n_85),
.B(n_86),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_368),
.A2(n_87),
.B(n_92),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_326),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_434)
);

AOI22x1_ASAP7_75t_L g435 ( 
.A1(n_348),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_334),
.B(n_105),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_316),
.B(n_106),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_332),
.A2(n_107),
.B(n_108),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

AO21x2_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_109),
.B(n_110),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_375),
.B(n_314),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_383),
.A2(n_316),
.B(n_114),
.Y(n_443)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_111),
.B(n_115),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_382),
.B(n_314),
.Y(n_445)
);

OA21x2_ASAP7_75t_L g446 ( 
.A1(n_389),
.A2(n_116),
.B(n_117),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_314),
.B(n_120),
.C(n_121),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_439),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_377),
.A2(n_125),
.B(n_126),
.Y(n_450)
);

AO31x2_ASAP7_75t_L g451 ( 
.A1(n_385),
.A2(n_127),
.A3(n_128),
.B(n_129),
.Y(n_451)
);

AO31x2_ASAP7_75t_L g452 ( 
.A1(n_397),
.A2(n_130),
.A3(n_131),
.B(n_132),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_408),
.B(n_134),
.Y(n_453)
);

AO31x2_ASAP7_75t_L g454 ( 
.A1(n_429),
.A2(n_135),
.A3(n_137),
.B(n_138),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_373),
.B(n_139),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_402),
.A2(n_140),
.B(n_142),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_386),
.B(n_143),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_401),
.B(n_147),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_149),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_372),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_371),
.A2(n_153),
.B(n_155),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_374),
.B(n_403),
.Y(n_462)
);

AO21x1_ASAP7_75t_L g463 ( 
.A1(n_417),
.A2(n_427),
.B(n_404),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_376),
.A2(n_409),
.B(n_381),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_411),
.A2(n_393),
.B(n_426),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_381),
.A2(n_409),
.B(n_370),
.Y(n_466)
);

AOI21xp33_ASAP7_75t_L g467 ( 
.A1(n_436),
.A2(n_390),
.B(n_387),
.Y(n_467)
);

AOI21xp33_ASAP7_75t_L g468 ( 
.A1(n_413),
.A2(n_434),
.B(n_416),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_381),
.A2(n_409),
.B1(n_421),
.B2(n_401),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_380),
.A2(n_398),
.B(n_391),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_421),
.A2(n_400),
.B1(n_426),
.B2(n_384),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_400),
.A2(n_425),
.B(n_422),
.C(n_399),
.Y(n_472)
);

AO31x2_ASAP7_75t_L g473 ( 
.A1(n_414),
.A2(n_407),
.A3(n_388),
.B(n_423),
.Y(n_473)
);

AO31x2_ASAP7_75t_L g474 ( 
.A1(n_415),
.A2(n_418),
.A3(n_438),
.B(n_406),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_392),
.B(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_430),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_395),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_433),
.A2(n_420),
.B(n_424),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_419),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_379),
.B(n_410),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_379),
.B(n_412),
.Y(n_482)
);

AOI221xp5_ASAP7_75t_SL g483 ( 
.A1(n_379),
.A2(n_408),
.B1(n_397),
.B2(n_237),
.C(n_373),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_376),
.A2(n_373),
.B(n_377),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_382),
.B(n_375),
.Y(n_485)
);

OAI211xp5_ASAP7_75t_L g486 ( 
.A1(n_374),
.A2(n_300),
.B(n_237),
.C(n_243),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_374),
.B(n_375),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_382),
.B(n_408),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_383),
.A2(n_378),
.B(n_405),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_376),
.A2(n_373),
.B(n_377),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_382),
.B(n_408),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_382),
.B(n_375),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_376),
.A2(n_373),
.B(n_377),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_383),
.A2(n_378),
.B(n_405),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_491),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_468),
.A2(n_469),
.B1(n_471),
.B2(n_441),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

AOI21xp33_ASAP7_75t_SL g498 ( 
.A1(n_487),
.A2(n_492),
.B(n_485),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_459),
.B(n_481),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_459),
.B(n_462),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_460),
.B(n_445),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_463),
.A2(n_450),
.B1(n_449),
.B2(n_458),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_472),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_460),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_478),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_483),
.A2(n_494),
.B(n_489),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_478),
.Y(n_507)
);

CKINVDCx6p67_ASAP7_75t_R g508 ( 
.A(n_480),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_453),
.A2(n_446),
.B1(n_444),
.B2(n_476),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_467),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_484),
.A2(n_493),
.B(n_490),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_447),
.A2(n_466),
.B1(n_455),
.B2(n_464),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_470),
.A2(n_479),
.B(n_443),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_452),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

NOR2x1_ASAP7_75t_SL g516 ( 
.A(n_482),
.B(n_457),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_465),
.Y(n_517)
);

AO31x2_ASAP7_75t_L g518 ( 
.A1(n_477),
.A2(n_452),
.A3(n_451),
.B(n_446),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_452),
.B(n_444),
.Y(n_519)
);

O2A1O1Ixp33_ASAP7_75t_SL g520 ( 
.A1(n_451),
.A2(n_454),
.B(n_440),
.C(n_473),
.Y(n_520)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_461),
.A2(n_456),
.B(n_473),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_451),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_456),
.A2(n_473),
.B1(n_454),
.B2(n_440),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_454),
.B(n_474),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_474),
.A2(n_490),
.B(n_484),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_468),
.A2(n_275),
.B1(n_382),
.B2(n_469),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_441),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_470),
.A2(n_494),
.B(n_489),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_408),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_459),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_470),
.A2(n_494),
.B(n_489),
.Y(n_531)
);

AO21x2_ASAP7_75t_L g532 ( 
.A1(n_465),
.A2(n_450),
.B(n_463),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g533 ( 
.A1(n_465),
.A2(n_450),
.B(n_463),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_459),
.B(n_462),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_465),
.A2(n_450),
.B(n_463),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_441),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_487),
.B(n_374),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_470),
.A2(n_494),
.B(n_489),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_500),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_495),
.B(n_529),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_504),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_497),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_513),
.A2(n_538),
.B(n_531),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_503),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_536),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_495),
.B(n_529),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_528),
.A2(n_521),
.B(n_511),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_527),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_500),
.B(n_534),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_510),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_505),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_514),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_499),
.B(n_526),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_508),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_501),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_515),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_530),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_506),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_507),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_522),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_522),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_498),
.B(n_502),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_525),
.B(n_516),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_496),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_502),
.B(n_517),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_512),
.A2(n_523),
.B(n_509),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_518),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_512),
.B(n_524),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_518),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_532),
.B(n_535),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_519),
.B(n_517),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_544),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_562),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_546),
.B(n_518),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_541),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_546),
.B(n_532),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_558),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_563),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_533),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_533),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_535),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_571),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_573),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_551),
.B(n_509),
.Y(n_591)
);

BUFx2_ASAP7_75t_SL g592 ( 
.A(n_564),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_575),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_540),
.B(n_523),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_568),
.B(n_520),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_561),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_551),
.B(n_563),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_539),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_550),
.B(n_555),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_567),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_553),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_560),
.B(n_556),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_559),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_548),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_542),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_553),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_569),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_549),
.B(n_554),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_549),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_604),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_588),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_588),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_581),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_577),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_576),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_585),
.B(n_574),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_585),
.B(n_574),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_554),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_586),
.B(n_572),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_586),
.B(n_559),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_583),
.B(n_566),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_579),
.B(n_552),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_590),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_596),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_580),
.B(n_570),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_583),
.B(n_566),
.Y(n_627)
);

INVxp67_ASAP7_75t_SL g628 ( 
.A(n_589),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_597),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_596),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_580),
.B(n_570),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_582),
.Y(n_632)
);

AND2x4_ASAP7_75t_SL g633 ( 
.A(n_582),
.B(n_551),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_601),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_602),
.B(n_566),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_578),
.B(n_547),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_603),
.A2(n_552),
.B1(n_557),
.B2(n_543),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_608),
.B(n_557),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_620),
.B(n_578),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_625),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_634),
.B(n_607),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_633),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_625),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_630),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_603),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_628),
.A2(n_591),
.B(n_594),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_630),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

BUFx2_ASAP7_75t_SL g650 ( 
.A(n_613),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_612),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_612),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_610),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_614),
.B(n_594),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_635),
.B(n_593),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_617),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_633),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_624),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_624),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_632),
.B(n_593),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_615),
.Y(n_662)
);

CKINVDCx14_ASAP7_75t_R g663 ( 
.A(n_629),
.Y(n_663)
);

AOI322xp5_ASAP7_75t_L g664 ( 
.A1(n_654),
.A2(n_637),
.A3(n_621),
.B1(n_618),
.B2(n_616),
.C1(n_626),
.C2(n_631),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_SL g665 ( 
.A1(n_645),
.A2(n_619),
.B1(n_638),
.B2(n_623),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_655),
.B(n_631),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_650),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_639),
.B(n_626),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_641),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_653),
.B(n_634),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_652),
.B(n_636),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_619),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_652),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_656),
.B(n_636),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_656),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_657),
.B(n_618),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_657),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_662),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_640),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_643),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_647),
.B(n_616),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_662),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_648),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_665),
.A2(n_646),
.B(n_661),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_680),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_669),
.B(n_646),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_681),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_684),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_673),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_667),
.A2(n_627),
.B1(n_622),
.B2(n_635),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_675),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_672),
.A2(n_601),
.B1(n_600),
.B2(n_629),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_678),
.Y(n_694)
);

AOI31xp33_ASAP7_75t_SL g695 ( 
.A1(n_679),
.A2(n_600),
.A3(n_595),
.B(n_663),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_666),
.B(n_663),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_683),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_683),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_685),
.B(n_687),
.C(n_664),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_690),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_692),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_691),
.A2(n_622),
.B1(n_627),
.B2(n_621),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_686),
.B(n_668),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_696),
.B(n_666),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_699),
.B(n_688),
.Y(n_705)
);

AOI222xp33_ASAP7_75t_L g706 ( 
.A1(n_700),
.A2(n_693),
.B1(n_689),
.B2(n_698),
.C1(n_668),
.C2(n_682),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_L g707 ( 
.A1(n_701),
.A2(n_693),
.B1(n_698),
.B2(n_682),
.C(n_697),
.Y(n_707)
);

AOI32xp33_ASAP7_75t_L g708 ( 
.A1(n_704),
.A2(n_671),
.A3(n_674),
.B1(n_695),
.B2(n_694),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_703),
.B(n_671),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_702),
.B(n_670),
.C(n_697),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_709),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_598),
.C(n_605),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_706),
.B(n_674),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_710),
.Y(n_714)
);

NOR4xp75_ASAP7_75t_L g715 ( 
.A(n_713),
.B(n_708),
.C(n_707),
.D(n_678),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_SL g716 ( 
.A(n_714),
.B(n_712),
.C(n_711),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_714),
.B(n_629),
.C(n_606),
.Y(n_717)
);

AND3x4_ASAP7_75t_L g718 ( 
.A(n_715),
.B(n_716),
.C(n_717),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_717),
.B(n_678),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_642),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_716),
.B(n_598),
.C(n_605),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_720),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_721),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_718),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_719),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_720),
.B(n_642),
.Y(n_726)
);

XNOR2xp5_ASAP7_75t_L g727 ( 
.A(n_718),
.B(n_609),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_722),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_724),
.A2(n_726),
.B(n_727),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_723),
.B(n_677),
.Y(n_730)
);

NAND4xp75_ASAP7_75t_L g731 ( 
.A(n_725),
.B(n_606),
.C(n_659),
.D(n_660),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_722),
.B(n_676),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_728),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_SL g734 ( 
.A1(n_730),
.A2(n_658),
.B1(n_592),
.B2(n_582),
.Y(n_734)
);

XNOR2xp5_ASAP7_75t_L g735 ( 
.A(n_729),
.B(n_609),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_732),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_733),
.A2(n_731),
.B1(n_658),
.B2(n_661),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_736),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_735),
.B(n_651),
.Y(n_739)
);

OAI21x1_ASAP7_75t_SL g740 ( 
.A1(n_738),
.A2(n_734),
.B(n_587),
.Y(n_740)
);

OAI21xp33_ASAP7_75t_L g741 ( 
.A1(n_739),
.A2(n_609),
.B(n_632),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_737),
.A2(n_589),
.B(n_587),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_740),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_742),
.A2(n_584),
.B(n_649),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_743),
.A2(n_741),
.B(n_744),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_582),
.B1(n_592),
.B2(n_597),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_746),
.A2(n_582),
.B1(n_597),
.B2(n_629),
.Y(n_747)
);


endmodule