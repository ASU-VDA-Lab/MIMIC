module real_aes_17141_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_1580, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_1580;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_1404;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_0), .A2(n_73), .B1(n_541), .B2(n_560), .Y(n_559) );
INVxp33_ASAP7_75t_SL g665 ( .A(n_0), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_1), .Y(n_864) );
XOR2xp5_ASAP7_75t_L g897 ( .A(n_2), .B(n_898), .Y(n_897) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_3), .A2(n_94), .B1(n_1093), .B2(n_1096), .Y(n_1292) );
INVxp67_ASAP7_75t_SL g1307 ( .A(n_3), .Y(n_1307) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_4), .Y(n_1033) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_5), .A2(n_87), .B1(n_834), .B2(n_836), .C(n_837), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_5), .A2(n_145), .B1(n_548), .B2(n_724), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g1338 ( .A(n_6), .Y(n_1338) );
INVx1_ASAP7_75t_L g1181 ( .A(n_7), .Y(n_1181) );
INVx1_ASAP7_75t_L g1143 ( .A(n_8), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g1163 ( .A1(n_8), .A2(n_156), .B1(n_1156), .B2(n_1159), .C(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_9), .A2(n_44), .B1(n_909), .B2(n_911), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_9), .A2(n_225), .B1(n_639), .B2(n_937), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_10), .A2(n_220), .B1(n_602), .B2(n_1004), .C(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1250 ( .A(n_10), .Y(n_1250) );
INVx1_ASAP7_75t_L g1275 ( .A(n_11), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1397 ( .A1(n_12), .A2(n_229), .B1(n_909), .B2(n_911), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_12), .A2(n_196), .B1(n_779), .B2(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1226 ( .A(n_13), .Y(n_1226) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_13), .A2(n_163), .B1(n_926), .B2(n_1254), .C(n_1255), .Y(n_1253) );
AOI21xp33_ASAP7_75t_L g1194 ( .A1(n_14), .A2(n_555), .B(n_738), .Y(n_1194) );
INVx1_ASAP7_75t_L g1214 ( .A(n_14), .Y(n_1214) );
INVx1_ASAP7_75t_L g509 ( .A(n_15), .Y(n_509) );
AND2x2_ASAP7_75t_L g621 ( .A(n_15), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g634 ( .A(n_15), .B(n_239), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_15), .B(n_519), .Y(n_693) );
AND2x2_ASAP7_75t_L g291 ( .A(n_16), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g294 ( .A(n_16), .B(n_112), .Y(n_294) );
INVx2_ASAP7_75t_L g298 ( .A(n_16), .Y(n_298) );
INVx1_ASAP7_75t_L g1392 ( .A(n_17), .Y(n_1392) );
OAI221xp5_ASAP7_75t_L g1419 ( .A1(n_17), .A2(n_175), .B1(n_1420), .B2(n_1421), .C(n_1422), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_18), .A2(n_242), .B1(n_743), .B2(n_1013), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g1167 ( .A(n_18), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1288 ( .A1(n_19), .A2(n_724), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1320 ( .A(n_19), .Y(n_1320) );
INVx1_ASAP7_75t_L g1337 ( .A(n_20), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1466 ( .A1(n_21), .A2(n_141), .B1(n_1467), .B2(n_1469), .Y(n_1466) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_21), .A2(n_141), .B1(n_511), .B2(n_1500), .Y(n_1499) );
OAI222xp33_ASAP7_75t_L g808 ( .A1(n_22), .A2(n_161), .B1(n_809), .B2(n_813), .C1(n_818), .C2(n_825), .Y(n_808) );
INVx1_ASAP7_75t_L g871 ( .A(n_22), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_23), .A2(n_164), .B1(n_884), .B2(n_885), .Y(n_1299) );
AOI32xp33_ASAP7_75t_L g1309 ( .A1(n_23), .A2(n_934), .A3(n_1310), .B1(n_1312), .B2(n_1580), .Y(n_1309) );
XNOR2x2_ASAP7_75t_L g1219 ( .A(n_24), .B(n_1220), .Y(n_1219) );
OAI21xp5_ASAP7_75t_L g942 ( .A1(n_25), .A2(n_943), .B(n_944), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_26), .A2(n_187), .B1(n_293), .B2(n_299), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_27), .A2(n_199), .B1(n_299), .B2(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g1189 ( .A(n_28), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_28), .A2(n_158), .B1(n_689), .B2(n_790), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_29), .B(n_1291), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1325 ( .A1(n_29), .A2(n_164), .B1(n_1054), .B2(n_1326), .C(n_1327), .Y(n_1325) );
INVx1_ASAP7_75t_L g1091 ( .A(n_30), .Y(n_1091) );
INVx1_ASAP7_75t_L g940 ( .A(n_31), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_32), .A2(n_79), .B1(n_563), .B2(n_564), .C(n_566), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_32), .A2(n_35), .B1(n_688), .B2(n_689), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_33), .Y(n_750) );
INVx1_ASAP7_75t_L g919 ( .A(n_34), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_35), .A2(n_143), .B1(n_532), .B2(n_541), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_36), .A2(n_214), .B1(n_288), .B2(n_296), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_37), .A2(n_186), .B1(n_534), .B2(n_1291), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_37), .A2(n_150), .B1(n_1367), .B2(n_1370), .Y(n_1369) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_38), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_39), .B(n_1286), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_39), .A2(n_276), .B1(n_1254), .B2(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g845 ( .A(n_40), .Y(n_845) );
INVx1_ASAP7_75t_L g580 ( .A(n_41), .Y(n_580) );
OA222x2_ASAP7_75t_L g627 ( .A1(n_41), .A2(n_182), .B1(n_275), .B2(n_628), .C1(n_635), .C2(n_643), .Y(n_627) );
INVx1_ASAP7_75t_L g1227 ( .A(n_42), .Y(n_1227) );
AOI221xp5_ASAP7_75t_L g1246 ( .A1(n_42), .A2(n_77), .B1(n_834), .B2(n_1247), .C(n_1249), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_43), .A2(n_219), .B1(n_548), .B2(n_550), .C(n_555), .Y(n_547) );
INVx1_ASAP7_75t_L g682 ( .A(n_43), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_44), .A2(n_132), .B1(n_926), .B2(n_927), .C(n_928), .Y(n_925) );
INVx1_ASAP7_75t_L g1343 ( .A(n_45), .Y(n_1343) );
INVx1_ASAP7_75t_L g1442 ( .A(n_46), .Y(n_1442) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_47), .A2(n_222), .B1(n_288), .B2(n_299), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_48), .A2(n_117), .B1(n_288), .B2(n_296), .Y(n_332) );
INVxp67_ASAP7_75t_SL g819 ( .A(n_49), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_49), .A2(n_87), .B1(n_548), .B2(n_724), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_50), .A2(n_106), .B1(n_288), .B2(n_296), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g1236 ( .A1(n_51), .A2(n_70), .B1(n_582), .B2(n_998), .C(n_999), .Y(n_1236) );
INVxp67_ASAP7_75t_SL g1242 ( .A(n_51), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1042 ( .A1(n_52), .A2(n_184), .B1(n_998), .B2(n_999), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_52), .A2(n_83), .B1(n_977), .B2(n_979), .Y(n_1059) );
OAI211xp5_ASAP7_75t_SL g1177 ( .A1(n_53), .A2(n_1178), .B(n_1179), .C(n_1182), .Y(n_1177) );
INVx1_ASAP7_75t_L g1200 ( .A(n_53), .Y(n_1200) );
INVx1_ASAP7_75t_L g816 ( .A(n_54), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_54), .A2(n_249), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g913 ( .A1(n_55), .A2(n_118), .B1(n_534), .B2(n_605), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_55), .A2(n_82), .B1(n_656), .B2(n_934), .C(n_935), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_56), .A2(n_124), .B1(n_1134), .B2(n_1135), .C(n_1136), .Y(n_1133) );
INVx1_ASAP7_75t_L g1161 ( .A(n_56), .Y(n_1161) );
INVx1_ASAP7_75t_L g540 ( .A(n_57), .Y(n_540) );
INVx1_ASAP7_75t_L g546 ( .A(n_57), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_58), .Y(n_959) );
CKINVDCx5p33_ASAP7_75t_R g973 ( .A(n_59), .Y(n_973) );
INVx1_ASAP7_75t_L g1082 ( .A(n_60), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_61), .A2(n_104), .B1(n_911), .B2(n_1141), .C(n_1142), .Y(n_1140) );
INVx1_ASAP7_75t_L g1166 ( .A(n_61), .Y(n_1166) );
INVx1_ASAP7_75t_L g290 ( .A(n_62), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_63), .A2(n_228), .B1(n_743), .B2(n_1013), .Y(n_1235) );
INVx1_ASAP7_75t_L g1245 ( .A(n_63), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_64), .A2(n_88), .B1(n_296), .B2(n_303), .Y(n_317) );
INVx2_ASAP7_75t_L g558 ( .A(n_65), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_66), .A2(n_249), .B1(n_639), .B2(n_839), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_66), .A2(n_167), .B1(n_885), .B2(n_887), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_67), .A2(n_231), .B1(n_550), .B2(n_1004), .Y(n_1545) );
AOI221xp5_ASAP7_75t_L g1561 ( .A1(n_67), .A2(n_179), .B1(n_1372), .B2(n_1375), .C(n_1562), .Y(n_1561) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_68), .A2(n_201), .B1(n_1093), .B2(n_1096), .Y(n_1223) );
INVx1_ASAP7_75t_L g1243 ( .A(n_68), .Y(n_1243) );
INVx1_ASAP7_75t_L g1031 ( .A(n_69), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_69), .A2(n_237), .B1(n_639), .B2(n_688), .Y(n_1053) );
INVx1_ASAP7_75t_L g1263 ( .A(n_70), .Y(n_1263) );
CKINVDCx5p33_ASAP7_75t_R g1041 ( .A(n_71), .Y(n_1041) );
AOI21xp33_ASAP7_75t_L g1086 ( .A1(n_72), .A2(n_552), .B(n_555), .Y(n_1086) );
INVxp67_ASAP7_75t_L g1111 ( .A(n_72), .Y(n_1111) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_73), .Y(n_686) );
INVx1_ASAP7_75t_L g985 ( .A(n_74), .Y(n_985) );
AOI22xp33_ASAP7_75t_SL g1548 ( .A1(n_75), .A2(n_125), .B1(n_853), .B2(n_1544), .Y(n_1548) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_75), .A2(n_153), .B1(n_1326), .B2(n_1327), .Y(n_1563) );
INVx1_ASAP7_75t_L g1144 ( .A(n_76), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g1228 ( .A1(n_77), .A2(n_221), .B1(n_1004), .B2(n_1229), .C(n_1230), .Y(n_1228) );
OAI211xp5_ASAP7_75t_L g1472 ( .A1(n_78), .A2(n_1473), .B(n_1475), .C(n_1477), .Y(n_1472) );
INVx1_ASAP7_75t_L g1514 ( .A(n_78), .Y(n_1514) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_79), .A2(n_219), .B1(n_656), .B2(n_658), .C(n_661), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_80), .A2(n_140), .B1(n_288), .B2(n_296), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_81), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_82), .A2(n_238), .B1(n_905), .B2(n_906), .Y(n_904) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_83), .A2(n_183), .B1(n_732), .B2(n_1039), .C(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1454 ( .A(n_84), .Y(n_1454) );
INVx1_ASAP7_75t_L g601 ( .A(n_85), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_85), .B(n_614), .Y(n_613) );
OAI222xp33_ASAP7_75t_L g993 ( .A1(n_86), .A2(n_138), .B1(n_250), .B2(n_745), .C1(n_994), .C2(n_995), .Y(n_993) );
INVx1_ASAP7_75t_L g1016 ( .A(n_86), .Y(n_1016) );
INVx1_ASAP7_75t_L g1197 ( .A(n_89), .Y(n_1197) );
XOR2x1_ASAP7_75t_L g1270 ( .A(n_90), .B(n_1271), .Y(n_1270) );
AOI22xp33_ASAP7_75t_SL g1346 ( .A1(n_91), .A2(n_99), .B1(n_906), .B2(n_1347), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1364 ( .A1(n_91), .A2(n_137), .B1(n_934), .B2(n_935), .C(n_1324), .Y(n_1364) );
CKINVDCx5p33_ASAP7_75t_R g1553 ( .A(n_92), .Y(n_1553) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_93), .A2(n_147), .B1(n_566), .B2(n_1002), .C(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_93), .A2(n_210), .B1(n_782), .B2(n_790), .Y(n_1215) );
INVx1_ASAP7_75t_L g1272 ( .A(n_94), .Y(n_1272) );
CKINVDCx5p33_ASAP7_75t_R g1539 ( .A(n_95), .Y(n_1539) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_96), .A2(n_195), .B1(n_1093), .B2(n_1096), .Y(n_1092) );
INVxp67_ASAP7_75t_SL g1099 ( .A(n_96), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_97), .A2(n_139), .B1(n_288), .B2(n_296), .Y(n_321) );
INVx1_ASAP7_75t_L g1439 ( .A(n_98), .Y(n_1439) );
AOI221xp5_ASAP7_75t_L g1371 ( .A1(n_99), .A2(n_224), .B1(n_1372), .B2(n_1373), .C(n_1375), .Y(n_1371) );
INVx1_ASAP7_75t_L g604 ( .A(n_100), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_100), .A2(n_198), .B1(n_699), .B2(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g972 ( .A(n_101), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_101), .A2(n_162), .B1(n_1002), .B2(n_1004), .C(n_1005), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_102), .A2(n_130), .B1(n_605), .B2(n_724), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1409 ( .A1(n_102), .A2(n_280), .B1(n_658), .B2(n_1410), .C(n_1413), .Y(n_1409) );
AOI22xp5_ASAP7_75t_SL g320 ( .A1(n_103), .A2(n_269), .B1(n_299), .B2(n_303), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g1155 ( .A1(n_104), .A2(n_205), .B1(n_1156), .B2(n_1159), .C(n_1160), .Y(n_1155) );
AND2x2_ASAP7_75t_L g289 ( .A(n_105), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_105), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_107), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_108), .A2(n_176), .B1(n_564), .B2(n_740), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_108), .A2(n_109), .B1(n_689), .B2(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g762 ( .A(n_109), .Y(n_762) );
OAI21xp5_ASAP7_75t_SL g1378 ( .A1(n_110), .A2(n_943), .B(n_1379), .Y(n_1378) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_111), .A2(n_121), .B1(n_293), .B2(n_299), .Y(n_331) );
INVx1_ASAP7_75t_L g292 ( .A(n_112), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_112), .B(n_298), .Y(n_300) );
XOR2x2_ASAP7_75t_L g1383 ( .A(n_113), .B(n_1384), .Y(n_1383) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_114), .A2(n_276), .B1(n_1294), .B2(n_1297), .C(n_1298), .Y(n_1293) );
INVx1_ASAP7_75t_L g1321 ( .A(n_114), .Y(n_1321) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_115), .A2(n_710), .B1(n_711), .B2(n_801), .Y(n_709) );
INVx1_ASAP7_75t_L g801 ( .A(n_115), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_116), .A2(n_274), .B1(n_288), .B2(n_293), .Y(n_287) );
XNOR2xp5_ASAP7_75t_L g1334 ( .A(n_116), .B(n_1335), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_118), .A2(n_238), .B1(n_689), .B2(n_839), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g1139 ( .A1(n_119), .A2(n_171), .B1(n_1093), .B2(n_1096), .Y(n_1139) );
INVxp67_ASAP7_75t_SL g1169 ( .A(n_119), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_120), .A2(n_270), .B1(n_743), .B2(n_1013), .Y(n_1277) );
INVxp33_ASAP7_75t_L g1329 ( .A(n_120), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g1535 ( .A(n_122), .Y(n_1535) );
AOI22xp33_ASAP7_75t_SL g1541 ( .A1(n_123), .A2(n_153), .B1(n_1542), .B2(n_1544), .Y(n_1541) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_123), .A2(n_125), .B1(n_935), .B2(n_1324), .C(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1165 ( .A(n_124), .Y(n_1165) );
INVx2_ASAP7_75t_L g557 ( .A(n_126), .Y(n_557) );
INVx1_ASAP7_75t_L g569 ( .A(n_126), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_126), .B(n_558), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_127), .Y(n_1026) );
INVx1_ASAP7_75t_L g988 ( .A(n_128), .Y(n_988) );
OAI22xp33_ASAP7_75t_L g997 ( .A1(n_128), .A2(n_173), .B1(n_998), .B2(n_999), .Y(n_997) );
INVx1_ASAP7_75t_L g1084 ( .A(n_129), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_130), .A2(n_272), .B1(n_839), .B2(n_1415), .Y(n_1425) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_131), .A2(n_245), .B1(n_288), .B2(n_296), .Y(n_304) );
XOR2xp5_ASAP7_75t_L g1431 ( .A(n_131), .B(n_1432), .Y(n_1431) );
CKINVDCx5p33_ASAP7_75t_R g1578 ( .A(n_131), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_132), .A2(n_225), .B1(n_909), .B2(n_911), .Y(n_908) );
INVxp67_ASAP7_75t_SL g1193 ( .A(n_133), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_133), .A2(n_147), .B1(n_1205), .B2(n_1207), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_134), .A2(n_165), .B1(n_715), .B2(n_848), .Y(n_1387) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_135), .A2(n_169), .B1(n_582), .B2(n_998), .C(n_999), .Y(n_1276) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_135), .B(n_987), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_136), .A2(n_196), .B1(n_909), .B2(n_1396), .Y(n_1395) );
AOI21xp33_ASAP7_75t_L g1424 ( .A1(n_136), .A2(n_928), .B(n_1410), .Y(n_1424) );
AOI221xp5_ASAP7_75t_L g1352 ( .A1(n_137), .A2(n_150), .B1(n_602), .B2(n_906), .C(n_1353), .Y(n_1352) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_138), .A2(n_173), .B1(n_694), .B2(n_977), .C(n_979), .Y(n_976) );
INVx1_ASAP7_75t_L g947 ( .A(n_139), .Y(n_947) );
OAI221xp5_ASAP7_75t_L g1130 ( .A1(n_142), .A2(n_208), .B1(n_582), .B2(n_998), .C(n_999), .Y(n_1130) );
OAI21xp33_ASAP7_75t_L g1151 ( .A1(n_142), .A2(n_643), .B(n_694), .Y(n_1151) );
INVxp67_ASAP7_75t_SL g662 ( .A(n_143), .Y(n_662) );
INVx1_ASAP7_75t_L g1448 ( .A(n_144), .Y(n_1448) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_145), .Y(n_822) );
INVx1_ASAP7_75t_L g1234 ( .A(n_146), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_148), .A2(n_1175), .B1(n_1217), .B2(n_1218), .Y(n_1174) );
INVx1_ASAP7_75t_L g1218 ( .A(n_148), .Y(n_1218) );
OAI211xp5_ASAP7_75t_SL g829 ( .A1(n_149), .A2(n_830), .B(n_832), .C(n_841), .Y(n_829) );
INVx1_ASAP7_75t_L g876 ( .A(n_149), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_151), .Y(n_1386) );
XOR2x2_ASAP7_75t_L g1065 ( .A(n_152), .B(n_1066), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g311 ( .A1(n_154), .A2(n_260), .B1(n_299), .B2(n_312), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_155), .A2(n_1013), .B1(n_1029), .B2(n_1032), .Y(n_1028) );
INVx1_ASAP7_75t_L g1048 ( .A(n_155), .Y(n_1048) );
INVx1_ASAP7_75t_L g1137 ( .A(n_156), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_157), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g1195 ( .A1(n_158), .A2(n_210), .B1(n_564), .B2(n_885), .Y(n_1195) );
INVx1_ASAP7_75t_L g1183 ( .A(n_159), .Y(n_1183) );
OAI221xp5_ASAP7_75t_L g1202 ( .A1(n_159), .A2(n_207), .B1(n_979), .B2(n_1153), .C(n_1203), .Y(n_1202) );
CKINVDCx5p33_ASAP7_75t_R g1552 ( .A(n_160), .Y(n_1552) );
INVx1_ASAP7_75t_L g867 ( .A(n_161), .Y(n_867) );
INVx1_ASAP7_75t_L g954 ( .A(n_162), .Y(n_954) );
INVx1_ASAP7_75t_L g1231 ( .A(n_163), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1406 ( .A1(n_165), .A2(n_1407), .B(n_1408), .C(n_1416), .Y(n_1406) );
BUFx3_ASAP7_75t_L g537 ( .A(n_166), .Y(n_537) );
INVx1_ASAP7_75t_L g815 ( .A(n_167), .Y(n_815) );
INVx1_ASAP7_75t_L g1184 ( .A(n_168), .Y(n_1184) );
INVxp67_ASAP7_75t_SL g1306 ( .A(n_169), .Y(n_1306) );
INVx1_ASAP7_75t_L g1129 ( .A(n_170), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_171), .A2(n_208), .B1(n_979), .B2(n_1153), .Y(n_1152) );
XNOR2x1_ASAP7_75t_L g804 ( .A(n_172), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g1069 ( .A(n_174), .Y(n_1069) );
INVx1_ASAP7_75t_L g1391 ( .A(n_175), .Y(n_1391) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_176), .A2(n_247), .B1(n_779), .B2(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g1486 ( .A(n_177), .Y(n_1486) );
OAI211xp5_ASAP7_75t_L g1503 ( .A1(n_177), .A2(n_1504), .B(n_1507), .C(n_1510), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_178), .A2(n_179), .B1(n_738), .B2(n_1291), .Y(n_1546) );
AOI22xp33_ASAP7_75t_SL g1559 ( .A1(n_178), .A2(n_231), .B1(n_1326), .B2(n_1327), .Y(n_1559) );
OAI21xp5_ASAP7_75t_SL g1564 ( .A1(n_180), .A2(n_943), .B(n_1565), .Y(n_1564) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_181), .Y(n_516) );
INVx1_ASAP7_75t_L g606 ( .A(n_182), .Y(n_606) );
OAI211xp5_ASAP7_75t_L g1045 ( .A1(n_183), .A2(n_1046), .B(n_1047), .C(n_1050), .Y(n_1045) );
INVx1_ASAP7_75t_L g1049 ( .A(n_184), .Y(n_1049) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_185), .Y(n_1025) );
AOI22xp33_ASAP7_75t_SL g1365 ( .A1(n_186), .A2(n_271), .B1(n_1366), .B2(n_1367), .Y(n_1365) );
INVx1_ASAP7_75t_L g939 ( .A(n_188), .Y(n_939) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_189), .A2(n_848), .B(n_851), .Y(n_847) );
INVx1_ASAP7_75t_L g917 ( .A(n_190), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g1076 ( .A1(n_191), .A2(n_566), .B(n_724), .Y(n_1076) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_191), .Y(n_1108) );
INVx1_ASAP7_75t_L g728 ( .A(n_192), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g783 ( .A1(n_192), .A2(n_643), .B1(n_784), .B2(n_792), .C(n_793), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g966 ( .A(n_193), .Y(n_966) );
INVx1_ASAP7_75t_L g1035 ( .A(n_194), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_194), .A2(n_204), .B1(n_688), .B2(n_782), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1121 ( .A1(n_195), .A2(n_223), .B1(n_694), .B2(n_977), .C(n_979), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_197), .A2(n_257), .B1(n_1400), .B2(n_1404), .Y(n_1399) );
INVx1_ASAP7_75t_L g1417 ( .A(n_197), .Y(n_1417) );
INVx1_ASAP7_75t_L g577 ( .A(n_198), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_200), .A2(n_203), .B1(n_293), .B2(n_299), .Y(n_342) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_201), .Y(n_1261) );
INVx1_ASAP7_75t_L g1090 ( .A(n_202), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_204), .A2(n_237), .B1(n_565), .B2(n_885), .C(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1138 ( .A(n_205), .Y(n_1138) );
INVx1_ASAP7_75t_L g1452 ( .A(n_206), .Y(n_1452) );
INVx1_ASAP7_75t_L g1198 ( .A(n_207), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_209), .Y(n_718) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_211), .Y(n_515) );
INVx1_ASAP7_75t_L g1079 ( .A(n_212), .Y(n_1079) );
INVx1_ASAP7_75t_L g1446 ( .A(n_213), .Y(n_1446) );
XNOR2x1_ASAP7_75t_L g1125 ( .A(n_214), .B(n_1126), .Y(n_1125) );
CKINVDCx5p33_ASAP7_75t_R g1538 ( .A(n_215), .Y(n_1538) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_216), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g962 ( .A(n_217), .Y(n_962) );
INVxp67_ASAP7_75t_SL g984 ( .A(n_218), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_218), .A2(n_1009), .B1(n_1011), .B2(n_1013), .Y(n_1008) );
INVx1_ASAP7_75t_L g1256 ( .A(n_220), .Y(n_1256) );
INVx1_ASAP7_75t_L g1259 ( .A(n_221), .Y(n_1259) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_223), .A2(n_244), .B1(n_582), .B2(n_998), .C(n_999), .Y(n_1070) );
AOI22xp33_ASAP7_75t_SL g1355 ( .A1(n_224), .A2(n_271), .B1(n_1135), .B2(n_1347), .Y(n_1355) );
INVx1_ASAP7_75t_L g1281 ( .A(n_226), .Y(n_1281) );
AOI22xp5_ASAP7_75t_L g1528 ( .A1(n_227), .A2(n_1529), .B1(n_1530), .B2(n_1531), .Y(n_1528) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_227), .Y(n_1529) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_228), .Y(n_1238) );
INVx1_ASAP7_75t_L g1423 ( .A(n_229), .Y(n_1423) );
INVx1_ASAP7_75t_L g1444 ( .A(n_230), .Y(n_1444) );
INVx1_ASAP7_75t_L g1359 ( .A(n_232), .Y(n_1359) );
INVx1_ASAP7_75t_L g1341 ( .A(n_233), .Y(n_1341) );
INVx1_ASAP7_75t_L g713 ( .A(n_234), .Y(n_713) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_235), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_235), .A2(n_582), .B1(n_743), .B2(n_746), .C(n_756), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_236), .Y(n_956) );
BUFx3_ASAP7_75t_L g519 ( .A(n_239), .Y(n_519) );
INVx1_ASAP7_75t_L g622 ( .A(n_239), .Y(n_622) );
INVx1_ASAP7_75t_L g707 ( .A(n_240), .Y(n_707) );
OAI22xp33_ASAP7_75t_L g1487 ( .A1(n_241), .A2(n_267), .B1(n_1488), .B2(n_1490), .Y(n_1487) );
OAI22xp5_ASAP7_75t_L g1515 ( .A1(n_241), .A2(n_267), .B1(n_1516), .B2(n_1518), .Y(n_1515) );
INVxp67_ASAP7_75t_SL g1146 ( .A(n_242), .Y(n_1146) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_243), .A2(n_555), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g776 ( .A(n_243), .Y(n_776) );
INVxp67_ASAP7_75t_SL g1123 ( .A(n_244), .Y(n_1123) );
INVx1_ASAP7_75t_L g1180 ( .A(n_246), .Y(n_1180) );
INVx1_ASAP7_75t_L g755 ( .A(n_247), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_248), .Y(n_725) );
INVx1_ASAP7_75t_L g990 ( .A(n_250), .Y(n_990) );
INVx2_ASAP7_75t_L g612 ( .A(n_251), .Y(n_612) );
INVx1_ASAP7_75t_L g619 ( .A(n_251), .Y(n_619) );
INVx1_ASAP7_75t_L g632 ( .A(n_251), .Y(n_632) );
INVx1_ASAP7_75t_L g1482 ( .A(n_252), .Y(n_1482) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_253), .A2(n_265), .B1(n_542), .B2(n_565), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1119 ( .A(n_253), .Y(n_1119) );
INVx1_ASAP7_75t_L g900 ( .A(n_254), .Y(n_900) );
INVx1_ASAP7_75t_L g1232 ( .A(n_255), .Y(n_1232) );
INVx1_ASAP7_75t_L g1361 ( .A(n_256), .Y(n_1361) );
INVx1_ASAP7_75t_L g1418 ( .A(n_257), .Y(n_1418) );
INVx1_ASAP7_75t_L g1019 ( .A(n_258), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_259), .A2(n_262), .B1(n_296), .B2(n_299), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_261), .Y(n_730) );
INVx1_ASAP7_75t_L g1037 ( .A(n_263), .Y(n_1037) );
INVx1_ASAP7_75t_L g1073 ( .A(n_264), .Y(n_1073) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_265), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_266), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g1187 ( .A(n_268), .Y(n_1187) );
INVxp67_ASAP7_75t_SL g1301 ( .A(n_270), .Y(n_1301) );
AOI22xp33_ASAP7_75t_SL g1398 ( .A1(n_272), .A2(n_280), .B1(n_605), .B2(n_724), .Y(n_1398) );
INVx1_ASAP7_75t_L g1438 ( .A(n_273), .Y(n_1438) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_275), .A2(n_279), .B1(n_594), .B2(n_595), .C(n_600), .Y(n_593) );
INVx1_ASAP7_75t_L g727 ( .A(n_277), .Y(n_727) );
INVx1_ASAP7_75t_L g843 ( .A(n_278), .Y(n_843) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_279), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_296), .B1(n_497), .B2(n_520), .C(n_1429), .Y(n_281) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_388), .B(n_409), .Y(n_283) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_305), .B(n_336), .C(n_374), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_301), .Y(n_285) );
INVx3_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
INVx3_ASAP7_75t_L g385 ( .A(n_286), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_286), .B(n_362), .Y(n_387) );
AND2x2_ASAP7_75t_L g407 ( .A(n_286), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g445 ( .A(n_286), .B(n_430), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_286), .B(n_301), .Y(n_449) );
AND2x2_ASAP7_75t_L g454 ( .A(n_286), .B(n_354), .Y(n_454) );
AND2x4_ASAP7_75t_SL g286 ( .A(n_287), .B(n_295), .Y(n_286) );
AND2x6_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
AND2x2_ASAP7_75t_L g293 ( .A(n_289), .B(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g296 ( .A(n_289), .B(n_297), .Y(n_296) );
AND2x6_ASAP7_75t_L g299 ( .A(n_289), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g303 ( .A(n_289), .B(n_294), .Y(n_303) );
AND2x2_ASAP7_75t_L g312 ( .A(n_289), .B(n_294), .Y(n_312) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_290), .Y(n_502) );
AND2x2_ASAP7_75t_L g297 ( .A(n_292), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g1575 ( .A(n_297), .Y(n_1575) );
AND2x2_ASAP7_75t_L g354 ( .A(n_301), .B(n_330), .Y(n_354) );
AND2x2_ASAP7_75t_L g384 ( .A(n_301), .B(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g393 ( .A(n_301), .B(n_329), .Y(n_393) );
OR2x2_ASAP7_75t_L g401 ( .A(n_301), .B(n_330), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_301), .B(n_416), .Y(n_424) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
AND2x4_ASAP7_75t_L g349 ( .A(n_302), .B(n_304), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_314), .B(n_322), .C(n_327), .Y(n_305) );
AND2x2_ASAP7_75t_L g365 ( .A(n_306), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_306), .B(n_361), .Y(n_431) );
AND2x2_ASAP7_75t_L g487 ( .A(n_306), .B(n_326), .Y(n_487) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .Y(n_306) );
INVx3_ASAP7_75t_L g325 ( .A(n_307), .Y(n_325) );
INVx2_ASAP7_75t_L g358 ( .A(n_307), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_307), .B(n_310), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_307), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g457 ( .A(n_307), .B(n_329), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_307), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_310), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_310), .B(n_335), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_310), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_310), .B(n_369), .Y(n_403) );
OR2x2_ASAP7_75t_L g466 ( .A(n_310), .B(n_376), .Y(n_466) );
AND2x2_ASAP7_75t_L g494 ( .A(n_310), .B(n_366), .Y(n_494) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x2_ASAP7_75t_L g338 ( .A(n_311), .B(n_313), .Y(n_338) );
INVx1_ASAP7_75t_L g361 ( .A(n_314), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_314), .B(n_325), .Y(n_461) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
AND2x2_ASAP7_75t_L g326 ( .A(n_315), .B(n_318), .Y(n_326) );
INVx1_ASAP7_75t_L g335 ( .A(n_315), .Y(n_335) );
AND2x2_ASAP7_75t_L g366 ( .A(n_315), .B(n_319), .Y(n_366) );
INVx1_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g334 ( .A(n_318), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
OR2x2_ASAP7_75t_L g351 ( .A(n_324), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g371 ( .A(n_324), .B(n_354), .Y(n_371) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_325), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g339 ( .A(n_325), .B(n_326), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_325), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_325), .B(n_421), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g446 ( .A1(n_325), .A2(n_437), .B(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_325), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_325), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g406 ( .A(n_326), .Y(n_406) );
AND2x2_ASAP7_75t_L g428 ( .A(n_326), .B(n_392), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_333), .Y(n_327) );
INVx1_ASAP7_75t_L g496 ( .A(n_328), .Y(n_496) );
AND2x2_ASAP7_75t_L g348 ( .A(n_329), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g363 ( .A(n_330), .Y(n_363) );
INVx1_ASAP7_75t_L g430 ( .A(n_330), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_333), .B(n_385), .C(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g417 ( .A(n_334), .B(n_370), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_334), .B(n_454), .Y(n_453) );
OAI32xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .A3(n_344), .B1(n_346), .B2(n_372), .Y(n_336) );
AOI332xp33_ASAP7_75t_L g462 ( .A1(n_337), .A2(n_345), .A3(n_402), .B1(n_408), .B2(n_430), .B3(n_463), .C1(n_465), .C2(n_467), .Y(n_462) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g360 ( .A(n_338), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g437 ( .A(n_338), .B(n_406), .Y(n_437) );
AOI22xp5_ASAP7_75t_SL g347 ( .A1(n_339), .A2(n_348), .B1(n_350), .B2(n_354), .Y(n_347) );
INVx1_ASAP7_75t_L g373 ( .A(n_340), .Y(n_373) );
AND2x2_ASAP7_75t_L g397 ( .A(n_340), .B(n_345), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_340), .A2(n_341), .B1(n_476), .B2(n_484), .Y(n_475) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g390 ( .A1(n_341), .A2(n_391), .B(n_393), .C(n_394), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_SL g432 ( .A1(n_341), .A2(n_433), .B(n_434), .C(n_435), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_341), .A2(n_440), .B(n_450), .C(n_458), .Y(n_439) );
INVx1_ASAP7_75t_L g468 ( .A(n_341), .Y(n_468) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_344), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_345), .A2(n_389), .B1(n_390), .B2(n_397), .C(n_398), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_345), .A2(n_474), .B1(n_475), .B2(n_488), .Y(n_473) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_346), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g346 ( .A(n_347), .B(n_355), .C(n_364), .D(n_367), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_348), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_348), .B(n_358), .Y(n_378) );
INVx1_ASAP7_75t_L g433 ( .A(n_348), .Y(n_433) );
INVx2_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
CKINVDCx6p67_ASAP7_75t_R g413 ( .A(n_349), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_349), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI21xp33_ASAP7_75t_L g482 ( .A1(n_351), .A2(n_357), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g442 ( .A(n_352), .Y(n_442) );
AND2x2_ASAP7_75t_L g381 ( .A(n_353), .B(n_370), .Y(n_381) );
CKINVDCx14_ASAP7_75t_R g483 ( .A(n_354), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_360), .B(n_362), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_356), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx2_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
AND2x2_ASAP7_75t_L g463 ( .A(n_358), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_358), .B(n_361), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g422 ( .A(n_359), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_360), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_361), .A2(n_368), .B(n_371), .Y(n_367) );
AND2x2_ASAP7_75t_L g391 ( .A(n_361), .B(n_392), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_361), .A2(n_371), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_362), .A2(n_407), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g486 ( .A(n_362), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_363), .A2(n_428), .B(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_365), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g421 ( .A(n_366), .B(n_370), .Y(n_421) );
INVx1_ASAP7_75t_L g478 ( .A(n_366), .Y(n_478) );
INVx1_ASAP7_75t_L g447 ( .A(n_368), .Y(n_447) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
OR2x2_ASAP7_75t_L g405 ( .A(n_370), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g460 ( .A(n_370), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g471 ( .A(n_370), .B(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_379), .C(n_382), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_376), .B(n_392), .Y(n_434) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g400 ( .A(n_385), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_393), .B(n_426), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_393), .A2(n_441), .B(n_443), .C(n_444), .Y(n_440) );
INVx2_ASAP7_75t_SL g481 ( .A(n_393), .Y(n_481) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g410 ( .A1(n_397), .A2(n_411), .B(n_432), .C(n_438), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_404), .B2(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_400), .B(n_405), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g458 ( .A1(n_400), .A2(n_459), .B(n_462), .C(n_469), .Y(n_458) );
INVx1_ASAP7_75t_L g464 ( .A(n_401), .Y(n_464) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_406), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g451 ( .A(n_407), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_408), .A2(n_431), .B(n_489), .C(n_490), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_408), .A2(n_481), .B1(n_491), .B2(n_492), .C(n_495), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_439), .C(n_473), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_418), .C(n_427), .Y(n_411) );
CKINVDCx6p67_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g484 ( .A1(n_415), .A2(n_430), .B(n_485), .C(n_486), .Y(n_484) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_416), .B(n_466), .Y(n_485) );
INVx1_ASAP7_75t_L g426 ( .A(n_417), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_423), .B(n_425), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g495 ( .A(n_421), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OAI211xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_453), .C(n_455), .Y(n_450) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_459), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI211xp5_ASAP7_75t_L g476 ( .A1(n_464), .A2(n_477), .B(n_479), .C(n_482), .Y(n_476) );
INVxp67_ASAP7_75t_L g474 ( .A(n_467), .Y(n_474) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g489 ( .A(n_486), .Y(n_489) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx4f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g1527 ( .A(n_500), .B(n_508), .Y(n_1527) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g1570 ( .A(n_502), .B(n_504), .Y(n_1570) );
INVx1_ASAP7_75t_L g1574 ( .A(n_502), .Y(n_1574) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g1577 ( .A(n_504), .B(n_1574), .Y(n_1577) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_510), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g1522 ( .A(n_508), .B(n_1523), .Y(n_1522) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_L g672 ( .A(n_509), .B(n_519), .Y(n_672) );
AND2x4_ASAP7_75t_L g817 ( .A(n_509), .B(n_518), .Y(n_817) );
AND2x4_ASAP7_75t_SL g1526 ( .A(n_510), .B(n_1527), .Y(n_1526) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_517), .Y(n_511) );
BUFx4f_ASAP7_75t_L g955 ( .A(n_512), .Y(n_955) );
INVxp67_ASAP7_75t_L g971 ( .A(n_512), .Y(n_971) );
INVx1_ASAP7_75t_L g1258 ( .A(n_512), .Y(n_1258) );
OR2x6_ASAP7_75t_L g1517 ( .A(n_512), .B(n_1502), .Y(n_1517) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx4f_ASAP7_75t_L g664 ( .A(n_513), .Y(n_664) );
INVx3_ASAP7_75t_L g1107 ( .A(n_513), .Y(n_1107) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g624 ( .A(n_515), .Y(n_624) );
INVx2_ASAP7_75t_L g642 ( .A(n_515), .Y(n_642) );
NAND2x1_ASAP7_75t_L g645 ( .A(n_515), .B(n_516), .Y(n_645) );
AND2x2_ASAP7_75t_L g652 ( .A(n_515), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g660 ( .A(n_515), .B(n_516), .Y(n_660) );
INVx1_ASAP7_75t_L g706 ( .A(n_515), .Y(n_706) );
INVx1_ASAP7_75t_L g625 ( .A(n_516), .Y(n_625) );
AND2x2_ASAP7_75t_L g641 ( .A(n_516), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g653 ( .A(n_516), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_516), .B(n_642), .Y(n_670) );
OR2x2_ASAP7_75t_L g681 ( .A(n_516), .B(n_624), .Y(n_681) );
BUFx2_ASAP7_75t_L g702 ( .A(n_516), .Y(n_702) );
INVxp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g1509 ( .A(n_518), .Y(n_1509) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g1512 ( .A(n_519), .Y(n_1512) );
AND2x4_ASAP7_75t_L g1513 ( .A(n_519), .B(n_705), .Y(n_1513) );
XOR2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_1061), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
XNOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_802), .Y(n_524) );
XNOR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_709), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_707), .B(n_708), .Y(n_526) );
AND3x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_626), .C(n_654), .Y(n_527) );
AOI31xp33_ASAP7_75t_L g708 ( .A1(n_528), .A2(n_626), .A3(n_654), .B(n_707), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_609), .B(n_613), .Y(n_528) );
NAND3xp33_ASAP7_75t_SL g529 ( .A(n_530), .B(n_571), .C(n_587), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_547), .B1(n_559), .B2(n_562), .Y(n_530) );
BUFx2_ASAP7_75t_SL g1134 ( .A(n_532), .Y(n_1134) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_534), .B(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1543 ( .A(n_534), .Y(n_1543) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g565 ( .A(n_535), .Y(n_565) );
INVx8_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g608 ( .A(n_535), .B(n_575), .Y(n_608) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_535), .Y(n_905) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_535), .B(n_1095), .Y(n_1094) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
AND2x4_ASAP7_75t_L g553 ( .A(n_536), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_537), .Y(n_543) );
AND2x4_ASAP7_75t_L g549 ( .A(n_537), .B(n_545), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_537), .B(n_546), .Y(n_599) );
OR2x2_ASAP7_75t_L g754 ( .A(n_537), .B(n_539), .Y(n_754) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_L g554 ( .A(n_540), .Y(n_554) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx5_ASAP7_75t_L g741 ( .A(n_542), .Y(n_741) );
AND2x4_ASAP7_75t_L g800 ( .A(n_542), .B(n_591), .Y(n_800) );
BUFx12f_ASAP7_75t_L g885 ( .A(n_542), .Y(n_885) );
BUFx3_ASAP7_75t_L g1004 ( .A(n_542), .Y(n_1004) );
BUFx3_ASAP7_75t_L g1291 ( .A(n_542), .Y(n_1291) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g574 ( .A(n_543), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_543), .B(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g1481 ( .A(n_543), .Y(n_1481) );
INVx1_ASAP7_75t_L g579 ( .A(n_544), .Y(n_579) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g585 ( .A(n_546), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_548), .A2(n_718), .B1(n_724), .B2(n_725), .Y(n_723) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g563 ( .A(n_549), .Y(n_563) );
BUFx2_ASAP7_75t_L g605 ( .A(n_549), .Y(n_605) );
BUFx2_ASAP7_75t_L g896 ( .A(n_549), .Y(n_896) );
INVx2_ASAP7_75t_L g907 ( .A(n_549), .Y(n_907) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_549), .B(n_1095), .Y(n_1097) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_549), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1476 ( .A(n_549), .B(n_570), .Y(n_1476) );
BUFx2_ASAP7_75t_L g1544 ( .A(n_549), .Y(n_1544) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g1225 ( .A1(n_551), .A2(n_749), .B1(n_1007), .B2(n_1226), .C(n_1227), .Y(n_1225) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g561 ( .A(n_552), .Y(n_561) );
INVx3_ASAP7_75t_L g594 ( .A(n_552), .Y(n_594) );
INVx5_ASAP7_75t_L g910 ( .A(n_552), .Y(n_910) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx8_ASAP7_75t_L g738 ( .A(n_553), .Y(n_738) );
INVx2_ASAP7_75t_L g745 ( .A(n_553), .Y(n_745) );
BUFx6f_ASAP7_75t_L g884 ( .A(n_553), .Y(n_884) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g1436 ( .A(n_556), .B(n_675), .Y(n_1436) );
NAND2xp33_ASAP7_75t_SL g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g576 ( .A(n_557), .Y(n_576) );
AND3x4_ASAP7_75t_L g880 ( .A(n_557), .B(n_766), .C(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_557), .B(n_881), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1495 ( .A(n_557), .Y(n_1495) );
INVx3_ASAP7_75t_L g570 ( .A(n_558), .Y(n_570) );
BUFx3_ASAP7_75t_L g881 ( .A(n_558), .Y(n_881) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g1003 ( .A(n_565), .Y(n_1003) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g746 ( .A1(n_567), .A2(n_747), .B1(n_750), .B2(n_751), .C(n_755), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_567), .A2(n_749), .B1(n_956), .B2(n_968), .C(n_1010), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_567), .A2(n_583), .B1(n_753), .B2(n_1030), .C(n_1031), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g1142 ( .A1(n_567), .A2(n_994), .B1(n_1085), .B2(n_1143), .C(n_1144), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g1230 ( .A1(n_567), .A2(n_749), .B1(n_753), .B2(n_1231), .C(n_1232), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_567), .B(n_1299), .Y(n_1298) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x6_ASAP7_75t_L g915 ( .A(n_568), .B(n_611), .Y(n_915) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND3x1_ASAP7_75t_L g892 ( .A(n_569), .B(n_570), .C(n_893), .Y(n_892) );
AND2x4_ASAP7_75t_L g575 ( .A(n_570), .B(n_576), .Y(n_575) );
OR2x4_ASAP7_75t_L g1468 ( .A(n_570), .B(n_754), .Y(n_1468) );
INVx1_ASAP7_75t_L g1471 ( .A(n_570), .Y(n_1471) );
OR2x6_ASAP7_75t_L g1492 ( .A(n_570), .B(n_598), .Y(n_1492) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B1(n_578), .B2(n_580), .C(n_581), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_572), .A2(n_578), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx4_ASAP7_75t_L g998 ( .A(n_572), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_572), .A2(n_578), .B1(n_581), .B2(n_1183), .C(n_1184), .Y(n_1182) );
AND2x6_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2x1_ASAP7_75t_L g869 ( .A(n_573), .B(n_870), .Y(n_869) );
AND2x2_ASAP7_75t_L g918 ( .A(n_573), .B(n_870), .Y(n_918) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_573), .B(n_870), .Y(n_1342) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_575), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g586 ( .A(n_575), .Y(n_586) );
AND2x4_ASAP7_75t_L g870 ( .A(n_575), .B(n_631), .Y(n_870) );
INVx2_ASAP7_75t_L g999 ( .A(n_578), .Y(n_999) );
INVx1_ASAP7_75t_L g874 ( .A(n_579), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g1000 ( .A(n_581), .B(n_1001), .C(n_1008), .Y(n_1000) );
NOR3xp33_ASAP7_75t_L g1022 ( .A(n_581), .B(n_1023), .C(n_1028), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_582), .Y(n_581) );
OR2x6_ASAP7_75t_L g582 ( .A(n_583), .B(n_586), .Y(n_582) );
INVx1_ASAP7_75t_L g1297 ( .A(n_583), .Y(n_1297) );
INVx1_ASAP7_75t_L g1474 ( .A(n_583), .Y(n_1474) );
BUFx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_584), .Y(n_734) );
BUFx3_ASAP7_75t_L g749 ( .A(n_584), .Y(n_749) );
BUFx2_ASAP7_75t_L g1485 ( .A(n_585), .Y(n_1485) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_593), .B1(n_606), .B2(n_607), .Y(n_587) );
INVxp67_ASAP7_75t_L g722 ( .A(n_588), .Y(n_722) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g996 ( .A(n_590), .Y(n_996) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g744 ( .A(n_591), .Y(n_744) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g850 ( .A(n_592), .B(n_675), .Y(n_850) );
INVx1_ASAP7_75t_L g1095 ( .A(n_592), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_594), .A2(n_1033), .B1(n_1034), .B2(n_1035), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_595), .A2(n_1442), .B1(n_1443), .B2(n_1444), .Y(n_1441) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g761 ( .A(n_599), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_600) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx8_ASAP7_75t_L g724 ( .A(n_603), .Y(n_724) );
INVx2_ASAP7_75t_L g853 ( .A(n_603), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_607), .A2(n_985), .B1(n_993), .B2(n_996), .C(n_997), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g1036 ( .A1(n_607), .A2(n_996), .B1(n_1037), .B2(n_1038), .C(n_1042), .Y(n_1036) );
AOI211xp5_ASAP7_75t_L g1068 ( .A1(n_607), .A2(n_1069), .B(n_1070), .C(n_1071), .Y(n_1068) );
AOI211xp5_ASAP7_75t_L g1128 ( .A1(n_607), .A2(n_1129), .B(n_1130), .C(n_1131), .Y(n_1128) );
INVx2_ASAP7_75t_L g1178 ( .A(n_607), .Y(n_1178) );
AOI211xp5_ASAP7_75t_SL g1233 ( .A1(n_607), .A2(n_1234), .B(n_1235), .C(n_1236), .Y(n_1233) );
AOI211xp5_ASAP7_75t_SL g1274 ( .A1(n_607), .A2(n_1275), .B(n_1276), .C(n_1277), .Y(n_1274) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g715 ( .A(n_608), .B(n_716), .Y(n_715) );
OR2x6_ASAP7_75t_L g878 ( .A(n_608), .B(n_716), .Y(n_878) );
INVx1_ASAP7_75t_L g846 ( .A(n_609), .Y(n_846) );
INVx2_ASAP7_75t_L g1014 ( .A(n_609), .Y(n_1014) );
OAI21xp5_ASAP7_75t_L g1176 ( .A1(n_609), .A2(n_1177), .B(n_1185), .Y(n_1176) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_610), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g692 ( .A(n_611), .B(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_612), .B(n_634), .Y(n_697) );
INVx2_ASAP7_75t_L g766 ( .A(n_612), .Y(n_766) );
INVx1_ASAP7_75t_L g1100 ( .A(n_614), .Y(n_1100) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI222xp33_ASAP7_75t_L g712 ( .A1(n_615), .A2(n_649), .B1(n_713), .B2(n_714), .C1(n_718), .C2(n_719), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_615), .B(n_990), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_615), .B(n_1041), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_615), .B(n_1169), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_615), .A2(n_1147), .B1(n_1180), .B2(n_1197), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_615), .B(n_1261), .Y(n_1260) );
AO211x2_ASAP7_75t_L g1271 ( .A1(n_615), .A2(n_1272), .B(n_1273), .C(n_1302), .Y(n_1271) );
AND2x4_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .Y(n_615) );
AND2x4_ASAP7_75t_L g649 ( .A(n_616), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g703 ( .A(n_617), .B(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g716 ( .A(n_617), .Y(n_716) );
OR2x2_ASAP7_75t_L g979 ( .A(n_617), .B(n_704), .Y(n_979) );
INVx1_ASAP7_75t_L g1523 ( .A(n_617), .Y(n_1523) );
BUFx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g675 ( .A(n_618), .Y(n_675) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_620), .Y(n_842) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_621), .B(n_632), .Y(n_638) );
AND2x2_ASAP7_75t_L g650 ( .A(n_621), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_SL g812 ( .A(n_621), .B(n_659), .Y(n_812) );
AND2x4_ASAP7_75t_L g831 ( .A(n_621), .B(n_782), .Y(n_831) );
AND2x4_ASAP7_75t_L g844 ( .A(n_621), .B(n_651), .Y(n_844) );
HB1xp67_ASAP7_75t_L g1502 ( .A(n_622), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_623), .B(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_623), .Y(n_688) );
INVx3_ASAP7_75t_L g780 ( .A(n_623), .Y(n_780) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_646), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_630), .B(n_799), .Y(n_798) );
AND2x4_ASAP7_75t_L g861 ( .A(n_630), .B(n_862), .Y(n_861) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g982 ( .A(n_631), .Y(n_982) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g893 ( .A(n_632), .Y(n_893) );
INVx1_ASAP7_75t_L g983 ( .A(n_633), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_634), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g828 ( .A(n_634), .Y(n_828) );
AND2x6_ASAP7_75t_L g840 ( .A(n_634), .B(n_659), .Y(n_840) );
AND2x2_ASAP7_75t_L g930 ( .A(n_634), .B(n_931), .Y(n_930) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g717 ( .A(n_636), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g980 ( .A1(n_636), .A2(n_981), .B1(n_984), .B2(n_985), .C1(n_986), .C2(n_988), .Y(n_980) );
AOI222xp33_ASAP7_75t_L g1122 ( .A1(n_636), .A2(n_981), .B1(n_986), .B2(n_1069), .C1(n_1091), .C2(n_1123), .Y(n_1122) );
AOI211xp5_ASAP7_75t_L g1150 ( .A1(n_636), .A2(n_1129), .B(n_1151), .C(n_1152), .Y(n_1150) );
AOI222xp33_ASAP7_75t_L g1199 ( .A1(n_636), .A2(n_981), .B1(n_986), .B2(n_1181), .C1(n_1184), .C2(n_1200), .Y(n_1199) );
AOI222xp33_ASAP7_75t_L g1241 ( .A1(n_636), .A2(n_794), .B1(n_795), .B2(n_1234), .C1(n_1242), .C2(n_1243), .Y(n_1241) );
INVx1_ASAP7_75t_L g1305 ( .A(n_636), .Y(n_1305) );
AND2x4_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AOI332xp33_ASAP7_75t_L g1047 ( .A1(n_637), .A2(n_639), .A3(n_982), .B1(n_983), .B2(n_986), .B3(n_1037), .C1(n_1048), .C2(n_1049), .Y(n_1047) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g643 ( .A(n_638), .B(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g987 ( .A(n_638), .B(n_644), .Y(n_987) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx3_ASAP7_75t_L g689 ( .A(n_641), .Y(n_689) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_641), .Y(n_782) );
BUFx3_ASAP7_75t_L g1326 ( .A(n_641), .Y(n_1326) );
BUFx3_ASAP7_75t_L g967 ( .A(n_644), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_644), .A2(n_1439), .B1(n_1454), .B2(n_1461), .Y(n_1460) );
BUFx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_645), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp33_ASAP7_75t_SL g1015 ( .A(n_649), .B(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1046 ( .A(n_649), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_649), .B(n_1090), .Y(n_1124) );
INVx1_ASAP7_75t_L g1148 ( .A(n_649), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_649), .B(n_1301), .Y(n_1300) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_651), .Y(n_836) );
INVx2_ASAP7_75t_L g1318 ( .A(n_651), .Y(n_1318) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g657 ( .A(n_652), .Y(n_657) );
BUFx3_ASAP7_75t_L g926 ( .A(n_652), .Y(n_926) );
AND2x4_ASAP7_75t_L g1501 ( .A(n_652), .B(n_1502), .Y(n_1501) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_671), .B(n_676), .C(n_698), .Y(n_654) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g1412 ( .A(n_657), .Y(n_1412) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g835 ( .A(n_659), .Y(n_835) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_659), .Y(n_927) );
BUFx3_ASAP7_75t_L g934 ( .A(n_659), .Y(n_934) );
BUFx3_ASAP7_75t_L g1254 ( .A(n_659), .Y(n_1254) );
BUFx3_ASAP7_75t_L g1372 ( .A(n_659), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_659), .B(n_1509), .Y(n_1508) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1158 ( .A(n_660), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_665), .B2(n_666), .Y(n_661) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_664), .Y(n_821) );
INVx4_ASAP7_75t_L g1251 ( .A(n_664), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_666), .A2(n_1444), .B1(n_1448), .B2(n_1464), .Y(n_1463) );
INVx6_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx5_ASAP7_75t_L g1322 ( .A(n_667), .Y(n_1322) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g824 ( .A(n_668), .Y(n_824) );
INVx2_ASAP7_75t_SL g957 ( .A(n_668), .Y(n_957) );
INVx4_ASAP7_75t_L g1252 ( .A(n_668), .Y(n_1252) );
INVx1_ASAP7_75t_L g1458 ( .A(n_668), .Y(n_1458) );
INVx8_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_669), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1520 ( .A(n_669), .B(n_1512), .Y(n_1520) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_671), .Y(n_792) );
AOI222xp33_ASAP7_75t_L g1154 ( .A1(n_671), .A2(n_981), .B1(n_1155), .B2(n_1162), .C1(n_1163), .C2(n_1167), .Y(n_1154) );
AOI222xp33_ASAP7_75t_L g1244 ( .A1(n_671), .A2(n_692), .B1(n_981), .B2(n_1245), .C1(n_1246), .C2(n_1253), .Y(n_1244) );
INVx2_ASAP7_75t_L g1462 ( .A(n_671), .Y(n_1462) );
AND2x4_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx4_ASAP7_75t_L g837 ( .A(n_672), .Y(n_837) );
INVx4_ASAP7_75t_L g935 ( .A(n_672), .Y(n_935) );
AND2x2_ASAP7_75t_SL g975 ( .A(n_672), .B(n_675), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_672), .B(n_673), .Y(n_1054) );
INVx1_ASAP7_75t_SL g1413 ( .A(n_672), .Y(n_1413) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g1497 ( .A(n_675), .Y(n_1497) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_690), .B(n_694), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_682), .B1(n_683), .B2(n_686), .C(n_687), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g813 ( .A1(n_678), .A2(n_814), .B1(n_815), .B2(n_816), .C(n_817), .Y(n_813) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_680), .A2(n_777), .B1(n_1026), .B2(n_1033), .C(n_1053), .Y(n_1052) );
BUFx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g775 ( .A(n_681), .Y(n_775) );
BUFx2_ASAP7_75t_L g787 ( .A(n_681), .Y(n_787) );
INVx1_ASAP7_75t_L g1113 ( .A(n_681), .Y(n_1113) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_681), .Y(n_1115) );
OAI221xp5_ASAP7_75t_L g1213 ( .A1(n_683), .A2(n_785), .B1(n_1187), .B2(n_1214), .C(n_1215), .Y(n_1213) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g960 ( .A(n_684), .Y(n_960) );
INVx4_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OR2x6_ASAP7_75t_L g694 ( .A(n_685), .B(n_695), .Y(n_694) );
BUFx4f_ASAP7_75t_L g777 ( .A(n_685), .Y(n_777) );
BUFx4f_ASAP7_75t_L g788 ( .A(n_685), .Y(n_788) );
BUFx4f_ASAP7_75t_L g814 ( .A(n_685), .Y(n_814) );
BUFx6f_ASAP7_75t_L g1057 ( .A(n_685), .Y(n_1057) );
BUFx4f_ASAP7_75t_L g1506 ( .A(n_685), .Y(n_1506) );
INVx3_ASAP7_75t_L g791 ( .A(n_688), .Y(n_791) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_688), .Y(n_839) );
INVx1_ASAP7_75t_L g1212 ( .A(n_690), .Y(n_1212) );
OAI33xp33_ASAP7_75t_L g1455 ( .A1(n_690), .A2(n_1456), .A3(n_1459), .B1(n_1460), .B2(n_1462), .B3(n_1463), .Y(n_1455) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx4_ASAP7_75t_L g772 ( .A(n_692), .Y(n_772) );
INVx2_ASAP7_75t_L g952 ( .A(n_692), .Y(n_952) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_692), .Y(n_1162) );
OAI21xp5_ASAP7_75t_SL g768 ( .A1(n_694), .A2(n_769), .B(n_773), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_694), .Y(n_1060) );
OAI21xp5_ASAP7_75t_L g1210 ( .A1(n_694), .A2(n_1211), .B(n_1213), .Y(n_1210) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2x2_ASAP7_75t_L g699 ( .A(n_696), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g794 ( .A(n_699), .Y(n_794) );
INVx2_ASAP7_75t_SL g978 ( .A(n_699), .Y(n_978) );
HB1xp67_ASAP7_75t_L g1153 ( .A(n_699), .Y(n_1153) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g827 ( .A(n_702), .Y(n_827) );
BUFx2_ASAP7_75t_L g931 ( .A(n_702), .Y(n_931) );
AND2x4_ASAP7_75t_L g1511 ( .A(n_702), .B(n_1512), .Y(n_1511) );
INVx2_ASAP7_75t_SL g795 ( .A(n_703), .Y(n_795) );
AND2x4_ASAP7_75t_L g848 ( .A(n_703), .B(n_849), .Y(n_848) );
AND2x4_ASAP7_75t_L g943 ( .A(n_703), .B(n_849), .Y(n_943) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_720), .C(n_767), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_742), .B(n_763), .Y(n_720) );
OAI211xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_726), .C(n_729), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_725), .A2(n_727), .B1(n_794), .B2(n_795), .Y(n_793) );
OAI211xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_735), .C(n_739), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_730), .A2(n_750), .B1(n_785), .B2(n_788), .C(n_789), .Y(n_784) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g1192 ( .A1(n_732), .A2(n_1193), .B(n_1194), .C(n_1195), .Y(n_1192) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g995 ( .A(n_733), .Y(n_995) );
INVx3_ASAP7_75t_L g1085 ( .A(n_733), .Y(n_1085) );
INVx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g849 ( .A(n_734), .B(n_850), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g1024 ( .A1(n_734), .A2(n_1007), .B1(n_1025), .B2(n_1026), .C(n_1027), .Y(n_1024) );
INVx4_ASAP7_75t_L g1075 ( .A(n_734), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1287 ( .A(n_734), .Y(n_1287) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_737), .A2(n_959), .B1(n_973), .B2(n_1012), .Y(n_1011) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g757 ( .A(n_738), .Y(n_757) );
INVx3_ASAP7_75t_L g888 ( .A(n_738), .Y(n_888) );
INVx2_ASAP7_75t_SL g1078 ( .A(n_738), .Y(n_1078) );
AND2x4_ASAP7_75t_L g1381 ( .A(n_738), .B(n_854), .Y(n_1381) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_R g911 ( .A(n_741), .Y(n_911) );
INVx2_ASAP7_75t_L g1396 ( .A(n_741), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_743), .Y(n_1089) );
OR2x6_ASAP7_75t_SL g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx3_ASAP7_75t_L g856 ( .A(n_745), .Y(n_856) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_745), .Y(n_1348) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI221xp5_ASAP7_75t_L g1005 ( .A1(n_749), .A2(n_962), .B1(n_966), .B2(n_1006), .C(n_1007), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1440 ( .A(n_749), .Y(n_1440) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
BUFx4f_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
BUFx3_ASAP7_75t_L g994 ( .A(n_754), .Y(n_994) );
BUFx3_ASAP7_75t_L g1010 ( .A(n_754), .Y(n_1010) );
INVx2_ASAP7_75t_L g1402 ( .A(n_754), .Y(n_1402) );
OR2x4_ASAP7_75t_L g1489 ( .A(n_754), .B(n_1471), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_759), .B2(n_762), .Y(n_756) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_757), .A2(n_1007), .B1(n_1085), .B2(n_1137), .C(n_1138), .Y(n_1136) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_758), .A2(n_774), .B1(n_776), .B2(n_777), .C(n_778), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g1445 ( .A1(n_759), .A2(n_1446), .B1(n_1447), .B2(n_1448), .Y(n_1445) );
CKINVDCx8_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
INVx3_ASAP7_75t_L g1012 ( .A(n_760), .Y(n_1012) );
INVx3_ASAP7_75t_L g1034 ( .A(n_760), .Y(n_1034) );
INVx3_ASAP7_75t_L g1188 ( .A(n_760), .Y(n_1188) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g863 ( .A(n_761), .Y(n_863) );
INVx1_ASAP7_75t_L g941 ( .A(n_763), .Y(n_941) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_SL g1067 ( .A1(n_764), .A2(n_1068), .B(n_1088), .C(n_1098), .Y(n_1067) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
HB1xp67_ASAP7_75t_L g1043 ( .A(n_765), .Y(n_1043) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_783), .C(n_796), .Y(n_767) );
INVxp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_SL g1313 ( .A(n_772), .Y(n_1313) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g965 ( .A(n_775), .Y(n_965) );
INVx2_ASAP7_75t_L g1056 ( .A(n_775), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1459 ( .A1(n_777), .A2(n_961), .B1(n_1442), .B2(n_1446), .Y(n_1459) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_SL g1327 ( .A(n_780), .Y(n_1327) );
INVx2_ASAP7_75t_L g1366 ( .A(n_780), .Y(n_1366) );
INVx1_ASAP7_75t_L g1370 ( .A(n_780), .Y(n_1370) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
HB1xp67_ASAP7_75t_L g1415 ( .A(n_782), .Y(n_1415) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx4_ASAP7_75t_L g961 ( .A(n_786), .Y(n_961) );
INVx2_ASAP7_75t_L g1461 ( .A(n_786), .Y(n_1461) );
INVx4_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g937 ( .A(n_791), .Y(n_937) );
AOI222xp33_ASAP7_75t_L g1303 ( .A1(n_794), .A2(n_795), .B1(n_1275), .B2(n_1304), .C1(n_1306), .C2(n_1307), .Y(n_1303) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx3_ASAP7_75t_L g1013 ( .A(n_800), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g1088 ( .A1(n_800), .A2(n_1089), .B1(n_1090), .B2(n_1091), .C(n_1092), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_800), .A2(n_1089), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
XNOR2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_945), .Y(n_802) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_897), .Y(n_803) );
NOR2x1p5_ASAP7_75t_L g805 ( .A(n_806), .B(n_858), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
O2A1O1Ixp33_ASAP7_75t_SL g807 ( .A1(n_808), .A2(n_829), .B(n_846), .C(n_847), .Y(n_807) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g1420 ( .A(n_810), .Y(n_1420) );
INVx4_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx3_ASAP7_75t_L g924 ( .A(n_812), .Y(n_924) );
INVx3_ASAP7_75t_L g928 ( .A(n_817), .Y(n_928) );
INVx1_ASAP7_75t_L g1375 ( .A(n_817), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B1(n_822), .B2(n_823), .Y(n_818) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g1457 ( .A(n_821), .Y(n_1457) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx2_ASAP7_75t_L g1421 ( .A(n_825), .Y(n_1421) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_831), .A2(n_840), .B1(n_900), .B2(n_933), .C(n_936), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g1363 ( .A1(n_831), .A2(n_840), .B1(n_1337), .B2(n_1364), .C(n_1365), .Y(n_1363) );
INVx2_ASAP7_75t_SL g1407 ( .A(n_831), .Y(n_1407) );
AOI221xp5_ASAP7_75t_L g1554 ( .A1(n_831), .A2(n_840), .B1(n_1534), .B2(n_1555), .C(n_1559), .Y(n_1554) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_838), .B(n_840), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
BUFx3_ASAP7_75t_L g1159 ( .A(n_836), .Y(n_1159) );
AOI21xp5_ASAP7_75t_L g1408 ( .A1(n_840), .A2(n_1409), .B(n_1414), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_842), .A2(n_844), .B1(n_939), .B2(n_940), .Y(n_938) );
HB1xp67_ASAP7_75t_L g1360 ( .A(n_842), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_842), .A2(n_844), .B1(n_1417), .B2(n_1418), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_842), .A2(n_1362), .B1(n_1552), .B2(n_1553), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_843), .A2(n_845), .B1(n_852), .B2(n_855), .Y(n_851) );
BUFx6f_ASAP7_75t_L g1362 ( .A(n_844), .Y(n_1362) );
A2O1A1Ixp33_ASAP7_75t_SL g1127 ( .A1(n_846), .A2(n_1128), .B(n_1132), .C(n_1145), .Y(n_1127) );
AOI21xp5_ASAP7_75t_SL g1549 ( .A1(n_846), .A2(n_1550), .B(n_1564), .Y(n_1549) );
INVx1_ASAP7_75t_L g854 ( .A(n_850), .Y(n_854) );
INVx1_ASAP7_75t_L g857 ( .A(n_850), .Y(n_857) );
OR2x2_ASAP7_75t_L g862 ( .A(n_850), .B(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_852), .A2(n_855), .B1(n_939), .B2(n_940), .Y(n_944) );
AND2x4_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
AND2x4_ASAP7_75t_L g1380 ( .A(n_853), .B(n_854), .Y(n_1380) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
INVx2_ASAP7_75t_L g1006 ( .A(n_856), .Y(n_1006) );
INVx2_ASAP7_75t_L g1039 ( .A(n_856), .Y(n_1039) );
INVxp67_ASAP7_75t_L g1403 ( .A(n_857), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_865), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_864), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_860), .A2(n_877), .B1(n_900), .B2(n_901), .C(n_902), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g1336 ( .A1(n_860), .A2(n_877), .B1(n_1337), .B2(n_1338), .C(n_1339), .Y(n_1336) );
AOI21xp33_ASAP7_75t_L g1385 ( .A1(n_860), .A2(n_1386), .B(n_1387), .Y(n_1385) );
AOI221xp5_ASAP7_75t_L g1533 ( .A1(n_860), .A2(n_877), .B1(n_1534), .B2(n_1535), .C(n_1536), .Y(n_1533) );
INVx8_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1081 ( .A(n_863), .Y(n_1081) );
AND4x1_ASAP7_75t_L g865 ( .A(n_866), .B(n_875), .C(n_879), .D(n_894), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B1(n_871), .B2(n_872), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_868), .A2(n_920), .B1(n_1538), .B2(n_1539), .Y(n_1537) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AND2x4_ASAP7_75t_SL g872 ( .A(n_870), .B(n_873), .Y(n_872) );
AND2x4_ASAP7_75t_L g895 ( .A(n_870), .B(n_896), .Y(n_895) );
AND2x4_ASAP7_75t_L g920 ( .A(n_870), .B(n_873), .Y(n_920) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
INVx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AOI33xp33_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_882), .A3(n_883), .B1(n_886), .B2(n_889), .B3(n_890), .Y(n_879) );
AOI33xp33_ASAP7_75t_L g903 ( .A1(n_880), .A2(n_904), .A3(n_908), .B1(n_912), .B2(n_913), .B3(n_914), .Y(n_903) );
BUFx3_ASAP7_75t_L g1354 ( .A(n_880), .Y(n_1354) );
AOI33xp33_ASAP7_75t_L g1393 ( .A1(n_880), .A2(n_914), .A3(n_1394), .B1(n_1395), .B2(n_1397), .B3(n_1398), .Y(n_1393) );
INVx3_ASAP7_75t_L g1480 ( .A(n_881), .Y(n_1480) );
INVx2_ASAP7_75t_L g1027 ( .A(n_884), .Y(n_1027) );
BUFx6f_ASAP7_75t_L g1141 ( .A(n_884), .Y(n_1141) );
BUFx6f_ASAP7_75t_L g1283 ( .A(n_884), .Y(n_1283) );
INVx1_ASAP7_75t_L g1447 ( .A(n_884), .Y(n_1447) );
AND2x4_ASAP7_75t_L g1470 ( .A(n_884), .B(n_1471), .Y(n_1470) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_885), .Y(n_1135) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
BUFx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
BUFx2_ASAP7_75t_L g1350 ( .A(n_891), .Y(n_1350) );
BUFx2_ASAP7_75t_L g1547 ( .A(n_891), .Y(n_1547) );
INVx3_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx3_ASAP7_75t_L g1450 ( .A(n_892), .Y(n_1450) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_894), .B(n_903), .C(n_916), .Y(n_902) );
INVx3_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx3_ASAP7_75t_L g1344 ( .A(n_895), .Y(n_1344) );
NOR3xp33_ASAP7_75t_L g1388 ( .A(n_895), .B(n_1389), .C(n_1399), .Y(n_1388) );
AND2x2_ASAP7_75t_L g898 ( .A(n_899), .B(n_921), .Y(n_898) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx8_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_910), .A2(n_1187), .B1(n_1188), .B2(n_1189), .C(n_1190), .Y(n_1186) );
BUFx3_ASAP7_75t_L g1443 ( .A(n_910), .Y(n_1443) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_916) );
AOI222xp33_ASAP7_75t_L g923 ( .A1(n_917), .A2(n_919), .B1(n_924), .B2(n_925), .C1(n_929), .C2(n_930), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_918), .A2(n_920), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_920), .A2(n_1341), .B1(n_1342), .B2(n_1343), .Y(n_1340) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_941), .B(n_942), .Y(n_921) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_932), .C(n_938), .Y(n_922) );
AOI222xp33_ASAP7_75t_L g1368 ( .A1(n_924), .A2(n_1341), .B1(n_1343), .B2(n_1369), .C1(n_1371), .C2(n_1376), .Y(n_1368) );
AOI222xp33_ASAP7_75t_L g1560 ( .A1(n_924), .A2(n_1376), .B1(n_1538), .B2(n_1539), .C1(n_1561), .C2(n_1563), .Y(n_1560) );
INVx1_ASAP7_75t_L g1206 ( .A(n_926), .Y(n_1206) );
INVx1_ASAP7_75t_L g1248 ( .A(n_926), .Y(n_1248) );
BUFx2_ASAP7_75t_L g1324 ( .A(n_926), .Y(n_1324) );
INVx1_ASAP7_75t_L g1377 ( .A(n_930), .Y(n_1377) );
OAI21xp5_ASAP7_75t_L g1405 ( .A1(n_941), .A2(n_1406), .B(n_1419), .Y(n_1405) );
XNOR2x1_ASAP7_75t_L g945 ( .A(n_946), .B(n_1017), .Y(n_945) );
XNOR2x1_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
NOR2x1_ASAP7_75t_L g948 ( .A(n_949), .B(n_991), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_980), .C(n_989), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g950 ( .A(n_951), .B(n_976), .Y(n_950) );
OAI33xp33_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .A3(n_958), .B1(n_963), .B2(n_969), .B3(n_974), .Y(n_951) );
OAI22xp5_ASAP7_75t_SL g1051 ( .A1(n_952), .A2(n_1052), .B1(n_1054), .B2(n_1055), .Y(n_1051) );
OAI33xp33_ASAP7_75t_L g1103 ( .A1(n_952), .A2(n_1104), .A3(n_1110), .B1(n_1114), .B2(n_1116), .B3(n_1120), .Y(n_1103) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_955), .A2(n_1109), .B1(n_1165), .B2(n_1166), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_955), .A2(n_1320), .B1(n_1321), .B2(n_1322), .Y(n_1319) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_957), .A2(n_970), .B1(n_972), .B2(n_973), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_957), .A2(n_1256), .B1(n_1257), .B2(n_1259), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_960), .B1(n_961), .B2(n_962), .Y(n_958) );
OAI211xp5_ASAP7_75t_SL g1422 ( .A1(n_960), .A2(n_1423), .B(n_1424), .C(n_1425), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_963) );
INVx4_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_967), .A2(n_1079), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1160 ( .A1(n_970), .A2(n_1109), .B1(n_1144), .B2(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g1120 ( .A(n_975), .Y(n_1120) );
INVx2_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AOI21xp33_ASAP7_75t_L g1328 ( .A1(n_981), .A2(n_1060), .B(n_1329), .Y(n_1328) );
AND2x4_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
AOI21xp5_ASAP7_75t_L g1262 ( .A1(n_986), .A2(n_1060), .B(n_1263), .Y(n_1262) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
A2O1A1Ixp33_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_1000), .B(n_1014), .C(n_1015), .Y(n_991) );
OAI22xp33_ASAP7_75t_L g1437 ( .A1(n_994), .A2(n_1438), .B1(n_1439), .B2(n_1440), .Y(n_1437) );
OAI22xp33_ASAP7_75t_L g1451 ( .A1(n_994), .A2(n_1452), .B1(n_1453), .B2(n_1454), .Y(n_1451) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1007), .Y(n_1289) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1010), .Y(n_1296) );
A2O1A1Ixp33_ASAP7_75t_L g1221 ( .A1(n_1014), .A2(n_1222), .B(n_1233), .C(n_1237), .Y(n_1221) );
AOI21xp5_ASAP7_75t_L g1356 ( .A1(n_1014), .A2(n_1357), .B(n_1378), .Y(n_1356) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
XNOR2x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1045), .Y(n_1020) );
A2O1A1Ixp33_ASAP7_75t_L g1021 ( .A1(n_1022), .A2(n_1036), .B(n_1043), .C(n_1044), .Y(n_1021) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_1025), .A2(n_1030), .B1(n_1056), .B2(n_1057), .C(n_1058), .Y(n_1055) );
A2O1A1Ixp33_ASAP7_75t_SL g1273 ( .A1(n_1043), .A2(n_1274), .B(n_1278), .C(n_1300), .Y(n_1273) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1046), .Y(n_1239) );
NOR3xp33_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1059), .C(n_1060), .Y(n_1050) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1054), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_1057), .A2(n_1073), .B1(n_1084), .B2(n_1115), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_1062), .A2(n_1266), .B1(n_1267), .B2(n_1428), .Y(n_1061) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1062), .Y(n_1428) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1172), .B1(n_1264), .B2(n_1265), .Y(n_1062) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1063), .Y(n_1264) );
OA22x2_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1125), .B1(n_1170), .B2(n_1171), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
BUFx2_ASAP7_75t_SL g1171 ( .A(n_1065), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1101), .Y(n_1066) );
OAI21xp33_ASAP7_75t_L g1071 ( .A1(n_1072), .A2(n_1077), .B(n_1083), .Y(n_1071) );
OAI21xp33_ASAP7_75t_L g1072 ( .A1(n_1073), .A2(n_1074), .B(n_1076), .Y(n_1072) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1075), .Y(n_1453) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1079), .B1(n_1080), .B2(n_1082), .Y(n_1077) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1078), .Y(n_1229) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_1082), .A2(n_1109), .B1(n_1117), .B2(n_1119), .Y(n_1116) );
OAI211xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1085), .B(n_1086), .C(n_1087), .Y(n_1083) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1094), .A2(n_1097), .B1(n_1197), .B2(n_1198), .Y(n_1196) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1100), .Y(n_1098) );
NAND3xp33_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1122), .C(n_1124), .Y(n_1101) );
NOR2xp33_ASAP7_75t_SL g1102 ( .A(n_1103), .B(n_1121), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1106), .B1(n_1108), .B2(n_1109), .Y(n_1104) );
BUFx6f_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1107), .Y(n_1118) );
BUFx3_ASAP7_75t_L g1464 ( .A(n_1107), .Y(n_1464) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1125), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1149), .Y(n_1126) );
NOR3xp33_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1139), .C(n_1140), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1147), .Y(n_1145) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
NAND3xp33_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1154), .C(n_1168), .Y(n_1149) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1157), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1158), .Y(n_1558) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1172), .Y(n_1265) );
XOR2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1219), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1175), .Y(n_1217) );
NAND4xp25_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1199), .C(n_1201), .D(n_1216), .Y(n_1175) );
NAND3xp33_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1192), .C(n_1196), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1210), .Y(n_1201) );
NAND3xp33_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1208), .C(n_1209), .Y(n_1203) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1240), .Y(n_1220) );
NOR3xp33_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .C(n_1228), .Y(n_1222) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_1232), .A2(n_1250), .B1(n_1251), .B2(n_1252), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1239), .Y(n_1237) );
NAND4xp25_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1244), .C(n_1260), .D(n_1262), .Y(n_1240) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1269), .B1(n_1330), .B2(n_1331), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
HB1xp67_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NOR3xp33_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1292), .C(n_1293), .Y(n_1278) );
NOR3xp33_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1284), .C(n_1290), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1281), .B(n_1311), .Y(n_1315) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1288), .Y(n_1284) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
NAND3xp33_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1308), .C(n_1328), .Y(n_1302) );
INVxp67_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1314), .B1(n_1323), .B2(n_1325), .Y(n_1308) );
AOI22xp5_ASAP7_75t_L g1314 ( .A1(n_1310), .A2(n_1315), .B1(n_1316), .B2(n_1319), .Y(n_1314) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1317), .Y(n_1374) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
BUFx3_ASAP7_75t_L g1367 ( .A(n_1326), .Y(n_1367) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AO22x1_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1382), .B1(n_1426), .B2(n_1427), .Y(n_1331) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1332), .Y(n_1426) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
NAND2xp67_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1356), .Y(n_1335) );
NAND3xp33_ASAP7_75t_SL g1339 ( .A(n_1340), .B(n_1344), .C(n_1345), .Y(n_1339) );
NAND3xp33_ASAP7_75t_SL g1536 ( .A(n_1344), .B(n_1537), .C(n_1540), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1349), .B1(n_1352), .B2(n_1355), .Y(n_1345) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
AOI33xp33_ASAP7_75t_L g1540 ( .A1(n_1354), .A2(n_1541), .A3(n_1545), .B1(n_1546), .B2(n_1547), .B3(n_1548), .Y(n_1540) );
NAND3xp33_ASAP7_75t_SL g1357 ( .A(n_1358), .B(n_1363), .C(n_1368), .Y(n_1357) );
AOI22xp5_ASAP7_75t_L g1358 ( .A1(n_1359), .A2(n_1360), .B1(n_1361), .B2(n_1362), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_1359), .A2(n_1361), .B1(n_1380), .B2(n_1381), .Y(n_1379) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_1380), .A2(n_1381), .B1(n_1552), .B2(n_1553), .Y(n_1565) );
INVx2_ASAP7_75t_L g1404 ( .A(n_1381), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1383), .Y(n_1427) );
NAND3xp33_ASAP7_75t_SL g1384 ( .A(n_1385), .B(n_1388), .C(n_1405), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1393), .Y(n_1389) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1403), .Y(n_1400) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_1402), .Y(n_1401) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx2_ASAP7_75t_L g1562 ( .A(n_1411), .Y(n_1562) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
OAI222xp33_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1524), .B1(n_1528), .B2(n_1566), .C1(n_1571), .C2(n_1578), .Y(n_1429) );
HB1xp67_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
NAND3xp33_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1465), .C(n_1498), .Y(n_1432) );
NOR2xp33_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1455), .Y(n_1433) );
OAI33xp33_ASAP7_75t_L g1434 ( .A1(n_1435), .A2(n_1437), .A3(n_1441), .B1(n_1445), .B2(n_1449), .B3(n_1451), .Y(n_1434) );
BUFx8_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
OAI22xp33_ASAP7_75t_L g1456 ( .A1(n_1438), .A2(n_1452), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_1450), .Y(n_1449) );
OAI31xp33_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1472), .A3(n_1487), .B(n_1493), .Y(n_1465) );
HB1xp67_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
CKINVDCx8_ASAP7_75t_R g1475 ( .A(n_1476), .Y(n_1475) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1482), .B1(n_1483), .B2(n_1486), .Y(n_1477) );
BUFx3_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1481), .Y(n_1479) );
AND2x4_ASAP7_75t_L g1484 ( .A(n_1480), .B(n_1485), .Y(n_1484) );
AOI22xp33_ASAP7_75t_SL g1510 ( .A1(n_1482), .A2(n_1511), .B1(n_1513), .B2(n_1514), .Y(n_1510) );
BUFx6f_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
BUFx3_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1496), .Y(n_1493) );
INVx1_ASAP7_75t_SL g1494 ( .A(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
OAI31xp33_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1503), .A3(n_1515), .B(n_1521), .Y(n_1498) );
INVx3_ASAP7_75t_SL g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
BUFx6f_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx2_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
BUFx2_ASAP7_75t_SL g1521 ( .A(n_1522), .Y(n_1521) );
INVx3_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
BUFx3_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
HB1xp67_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1549), .Y(n_1532) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
NAND3xp33_ASAP7_75t_SL g1550 ( .A(n_1551), .B(n_1554), .C(n_1560), .Y(n_1550) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
CKINVDCx5p33_ASAP7_75t_R g1566 ( .A(n_1567), .Y(n_1566) );
HB1xp67_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
BUFx3_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
BUFx3_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
HB1xp67_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
OAI21xp5_ASAP7_75t_L g1573 ( .A1(n_1574), .A2(n_1575), .B(n_1576), .Y(n_1573) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
endmodule