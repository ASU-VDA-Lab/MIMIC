module fake_jpeg_11897_n_197 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_86),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_71),
.B1(n_74),
.B2(n_63),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_80),
.B1(n_69),
.B2(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_101),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_80),
.B1(n_69),
.B2(n_75),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_65),
.B1(n_71),
.B2(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_63),
.B1(n_77),
.B2(n_54),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_77),
.B1(n_58),
.B2(n_62),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_81),
.B1(n_79),
.B2(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_59),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_59),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_90),
.B1(n_60),
.B2(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_116),
.B1(n_115),
.B2(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_118),
.B1(n_6),
.B2(n_8),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_92),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_98),
.B(n_5),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_126),
.Y(n_139)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_24),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_132),
.B(n_145),
.Y(n_166)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_11),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_12),
.B(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_14),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_148),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_23),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_25),
.C(n_26),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_29),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_32),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_33),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_34),
.B(n_36),
.C(n_37),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_131),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_176),
.Y(n_183)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_147),
.B(n_141),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_179),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_38),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_151),
.B1(n_165),
.B2(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_181),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_151),
.B1(n_130),
.B2(n_145),
.Y(n_181)
);

INVxp33_ASAP7_75t_SL g182 ( 
.A(n_172),
.Y(n_182)
);

OAI31xp33_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_170),
.A3(n_175),
.B(n_158),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_155),
.B(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_177),
.C(n_169),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_183),
.B1(n_186),
.B2(n_182),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_184),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_40),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_41),
.B(n_44),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_48),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_49),
.Y(n_197)
);


endmodule