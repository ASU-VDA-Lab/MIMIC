module fake_jpeg_28001_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_SL g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_57),
.Y(n_81)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_37),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_73),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_71),
.B(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_28),
.B1(n_19),
.B2(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_74),
.B1(n_84),
.B2(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_20),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_28),
.B1(n_19),
.B2(n_33),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_31),
.B1(n_39),
.B2(n_22),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_88),
.B1(n_21),
.B2(n_46),
.Y(n_122)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_83),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_31),
.B1(n_25),
.B2(n_29),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_92),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_32),
.B1(n_29),
.B2(n_21),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_41),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_102),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_37),
.C(n_49),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_76),
.B1(n_86),
.B2(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_126),
.B1(n_83),
.B2(n_87),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_40),
.C(n_41),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_112),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_18),
.B1(n_26),
.B2(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_115),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_64),
.B1(n_63),
.B2(n_60),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_122),
.B1(n_46),
.B2(n_35),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_26),
.B(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_69),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_127),
.B(n_133),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_134),
.B1(n_137),
.B2(n_98),
.Y(n_170)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_75),
.B1(n_89),
.B2(n_66),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_139),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_10),
.Y(n_136)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_11),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_70),
.B1(n_92),
.B2(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_24),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_93),
.B1(n_70),
.B2(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_59),
.B1(n_68),
.B2(n_120),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_155),
.B1(n_99),
.B2(n_97),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_23),
.B1(n_32),
.B2(n_17),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_119),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_126),
.C(n_100),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_166),
.C(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_176),
.B1(n_145),
.B2(n_146),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_106),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_183),
.B(n_143),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_122),
.B1(n_114),
.B2(n_103),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_16),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_114),
.C(n_108),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_97),
.B1(n_115),
.B2(n_121),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_125),
.B1(n_116),
.B2(n_98),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_177),
.B1(n_186),
.B2(n_172),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_127),
.B(n_15),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_184),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_116),
.B1(n_23),
.B2(n_69),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_42),
.C(n_96),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_42),
.C(n_80),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_152),
.A2(n_46),
.B(n_27),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_153),
.C(n_139),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_32),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_189),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_143),
.A2(n_59),
.B1(n_43),
.B2(n_17),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_43),
.A3(n_35),
.B1(n_24),
.B2(n_27),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_80),
.C(n_61),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_148),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_190),
.B(n_204),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_193),
.B(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_169),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_203),
.B1(n_211),
.B2(n_217),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_218),
.B1(n_186),
.B2(n_160),
.Y(n_227)
);

CKINVDCx10_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_210),
.B(n_213),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_145),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_205),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_182),
.B(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_129),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_209),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_156),
.B(n_130),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_164),
.B(n_149),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_140),
.B1(n_61),
.B2(n_80),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_212),
.B(n_215),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_140),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_12),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_27),
.B1(n_16),
.B2(n_12),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_243),
.B1(n_189),
.B2(n_217),
.Y(n_264)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_234),
.Y(n_260)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_183),
.B(n_165),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_158),
.B1(n_178),
.B2(n_188),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_196),
.B1(n_157),
.B2(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_239),
.Y(n_262)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_210),
.A2(n_195),
.B(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_218),
.B1(n_196),
.B2(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_255),
.B1(n_264),
.B2(n_223),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_191),
.C(n_206),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_254),
.C(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_257),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_191),
.C(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_205),
.C(n_179),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_194),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_239),
.B(n_219),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_265),
.B(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_202),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_228),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_269),
.B(n_271),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_228),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_282),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_234),
.C(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_279),
.C(n_283),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_280),
.B1(n_286),
.B2(n_2),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_226),
.C(n_238),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_232),
.B1(n_229),
.B2(n_226),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_224),
.B(n_222),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_1),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_260),
.B(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_231),
.C(n_227),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_222),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_266),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_262),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_1),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_240),
.B1(n_194),
.B2(n_242),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_268),
.B1(n_248),
.B2(n_263),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_300),
.B1(n_5),
.B2(n_7),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_2),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_253),
.C(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_298),
.Y(n_303)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_252),
.B(n_261),
.C(n_262),
.D(n_248),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

AO221x1_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_251),
.B1(n_249),
.B2(n_161),
.C(n_180),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_293),
.B(n_295),
.Y(n_306)
);

OAI322xp33_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_251),
.A3(n_161),
.B1(n_159),
.B2(n_11),
.C1(n_4),
.C2(n_5),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_11),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_299),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_270),
.B1(n_276),
.B2(n_272),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_3),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_274),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_289),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_284),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_298),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_313),
.B1(n_291),
.B2(n_7),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_9),
.C(n_6),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_5),
.C(n_7),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_320),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_294),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_7),
.B(n_8),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_307),
.B(n_304),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_306),
.B(n_309),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_314),
.B1(n_302),
.B2(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_8),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_331),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_328),
.C(n_324),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_325),
.C(n_330),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

XNOR2x2_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_9),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_9),
.Y(n_338)
);


endmodule