module real_jpeg_10649_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_48),
.B1(n_52),
.B2(n_64),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_45),
.B1(n_50),
.B2(n_53),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_4),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_50),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_4),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_4),
.A2(n_45),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_6),
.B(n_23),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_6),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_24),
.B(n_42),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_82),
.B1(n_84),
.B2(n_109),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_31),
.B(n_58),
.C(n_66),
.D(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_6),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_6),
.B(n_27),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_6),
.A2(n_46),
.B(n_135),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_23),
.B(n_36),
.C(n_71),
.D(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_10),
.A2(n_48),
.B1(n_52),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_10),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_28),
.B1(n_31),
.B2(n_51),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_13),
.A2(n_35),
.B1(n_48),
.B2(n_52),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_13),
.A2(n_35),
.B1(n_84),
.B2(n_109),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_14),
.A2(n_25),
.B1(n_48),
.B2(n_52),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_115),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_77),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_18),
.B(n_77),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_56),
.C(n_69),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_19),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_38),
.B2(n_55),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_39),
.C(n_44),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_32),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_22),
.A2(n_26),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_27),
.B(n_29),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_26),
.B(n_34),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_28),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_59),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_31),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_40),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_41),
.A2(n_43),
.B(n_84),
.C(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_82),
.B(n_83),
.C(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_43),
.B(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_47),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_46),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_47),
.A2(n_141),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_47),
.B(n_82),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_48),
.A2(n_61),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_52),
.B(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_52),
.B(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_53),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_56),
.B(n_69),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_63),
.B(n_65),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_57),
.A2(n_63),
.B1(n_67),
.B2(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_97),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_67),
.B(n_82),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_70),
.B(n_74),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_75),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_93),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_90),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_110),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_170),
.B(n_174),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_157),
.B(n_169),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_137),
.B(n_156),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_119),
.B(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_131),
.C(n_133),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_134),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_145),
.B(n_155),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_154),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_159),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_167),
.B2(n_168),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_171),
.B(n_172),
.Y(n_174)
);


endmodule