module real_jpeg_32990_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_666;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_605;
wire n_216;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_689;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_431;
wire n_357;
wire n_420;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_686;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_468;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_0),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_0),
.Y(n_401)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_0),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_1),
.A2(n_121),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_1),
.A2(n_121),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_1),
.A2(n_121),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_2),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_2),
.A2(n_131),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_2),
.A2(n_131),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_2),
.A2(n_131),
.B1(n_344),
.B2(n_347),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_3),
.A2(n_123),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_3),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_3),
.A2(n_362),
.B1(n_464),
.B2(n_468),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_3),
.A2(n_362),
.B1(n_558),
.B2(n_560),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_3),
.A2(n_362),
.B1(n_626),
.B2(n_630),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_5),
.A2(n_27),
.B1(n_138),
.B2(n_145),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_5),
.A2(n_27),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_5),
.A2(n_27),
.B1(n_303),
.B2(n_306),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_6),
.A2(n_285),
.B1(n_286),
.B2(n_289),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_6),
.A2(n_285),
.B1(n_390),
.B2(n_394),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_6),
.A2(n_232),
.B1(n_285),
.B2(n_512),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_6),
.A2(n_285),
.B1(n_604),
.B2(n_605),
.Y(n_603)
);

OAI22x1_ASAP7_75t_SL g268 ( 
.A1(n_7),
.A2(n_129),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_7),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_7),
.A2(n_269),
.B1(n_369),
.B2(n_371),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_7),
.A2(n_269),
.B1(n_448),
.B2(n_451),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_7),
.A2(n_269),
.B1(n_539),
.B2(n_544),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_67),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_60),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_8),
.A2(n_60),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

AO22x1_ASAP7_75t_SL g250 ( 
.A1(n_8),
.A2(n_60),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_11),
.Y(n_247)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_11),
.Y(n_543)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_12),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_13),
.A2(n_208),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_13),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_13),
.A2(n_212),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_13),
.A2(n_212),
.B1(n_355),
.B2(n_357),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_13),
.A2(n_212),
.B1(n_483),
.B2(n_486),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_14),
.B(n_678),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_14),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_15),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_16),
.B(n_47),
.Y(n_422)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_16),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_16),
.B(n_72),
.Y(n_490)
);

OAI32xp33_ASAP7_75t_L g516 ( 
.A1(n_16),
.A2(n_517),
.A3(n_520),
.B1(n_522),
.B2(n_529),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_16),
.A2(n_459),
.B1(n_552),
.B2(n_555),
.Y(n_551)
);

OAI21xp33_ASAP7_75t_L g641 ( 
.A1(n_16),
.A2(n_307),
.B(n_607),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_18),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_18),
.Y(n_148)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_18),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_681),
.C(n_686),
.Y(n_19)
);

AOI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_190),
.A3(n_666),
.B1(n_679),
.B2(n_680),
.Y(n_20)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_21),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_21),
.A2(n_676),
.B1(n_687),
.B2(n_689),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_189),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_73),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_25),
.B(n_73),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B1(n_59),
.B2(n_72),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_26),
.A2(n_35),
.B1(n_72),
.B2(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_31),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_31),
.Y(n_130)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_31),
.Y(n_274)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_34),
.Y(n_417)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_35),
.A2(n_72),
.B1(n_117),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_37),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_37),
.B(n_284),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g360 ( 
.A1(n_37),
.A2(n_72),
.B1(n_284),
.B2(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_37),
.B(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_46),
.Y(n_37)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

AOI22x1_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_38)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_40),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_40),
.Y(n_393)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_42),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_42),
.Y(n_428)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_45),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_53),
.B2(n_57),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_54),
.Y(n_365)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_56),
.Y(n_211)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_72),
.B(n_207),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_72),
.B(n_268),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_72),
.B(n_361),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_185),
.C(n_187),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_74),
.B(n_671),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_115),
.C(n_135),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_75),
.A2(n_76),
.B1(n_135),
.B2(n_136),
.Y(n_217)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_76),
.B(n_196),
.C(n_205),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_76),
.B(n_196),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_93),
.B(n_106),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_77),
.A2(n_93),
.B1(n_106),
.B2(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_77),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_77),
.A2(n_93),
.B1(n_447),
.B2(n_453),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_77),
.B(n_447),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_95),
.Y(n_94)
);

OAI22x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_81),
.Y(n_251)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_81),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_86),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_86),
.Y(n_408)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_86),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_87),
.Y(n_254)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_87),
.Y(n_406)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_87),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_87),
.Y(n_546)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_93),
.B(n_596),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_93),
.B(n_447),
.Y(n_612)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_94),
.A2(n_231),
.B1(n_257),
.B2(n_264),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_94),
.A2(n_257),
.B1(n_264),
.B2(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_94),
.A2(n_264),
.B1(n_312),
.B2(n_354),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_94),
.A2(n_511),
.B(n_514),
.Y(n_510)
);

OAI22xp33_ASAP7_75t_L g556 ( 
.A1(n_94),
.A2(n_264),
.B1(n_511),
.B2(n_557),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_96),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_98),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_98),
.Y(n_521)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_103),
.Y(n_313)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_104),
.Y(n_450)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_105),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_105),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_108),
.Y(n_356)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_108),
.Y(n_452)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_114),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_115),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_126),
.B1(n_127),
.B2(n_134),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_125),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx4f_ASAP7_75t_SL g213 ( 
.A(n_130),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22x1_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_149),
.B1(n_174),
.B2(n_181),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_137),
.A2(n_151),
.B1(n_181),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_143),
.Y(n_228)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_143),
.Y(n_296)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_143),
.Y(n_370)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_144),
.Y(n_554)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_147),
.Y(n_555)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_148),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_174),
.B(n_181),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_149),
.A2(n_181),
.B1(n_197),
.B2(n_225),
.Y(n_224)
);

AOI22x1_ASAP7_75t_L g461 ( 
.A1(n_149),
.A2(n_181),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g366 ( 
.A1(n_150),
.A2(n_182),
.B1(n_367),
.B2(n_372),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_150),
.A2(n_389),
.B(n_396),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_150),
.A2(n_396),
.B(n_551),
.Y(n_550)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_151),
.A2(n_183),
.B1(n_225),
.B2(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_151),
.B(n_368),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_161),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_157),
.B1(n_159),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_156),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_168),
.B2(n_173),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_163),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_164),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_164),
.Y(n_472)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_182),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_182),
.B(n_459),
.Y(n_610)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_183),
.B(n_368),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g671 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_672),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_185),
.Y(n_672)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_190),
.Y(n_685)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_328),
.B(n_661),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_276),
.Y(n_192)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_193),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_219),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_194),
.B(n_219),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_214),
.Y(n_194)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_195),
.Y(n_675)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_221),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_206),
.A2(n_221),
.B(n_222),
.C(n_326),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_206),
.Y(n_327)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_216),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_218),
.B(n_674),
.C(n_675),
.Y(n_673)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_238),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_220),
.A2(n_222),
.B(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_221),
.A2(n_223),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_224),
.B(n_229),
.Y(n_279)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx4f_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_255),
.B(n_265),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_239),
.A2(n_240),
.B1(n_266),
.B2(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_239),
.A2(n_240),
.B1(n_256),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_256),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_244),
.B(n_250),
.Y(n_240)
);

BUFx2_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_242),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_243),
.Y(n_639)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

AO22x1_ASAP7_75t_SL g399 ( 
.A1(n_244),
.A2(n_343),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_244),
.B(n_538),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_244),
.A2(n_400),
.B1(n_624),
.B2(n_632),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_246),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_247),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_247),
.Y(n_488)
);

INVx4_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g536 ( 
.A(n_249),
.Y(n_536)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_256),
.Y(n_374)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_262),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_263),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_263),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_264),
.A2(n_557),
.B(n_612),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_264),
.B(n_459),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_266),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_275),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_267),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_323),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_277),
.B(n_323),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_319),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_279),
.B(n_320),
.Y(n_376)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g375 ( 
.A(n_281),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_292),
.C(n_299),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_282),
.A2(n_293),
.B1(n_294),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_291),
.Y(n_282)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_291),
.B(n_455),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_311),
.Y(n_300)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_301),
.B(n_430),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_307),
.B1(n_342),
.B2(n_350),
.Y(n_341)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_303),
.Y(n_586)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_307),
.A2(n_350),
.B1(n_403),
.B2(n_482),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_307),
.A2(n_603),
.B(n_607),
.Y(n_602)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_309),
.Y(n_608)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_311),
.Y(n_430)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_318),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2x1_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_500),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_434),
.B(n_496),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_331),
.B(n_658),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_375),
.B(n_377),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_332),
.B(n_375),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_332),
.B(n_375),
.Y(n_499)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.C(n_373),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_335),
.B1(n_373),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_360),
.C(n_366),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_340),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_353),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_341),
.B(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_360),
.B(n_366),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_369),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_373),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_378),
.B(n_381),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_429),
.C(n_431),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.C(n_397),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_383),
.A2(n_384),
.B1(n_387),
.B2(n_388),
.Y(n_441)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_397),
.A2(n_398),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_409),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_399),
.A2(n_409),
.B1(n_410),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_406),
.Y(n_649)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AOI32xp33_ASAP7_75t_SL g410 ( 
.A1(n_411),
.A2(n_414),
.A3(n_418),
.B1(n_422),
.B2(n_423),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_432),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_438),
.C(n_473),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_SL g658 ( 
.A1(n_436),
.A2(n_659),
.B(n_660),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_438),
.Y(n_659)
);

MAJx2_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.C(n_444),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_439),
.B(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.Y(n_495)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_454),
.C(n_461),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_461),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_476),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_459),
.B(n_460),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_459),
.B(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_459),
.B(n_520),
.Y(n_584)
);

OAI21xp33_ASAP7_75t_SL g596 ( 
.A1(n_459),
.A2(n_584),
.B(n_597),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_459),
.B(n_644),
.Y(n_643)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_494),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_474),
.B(n_494),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_477),
.C(n_479),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_475),
.B(n_567),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_477),
.A2(n_479),
.B1(n_480),
.B2(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_477),
.Y(n_568)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_489),
.C(n_491),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_481),
.A2(n_489),
.B1(n_490),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_481),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_482),
.A2(n_534),
.B(n_537),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_488),
.Y(n_631)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XOR2x2_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_498),
.B(n_499),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_657),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_569),
.B(n_655),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_562),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_547),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_504),
.B(n_547),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_508),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_505),
.B(n_509),
.C(n_565),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_515),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_514),
.B(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_533),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_516),
.B(n_533),
.Y(n_548)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx2_ASAP7_75t_SL g518 ( 
.A(n_519),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_521),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx3_ASAP7_75t_SL g530 ( 
.A(n_531),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_535),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_537),
.A2(n_625),
.B(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_538),
.B(n_608),
.Y(n_607)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

MAJx2_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_549),
.C(n_556),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_548),
.B(n_619),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_550),
.B(n_556),
.Y(n_619)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_566),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_564),
.B(n_656),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

AOI211x1_ASAP7_75t_L g569 ( 
.A1(n_570),
.A2(n_620),
.B(n_652),
.C(n_654),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_571),
.A2(n_613),
.B(n_614),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_571),
.B(n_621),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_601),
.Y(n_571)
);

NOR2x1_ASAP7_75t_SL g613 ( 
.A(n_572),
.B(n_601),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_594),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_594),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_574),
.A2(n_583),
.B1(n_585),
.B2(n_587),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_579),
.Y(n_574)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_580),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_582),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_591),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_598),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

XNOR2x1_ASAP7_75t_L g601 ( 
.A(n_602),
.B(n_609),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_616),
.C(n_617),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_603),
.Y(n_632)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_611),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_610),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_611),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_615),
.B(n_618),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_615),
.B(n_618),
.Y(n_653)
);

AOI21xp33_ASAP7_75t_L g621 ( 
.A1(n_622),
.A2(n_634),
.B(n_651),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_633),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_623),
.B(n_633),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

BUFx2_ASAP7_75t_SL g628 ( 
.A(n_629),
.Y(n_628)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_635),
.A2(n_640),
.B(n_650),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_636),
.B(n_637),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_636),
.B(n_637),
.Y(n_650)
);

INVx8_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_641),
.B(n_642),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_643),
.B(n_648),
.Y(n_642)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_662),
.A2(n_663),
.B(n_664),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g664 ( 
.A(n_665),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_667),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_667),
.B(n_688),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_668),
.B(n_676),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_668),
.B(n_677),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_669),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_670),
.B(n_673),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_670),
.B(n_673),
.Y(n_684)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_677),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_677),
.B(n_683),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_679),
.B(n_682),
.C(n_685),
.Y(n_681)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_683),
.Y(n_688)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_684),
.Y(n_683)
);


endmodule