module fake_jpeg_4240_n_278 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_227;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_43),
.B(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_9),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_55),
.B(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_7),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_7),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_59),
.B(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_31),
.B(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_11),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_22),
.B1(n_25),
.B2(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_102),
.B1(n_20),
.B2(n_27),
.Y(n_118)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_78),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_76),
.B(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_25),
.B1(n_22),
.B2(n_33),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_84),
.B1(n_12),
.B2(n_3),
.Y(n_133)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_85),
.Y(n_128)
);

NAND2x1_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_19),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_20),
.B(n_41),
.C(n_27),
.D(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_29),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_83),
.A2(n_91),
.B1(n_106),
.B2(n_3),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_29),
.B1(n_40),
.B2(n_36),
.Y(n_84)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_32),
.B1(n_61),
.B2(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_107),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_53),
.A2(n_30),
.B1(n_13),
.B2(n_2),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_66),
.B1(n_61),
.B2(n_41),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_111),
.B1(n_118),
.B2(n_123),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_109),
.B(n_95),
.Y(n_158)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_134),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_138),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_64),
.B(n_63),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_68),
.B(n_75),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_27),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_24),
.B1(n_20),
.B2(n_2),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_24),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_88),
.C(n_73),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_69),
.A2(n_24),
.B1(n_1),
.B2(n_0),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_129),
.B1(n_130),
.B2(n_141),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_20),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_12),
.B1(n_3),
.B2(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_97),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_100),
.Y(n_142)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_78),
.A2(n_1),
.B1(n_6),
.B2(n_11),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_149),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_162),
.B(n_168),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_99),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_140),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_154),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_112),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_77),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_164),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_99),
.B1(n_103),
.B2(n_87),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_124),
.B1(n_135),
.B2(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_122),
.B(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_70),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_72),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_72),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_88),
.B1(n_73),
.B2(n_96),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_136),
.B1(n_127),
.B2(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_101),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_189),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_182),
.B(n_191),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_145),
.B1(n_163),
.B2(n_164),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_170),
.B1(n_155),
.B2(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_163),
.B1(n_148),
.B2(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_117),
.C(n_139),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_120),
.C(n_132),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_190),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_195),
.B1(n_163),
.B2(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_133),
.B1(n_109),
.B2(n_114),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_128),
.B1(n_124),
.B2(n_135),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_179),
.B1(n_176),
.B2(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_206),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_165),
.B(n_146),
.C(n_157),
.D(n_149),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_209),
.B(n_210),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_157),
.B1(n_155),
.B2(n_159),
.Y(n_210)
);

AOI221xp5_ASAP7_75t_SL g211 ( 
.A1(n_175),
.A2(n_156),
.B1(n_141),
.B2(n_160),
.C(n_89),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_104),
.B(n_120),
.C(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_177),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_147),
.B(n_16),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_177),
.B(n_176),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_134),
.C(n_137),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_169),
.C(n_101),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_199),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_235),
.A3(n_173),
.B1(n_206),
.B2(n_179),
.C1(n_211),
.C2(n_194),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_198),
.C(n_193),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_228),
.C(n_210),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_190),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_227),
.B1(n_200),
.B2(n_209),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_215),
.C(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_204),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_216),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_230),
.B(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_247),
.C(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_197),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_203),
.B1(n_202),
.B2(n_207),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_244),
.A2(n_246),
.B1(n_201),
.B2(n_233),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_201),
.B1(n_194),
.B2(n_192),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_207),
.B1(n_188),
.B2(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_208),
.C(n_188),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_219),
.C(n_189),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_220),
.B(n_213),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_231),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_238),
.C(n_247),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_254),
.C(n_191),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_252),
.B(n_255),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_256),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_228),
.C(n_224),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_197),
.B1(n_195),
.B2(n_184),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_240),
.B1(n_249),
.B2(n_217),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_243),
.B(n_240),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_262),
.C(n_250),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_154),
.C(n_150),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_250),
.C(n_253),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_271)
);

AOI31xp33_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_265),
.A3(n_262),
.B(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_263),
.A2(n_154),
.B1(n_89),
.B2(n_150),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_SL g272 ( 
.A1(n_267),
.A2(n_17),
.B(n_93),
.C(n_270),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_266),
.C(n_93),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_272),
.B(n_17),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_271),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_277),
.Y(n_278)
);


endmodule