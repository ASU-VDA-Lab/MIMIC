module real_aes_92_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_785, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_785;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g222 ( .A(n_0), .B(n_159), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_1), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_2), .B(n_135), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_3), .B(n_157), .Y(n_472) );
INVx1_ASAP7_75t_L g131 ( .A(n_4), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_5), .B(n_135), .Y(n_180) );
NAND2xp33_ASAP7_75t_SL g242 ( .A(n_6), .B(n_141), .Y(n_242) );
INVx1_ASAP7_75t_L g234 ( .A(n_7), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_8), .A2(n_57), .B1(n_770), .B2(n_771), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_8), .Y(n_770) );
CKINVDCx16_ASAP7_75t_R g780 ( .A(n_9), .Y(n_780) );
AND2x2_ASAP7_75t_L g178 ( .A(n_10), .B(n_164), .Y(n_178) );
AND2x2_ASAP7_75t_L g465 ( .A(n_11), .B(n_240), .Y(n_465) );
AND2x2_ASAP7_75t_L g474 ( .A(n_12), .B(n_121), .Y(n_474) );
INVx2_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_14), .B(n_157), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_15), .Y(n_108) );
AOI221x1_ASAP7_75t_L g237 ( .A1(n_16), .A2(n_143), .B1(n_238), .B2(n_240), .C(n_241), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_17), .B(n_135), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_18), .A2(n_69), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_18), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_19), .B(n_135), .Y(n_514) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_21), .A2(n_90), .B1(n_126), .B2(n_135), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_22), .A2(n_143), .B(n_182), .Y(n_181) );
AOI221xp5_ASAP7_75t_SL g211 ( .A1(n_23), .A2(n_37), .B1(n_135), .B2(n_143), .C(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_24), .B(n_159), .Y(n_183) );
OA21x2_ASAP7_75t_L g122 ( .A1(n_25), .A2(n_89), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g165 ( .A(n_25), .B(n_89), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_26), .B(n_157), .Y(n_206) );
INVxp67_ASAP7_75t_L g236 ( .A(n_27), .Y(n_236) );
AND2x2_ASAP7_75t_L g175 ( .A(n_28), .B(n_163), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_29), .A2(n_143), .B(n_221), .Y(n_220) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_30), .A2(n_240), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_31), .B(n_157), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_32), .A2(n_143), .B(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_33), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_34), .B(n_157), .Y(n_528) );
AND2x2_ASAP7_75t_L g133 ( .A(n_35), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g141 ( .A(n_35), .B(n_131), .Y(n_141) );
INVx1_ASAP7_75t_L g147 ( .A(n_35), .Y(n_147) );
OR2x6_ASAP7_75t_L g109 ( .A(n_36), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_38), .B(n_135), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g142 ( .A1(n_39), .A2(n_82), .B1(n_143), .B2(n_145), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_40), .B(n_157), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_41), .B(n_135), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_42), .B(n_159), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_43), .A2(n_143), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g225 ( .A(n_44), .B(n_163), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_45), .B(n_159), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_46), .B(n_163), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_47), .B(n_135), .Y(n_496) );
INVx1_ASAP7_75t_L g129 ( .A(n_48), .Y(n_129) );
INVx1_ASAP7_75t_L g138 ( .A(n_48), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_49), .B(n_157), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_50), .Y(n_782) );
AND2x2_ASAP7_75t_L g504 ( .A(n_51), .B(n_163), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_52), .B(n_135), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_53), .B(n_159), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_54), .B(n_159), .Y(n_527) );
AND2x2_ASAP7_75t_L g166 ( .A(n_55), .B(n_163), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_56), .B(n_135), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_57), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_58), .B(n_157), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_59), .B(n_135), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_60), .A2(n_143), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_61), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_62), .B(n_164), .Y(n_207) );
AND2x2_ASAP7_75t_L g520 ( .A(n_63), .B(n_164), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_64), .A2(n_143), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_65), .B(n_157), .Y(n_184) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_66), .B(n_121), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_67), .B(n_159), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_68), .B(n_159), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_69), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_70), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_71), .A2(n_92), .B1(n_143), .B2(n_145), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_72), .B(n_157), .Y(n_517) );
INVx1_ASAP7_75t_L g134 ( .A(n_73), .Y(n_134) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_74), .B(n_159), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_75), .A2(n_143), .B(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_76), .A2(n_143), .B(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_77), .A2(n_143), .B(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g530 ( .A(n_78), .B(n_164), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_79), .B(n_163), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_80), .A2(n_84), .B1(n_126), .B2(n_135), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_81), .B(n_135), .Y(n_161) );
INVx1_ASAP7_75t_L g112 ( .A(n_83), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_85), .B(n_159), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_86), .B(n_159), .Y(n_214) );
AND2x2_ASAP7_75t_L g486 ( .A(n_87), .B(n_121), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_88), .A2(n_143), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_91), .B(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_93), .A2(n_143), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_94), .B(n_157), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_95), .B(n_135), .Y(n_224) );
INVxp67_ASAP7_75t_L g239 ( .A(n_96), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_97), .B(n_157), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_98), .A2(n_143), .B(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g519 ( .A(n_99), .Y(n_519) );
BUFx2_ASAP7_75t_L g761 ( .A(n_100), .Y(n_761) );
INVx1_ASAP7_75t_SL g764 ( .A(n_100), .Y(n_764) );
AOI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_772), .B(n_781), .Y(n_101) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_762), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_750), .B(n_758), .Y(n_103) );
AOI221xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_739), .B1(n_742), .B2(n_743), .C(n_745), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_113), .B1(n_442), .B2(n_735), .Y(n_105) );
INVx3_ASAP7_75t_SL g744 ( .A(n_106), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OR2x6_ASAP7_75t_SL g737 ( .A(n_108), .B(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g749 ( .A(n_108), .B(n_109), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_108), .B(n_738), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_109), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AO22x1_ASAP7_75t_L g743 ( .A1(n_113), .A2(n_442), .B1(n_736), .B2(n_744), .Y(n_743) );
XNOR2x1_ASAP7_75t_L g768 ( .A(n_113), .B(n_769), .Y(n_768) );
AND3x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_313), .C(n_387), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_255), .C(n_286), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_188), .B(n_197), .C(n_226), .Y(n_115) );
AOI21x1_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_167), .B(n_186), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_117), .A2(n_289), .B1(n_295), .B2(n_298), .Y(n_288) );
AND2x2_ASAP7_75t_L g422 ( .A(n_117), .B(n_190), .Y(n_422) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_151), .Y(n_117) );
BUFx2_ASAP7_75t_L g193 ( .A(n_118), .Y(n_193) );
AND2x2_ASAP7_75t_L g281 ( .A(n_118), .B(n_152), .Y(n_281) );
AND2x2_ASAP7_75t_L g352 ( .A(n_118), .B(n_196), .Y(n_352) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_119), .Y(n_246) );
AOI21x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_150), .Y(n_119) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_121), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_121), .A2(n_514), .B(n_515), .Y(n_513) );
BUFx4f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g218 ( .A(n_122), .Y(n_218) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_123), .B(n_165), .Y(n_164) );
AND2x4_ASAP7_75t_L g185 ( .A(n_123), .B(n_165), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_142), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_126), .A2(n_145), .B1(n_233), .B2(n_235), .Y(n_232) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_132), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g144 ( .A(n_129), .B(n_131), .Y(n_144) );
AND2x4_ASAP7_75t_L g157 ( .A(n_129), .B(n_139), .Y(n_157) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_L g143 ( .A(n_133), .B(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g149 ( .A(n_134), .Y(n_149) );
AND2x6_ASAP7_75t_L g159 ( .A(n_134), .B(n_137), .Y(n_159) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_141), .Y(n_135) );
INVx1_ASAP7_75t_L g243 ( .A(n_136), .Y(n_243) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx5_ASAP7_75t_L g160 ( .A(n_141), .Y(n_160) );
AND2x4_ASAP7_75t_L g145 ( .A(n_144), .B(n_146), .Y(n_145) );
NOR2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g245 ( .A(n_151), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g187 ( .A(n_152), .B(n_177), .Y(n_187) );
OR2x2_ASAP7_75t_L g195 ( .A(n_152), .B(n_196), .Y(n_195) );
AND2x4_ASAP7_75t_L g250 ( .A(n_152), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g297 ( .A(n_152), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_152), .B(n_196), .Y(n_305) );
AND2x2_ASAP7_75t_L g342 ( .A(n_152), .B(n_246), .Y(n_342) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_152), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_152), .B(n_176), .Y(n_383) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_162), .B(n_166), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_161), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_160), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_159), .B(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_160), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_160), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_160), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_160), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_160), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_160), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_160), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_160), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_160), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_160), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_160), .A2(n_527), .B(n_528), .Y(n_526) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_162), .A2(n_169), .B(n_175), .Y(n_168) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_162), .A2(n_169), .B(n_175), .Y(n_196) );
AOI21x1_ASAP7_75t_L g467 ( .A1(n_162), .A2(n_468), .B(n_474), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_163), .Y(n_162) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_163), .A2(n_211), .B(n_215), .Y(n_210) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_163), .A2(n_453), .B(n_454), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_163), .A2(n_481), .B(n_482), .Y(n_480) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_167), .B(n_245), .Y(n_340) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_167), .Y(n_441) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_176), .Y(n_167) );
AND2x2_ASAP7_75t_L g186 ( .A(n_168), .B(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g266 ( .A(n_168), .B(n_177), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_168), .B(n_297), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_174), .Y(n_169) );
AND2x2_ASAP7_75t_L g333 ( .A(n_176), .B(n_250), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_176), .B(n_245), .Y(n_389) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g191 ( .A(n_177), .Y(n_191) );
AND2x2_ASAP7_75t_L g260 ( .A(n_177), .B(n_251), .Y(n_260) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_177), .Y(n_280) );
AND2x4_ASAP7_75t_L g287 ( .A(n_177), .B(n_196), .Y(n_287) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_177), .B(n_246), .Y(n_434) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_185), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_185), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_185), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_185), .B(n_239), .Y(n_238) );
NOR3xp33_ASAP7_75t_L g241 ( .A(n_185), .B(n_242), .C(n_243), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_185), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_185), .A2(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g413 ( .A(n_186), .Y(n_413) );
INVx1_ASAP7_75t_L g355 ( .A(n_187), .Y(n_355) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_192), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g277 ( .A(n_191), .B(n_195), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_191), .B(n_246), .Y(n_370) );
AND2x2_ASAP7_75t_L g372 ( .A(n_191), .B(n_194), .Y(n_372) );
AOI32xp33_ASAP7_75t_L g438 ( .A1(n_191), .A2(n_254), .A3(n_409), .B1(n_439), .B2(n_441), .Y(n_438) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AND2x2_ASAP7_75t_L g264 ( .A(n_193), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g382 ( .A(n_193), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g405 ( .A(n_193), .B(n_266), .Y(n_405) );
AND2x2_ASAP7_75t_L g432 ( .A(n_193), .B(n_333), .Y(n_432) );
AND2x2_ASAP7_75t_L g358 ( .A(n_194), .B(n_246), .Y(n_358) );
AND2x2_ASAP7_75t_L g433 ( .A(n_194), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
NOR2x1p5_ASAP7_75t_L g291 ( .A(n_199), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g309 ( .A(n_199), .Y(n_309) );
OR2x2_ASAP7_75t_L g337 ( .A(n_199), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_SL g254 ( .A(n_200), .B(n_231), .Y(n_254) );
AND2x4_ASAP7_75t_L g270 ( .A(n_200), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g273 ( .A(n_200), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g301 ( .A(n_200), .B(n_210), .Y(n_301) );
OR2x2_ASAP7_75t_L g326 ( .A(n_200), .B(n_275), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_200), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_200), .B(n_210), .Y(n_361) );
INVx2_ASAP7_75t_L g377 ( .A(n_200), .Y(n_377) );
AND2x2_ASAP7_75t_L g392 ( .A(n_200), .B(n_230), .Y(n_392) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_200), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_200), .Y(n_421) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_207), .Y(n_200) );
AND2x2_ASAP7_75t_L g285 ( .A(n_208), .B(n_270), .Y(n_285) );
AND2x2_ASAP7_75t_L g306 ( .A(n_208), .B(n_254), .Y(n_306) );
INVx1_ASAP7_75t_L g338 ( .A(n_208), .Y(n_338) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_216), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g229 ( .A(n_210), .Y(n_229) );
INVx2_ASAP7_75t_L g275 ( .A(n_210), .Y(n_275) );
BUFx3_ASAP7_75t_L g292 ( .A(n_210), .Y(n_292) );
AND2x2_ASAP7_75t_L g331 ( .A(n_210), .B(n_216), .Y(n_331) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_210), .Y(n_429) );
INVx2_ASAP7_75t_L g244 ( .A(n_216), .Y(n_244) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
INVx1_ASAP7_75t_L g269 ( .A(n_216), .Y(n_269) );
OR2x2_ASAP7_75t_L g274 ( .A(n_216), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g294 ( .A(n_216), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_216), .B(n_271), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_216), .B(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AOI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_217) );
INVx4_ASAP7_75t_L g240 ( .A(n_218), .Y(n_240) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_218), .A2(n_459), .B(n_465), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_245), .B(n_247), .Y(n_226) );
AND2x2_ASAP7_75t_SL g227 ( .A(n_228), .B(n_230), .Y(n_227) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_228), .Y(n_437) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_SL g263 ( .A(n_229), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_229), .B(n_269), .Y(n_311) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_229), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_230), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g316 ( .A(n_230), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g367 ( .A(n_230), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_230), .A2(n_372), .B1(n_373), .B2(n_378), .C(n_381), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_230), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_244), .Y(n_230) );
INVx3_ASAP7_75t_L g271 ( .A(n_231), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_231), .B(n_275), .Y(n_375) );
AND2x2_ASAP7_75t_L g404 ( .A(n_231), .B(n_377), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_231), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g231 ( .A(n_232), .B(n_237), .Y(n_231) );
INVx3_ASAP7_75t_L g523 ( .A(n_240), .Y(n_523) );
AND2x2_ASAP7_75t_L g312 ( .A(n_245), .B(n_287), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_245), .A2(n_265), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g249 ( .A(n_246), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g258 ( .A(n_246), .Y(n_258) );
OR2x2_ASAP7_75t_L g304 ( .A(n_246), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_246), .B(n_287), .Y(n_396) );
OR2x2_ASAP7_75t_L g428 ( .A(n_246), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g440 ( .A(n_246), .B(n_346), .Y(n_440) );
INVxp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
INVx2_ASAP7_75t_L g318 ( .A(n_249), .Y(n_318) );
INVx3_ASAP7_75t_SL g384 ( .A(n_250), .Y(n_384) );
INVxp67_ASAP7_75t_L g334 ( .A(n_252), .Y(n_334) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AOI322xp5_ASAP7_75t_L g256 ( .A1(n_254), .A2(n_257), .A3(n_261), .B1(n_264), .B2(n_267), .C1(n_272), .C2(n_276), .Y(n_256) );
INVx1_ASAP7_75t_SL g345 ( .A(n_254), .Y(n_345) );
AND2x4_ASAP7_75t_L g430 ( .A(n_254), .B(n_317), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_278), .Y(n_255) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR2x2_ASAP7_75t_L g283 ( .A(n_258), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g379 ( .A(n_258), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g407 ( .A(n_258), .B(n_260), .Y(n_407) );
AOI32xp33_ASAP7_75t_L g408 ( .A1(n_258), .A2(n_259), .A3(n_409), .B1(n_411), .B2(n_414), .Y(n_408) );
OR2x2_ASAP7_75t_L g412 ( .A(n_258), .B(n_305), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_259), .B(n_284), .C(n_369), .Y(n_368) );
OAI22xp33_ASAP7_75t_SL g388 ( .A1(n_259), .A2(n_325), .B1(n_389), .B2(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g391 ( .A(n_262), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_266), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OAI322xp33_ASAP7_75t_L g314 ( .A1(n_270), .A2(n_274), .A3(n_283), .B1(n_315), .B2(n_318), .C1(n_319), .C2(n_320), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_270), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_270), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g293 ( .A(n_271), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g325 ( .A(n_271), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_271), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g386 ( .A(n_274), .Y(n_386) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_275), .Y(n_317) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B(n_285), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_281), .B(n_329), .Y(n_328) );
AOI322xp5_ASAP7_75t_SL g423 ( .A1(n_281), .A2(n_287), .A3(n_404), .B1(n_422), .B2(n_424), .C1(n_427), .C2(n_430), .Y(n_423) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_302), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_287), .B(n_297), .Y(n_319) );
INVx2_ASAP7_75t_SL g329 ( .A(n_287), .Y(n_329) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_SL g354 ( .A(n_293), .Y(n_354) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g399 ( .A(n_300), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g353 ( .A(n_301), .B(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B1(n_307), .B2(n_312), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR4xp75_ASAP7_75t_L g313 ( .A(n_314), .B(n_327), .C(n_347), .D(n_363), .Y(n_313) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_325), .A2(n_402), .B1(n_405), .B2(n_406), .Y(n_401) );
OR2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g410 ( .A(n_326), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B1(n_332), .B2(n_334), .C(n_335), .Y(n_327) );
INVx2_ASAP7_75t_L g346 ( .A(n_331), .Y(n_346) );
AND2x2_ASAP7_75t_L g403 ( .A(n_331), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_339), .B1(n_341), .B2(n_343), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g398 ( .A(n_342), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_343), .A2(n_349), .B1(n_365), .B2(n_368), .Y(n_364) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_353), .B1(n_355), .B2(n_356), .C(n_785), .Y(n_347) );
AND2x2_ASAP7_75t_SL g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g415 ( .A(n_354), .B(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g400 ( .A(n_362), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_371), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_385), .Y(n_381) );
NOR3xp33_ASAP7_75t_SL g387 ( .A(n_388), .B(n_393), .C(n_417), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_408), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B(n_399), .C(n_401), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g409 ( .A(n_400), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_413), .Y(n_411) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NAND4xp25_ASAP7_75t_SL g417 ( .A(n_418), .B(n_423), .C(n_431), .D(n_438), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_433), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g442 ( .A(n_443), .B(n_660), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_596), .C(n_643), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_531), .C(n_549), .D(n_575), .Y(n_444) );
OAI21xp33_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_490), .B(n_491), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_475), .Y(n_446) );
INVx1_ASAP7_75t_L g711 ( .A(n_447), .Y(n_711) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_455), .Y(n_447) );
INVx2_ASAP7_75t_L g535 ( .A(n_448), .Y(n_535) );
AND2x2_ASAP7_75t_L g555 ( .A(n_448), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g657 ( .A(n_448), .B(n_477), .Y(n_657) );
AND2x2_ASAP7_75t_L g717 ( .A(n_448), .B(n_536), .Y(n_717) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_449), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g601 ( .A(n_450), .B(n_458), .Y(n_601) );
BUFx3_ASAP7_75t_L g611 ( .A(n_450), .Y(n_611) );
AND2x2_ASAP7_75t_L g674 ( .A(n_450), .B(n_675), .Y(n_674) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AND2x4_ASAP7_75t_L g489 ( .A(n_451), .B(n_452), .Y(n_489) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g720 ( .A(n_456), .Y(n_720) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
AND2x2_ASAP7_75t_L g488 ( .A(n_457), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g675 ( .A(n_457), .Y(n_675) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g490 ( .A(n_458), .B(n_479), .Y(n_490) );
AND2x2_ASAP7_75t_L g552 ( .A(n_458), .B(n_466), .Y(n_552) );
INVx2_ASAP7_75t_L g557 ( .A(n_458), .Y(n_557) );
AND2x2_ASAP7_75t_L g559 ( .A(n_458), .B(n_467), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
INVx1_ASAP7_75t_L g537 ( .A(n_466), .Y(n_537) );
INVx2_ASAP7_75t_L g541 ( .A(n_466), .Y(n_541) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_466), .B(n_479), .Y(n_572) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_466), .Y(n_604) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_467), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_488), .Y(n_475) );
AND2x2_ASAP7_75t_L g638 ( .A(n_476), .B(n_583), .Y(n_638) );
INVx2_ASAP7_75t_SL g726 ( .A(n_476), .Y(n_726) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_478), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g646 ( .A(n_478), .B(n_559), .Y(n_646) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g534 ( .A(n_479), .Y(n_534) );
AND2x4_ASAP7_75t_L g536 ( .A(n_479), .B(n_537), .Y(n_536) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_479), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g629 ( .A(n_479), .Y(n_629) );
AND2x2_ASAP7_75t_L g648 ( .A(n_479), .B(n_587), .Y(n_648) );
AND2x2_ASAP7_75t_L g679 ( .A(n_479), .B(n_588), .Y(n_679) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
AND2x2_ASAP7_75t_L g618 ( .A(n_488), .B(n_572), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_488), .B(n_629), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_488), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_728) );
AND2x2_ASAP7_75t_L g731 ( .A(n_488), .B(n_538), .Y(n_731) );
INVx3_ASAP7_75t_L g584 ( .A(n_489), .Y(n_584) );
AND2x2_ASAP7_75t_L g587 ( .A(n_489), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g603 ( .A(n_490), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g612 ( .A(n_490), .Y(n_612) );
AND2x4_ASAP7_75t_SL g491 ( .A(n_492), .B(n_501), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_492), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g663 ( .A(n_492), .B(n_664), .Y(n_663) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_492), .B(n_625), .C(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g733 ( .A(n_492), .B(n_627), .Y(n_733) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g548 ( .A(n_494), .B(n_512), .Y(n_548) );
INVx1_ASAP7_75t_L g565 ( .A(n_494), .Y(n_565) );
INVx2_ASAP7_75t_L g578 ( .A(n_494), .Y(n_578) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_494), .Y(n_593) );
AND2x2_ASAP7_75t_L g607 ( .A(n_494), .B(n_580), .Y(n_607) );
AND2x2_ASAP7_75t_L g686 ( .A(n_494), .B(n_503), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_501), .A2(n_550), .B1(n_553), .B2(n_560), .C(n_566), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_501), .A2(n_679), .B1(n_680), .B2(n_681), .C(n_682), .Y(n_678) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
INVx2_ASAP7_75t_L g620 ( .A(n_502), .Y(n_620) );
AND2x2_ASAP7_75t_L g680 ( .A(n_502), .B(n_564), .Y(n_680) );
AND2x2_ASAP7_75t_L g690 ( .A(n_502), .B(n_576), .Y(n_690) );
OR2x2_ASAP7_75t_L g730 ( .A(n_502), .B(n_614), .Y(n_730) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_SL g547 ( .A(n_503), .B(n_548), .Y(n_547) );
NAND2x1_ASAP7_75t_L g563 ( .A(n_503), .B(n_512), .Y(n_563) );
INVx4_ASAP7_75t_L g592 ( .A(n_503), .Y(n_592) );
OR2x2_ASAP7_75t_L g634 ( .A(n_503), .B(n_521), .Y(n_634) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AND2x2_ASAP7_75t_L g685 ( .A(n_511), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
INVx2_ASAP7_75t_SL g573 ( .A(n_512), .Y(n_573) );
NOR2x1_ASAP7_75t_SL g579 ( .A(n_512), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g594 ( .A(n_512), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g625 ( .A(n_512), .B(n_592), .Y(n_625) );
AND2x2_ASAP7_75t_L g632 ( .A(n_512), .B(n_578), .Y(n_632) );
BUFx2_ASAP7_75t_L g666 ( .A(n_512), .Y(n_666) );
AND2x2_ASAP7_75t_L g677 ( .A(n_512), .B(n_592), .Y(n_677) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_521), .Y(n_545) );
AND2x2_ASAP7_75t_L g564 ( .A(n_521), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g595 ( .A(n_521), .Y(n_595) );
AND2x2_ASAP7_75t_L g621 ( .A(n_521), .B(n_577), .Y(n_621) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_530), .Y(n_522) );
AO21x1_ASAP7_75t_SL g580 ( .A1(n_523), .A2(n_524), .B(n_530), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
OAI31xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_536), .A3(n_538), .B(n_542), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g640 ( .A(n_534), .Y(n_640) );
NOR2xp67_ASAP7_75t_L g550 ( .A(n_535), .B(n_551), .Y(n_550) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_535), .A2(n_624), .A3(n_631), .B1(n_635), .B2(n_636), .C1(n_638), .C2(n_639), .Y(n_630) );
AND2x2_ASAP7_75t_L g702 ( .A(n_535), .B(n_679), .Y(n_702) );
AOI221xp5_ASAP7_75t_SL g615 ( .A1(n_536), .A2(n_616), .B1(n_618), .B2(n_619), .C(n_622), .Y(n_615) );
INVx2_ASAP7_75t_L g635 ( .A(n_536), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_538), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_538), .B(n_631), .Y(n_734) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_584), .Y(n_609) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g588 ( .A(n_541), .B(n_557), .Y(n_588) );
AND2x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g659 ( .A(n_545), .Y(n_659) );
O2A1O1Ixp5_ASAP7_75t_L g650 ( .A1(n_546), .A2(n_651), .B(n_653), .C(n_655), .Y(n_650) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_547), .A2(n_683), .B1(n_684), .B2(n_687), .Y(n_682) );
OR2x2_ASAP7_75t_L g637 ( .A(n_548), .B(n_634), .Y(n_637) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_554), .B(n_558), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g570 ( .A(n_557), .Y(n_570) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_559), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g613 ( .A(n_563), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_563), .B(n_564), .Y(n_656) );
OR2x2_ASAP7_75t_L g658 ( .A(n_563), .B(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_563), .B(n_707), .Y(n_706) );
BUFx2_ASAP7_75t_L g574 ( .A(n_565), .Y(n_574) );
NOR4xp25_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .C(n_573), .D(n_574), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g694 ( .A(n_568), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g722 ( .A(n_568), .B(n_571), .Y(n_722) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g652 ( .A(n_570), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_571), .B(n_600), .Y(n_687) );
AOI321xp33_ASAP7_75t_L g689 ( .A1(n_571), .A2(n_690), .A3(n_691), .B1(n_692), .B2(n_694), .C(n_697), .Y(n_689) );
INVx2_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_572), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_572), .B(n_611), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_573), .B(n_595), .Y(n_700) );
OR2x2_ASAP7_75t_L g727 ( .A(n_574), .B(n_611), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_581), .B(n_585), .Y(n_575) );
AND2x2_ASAP7_75t_L g616 ( .A(n_576), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g642 ( .A(n_578), .B(n_580), .Y(n_642) );
INVx2_ASAP7_75t_L g627 ( .A(n_579), .Y(n_627) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_582), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g683 ( .A(n_583), .B(n_635), .Y(n_683) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g641 ( .A(n_584), .B(n_642), .Y(n_641) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_584), .B(n_720), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g670 ( .A(n_588), .Y(n_670) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
NOR2xp67_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_592), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g617 ( .A(n_592), .Y(n_617) );
BUFx2_ASAP7_75t_L g699 ( .A(n_592), .Y(n_699) );
INVxp67_ASAP7_75t_L g707 ( .A(n_595), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_615), .C(n_630), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_605), .B(n_608), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g628 ( .A(n_601), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g681 ( .A(n_602), .Y(n_681) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g696 ( .A(n_604), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_605), .A2(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_SL g614 ( .A(n_607), .Y(n_614) );
AND2x2_ASAP7_75t_L g676 ( .A(n_607), .B(n_677), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_613), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_609), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g645 ( .A(n_611), .Y(n_645) );
OR2x2_ASAP7_75t_L g693 ( .A(n_614), .B(n_625), .Y(n_693) );
NOR4xp25_ASAP7_75t_L g725 ( .A(n_617), .B(n_666), .C(n_726), .D(n_727), .Y(n_725) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
OR2x2_ASAP7_75t_L g626 ( .A(n_620), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_620), .B(n_642), .Y(n_724) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_626), .B(n_628), .Y(n_622) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g713 ( .A(n_625), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g721 ( .A(n_627), .Y(n_721) );
AND2x4_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVxp67_ASAP7_75t_L g649 ( .A(n_632), .Y(n_649) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g665 ( .A(n_634), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g668 ( .A(n_640), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g714 ( .A(n_642), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B(n_649), .C(n_650), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g704 ( .A(n_646), .Y(n_704) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g708 ( .A(n_651), .Y(n_708) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_688), .C(n_709), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_667), .B(n_671), .C(n_678), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_674), .B(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g710 ( .A1(n_674), .A2(n_711), .B(n_712), .C(n_715), .Y(n_710) );
BUFx2_ASAP7_75t_L g691 ( .A(n_675), .Y(n_691) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_701), .Y(n_688) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_698), .A2(n_704), .B1(n_705), .B2(n_708), .Y(n_703) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_710), .B(n_718), .C(n_728), .D(n_734), .Y(n_709) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_722), .B2(n_723), .C(n_725), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
CKINVDCx11_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g742 ( .A(n_739), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx3_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVxp33_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_751), .A2(n_766), .B(n_767), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_R g766 ( .A(n_757), .Y(n_766) );
BUFx2_ASAP7_75t_L g777 ( .A(n_757), .Y(n_777) );
BUFx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NOR2xp67_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_774), .Y(n_783) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_776), .B(n_778), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
endmodule