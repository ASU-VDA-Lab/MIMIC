module real_jpeg_8680_n_11 (n_5, n_4, n_8, n_0, n_245, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_245;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_0),
.A2(n_1),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_10),
.B1(n_17),
.B2(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_0),
.A2(n_8),
.B1(n_23),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_33),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_1),
.A2(n_18),
.B(n_21),
.C(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_18),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_2),
.B(n_189),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_4),
.A2(n_9),
.B(n_46),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_5),
.A2(n_23),
.B(n_38),
.C(n_39),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_5),
.B(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_6),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_6),
.A3(n_23),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_6),
.A2(n_44),
.B(n_47),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_6),
.B(n_47),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_8),
.B1(n_26),
.B2(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_9),
.B1(n_34),
.B2(n_41),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_34),
.B(n_47),
.C(n_114),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_6),
.A2(n_10),
.B1(n_17),
.B2(n_41),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_10),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_7),
.A2(n_8),
.B1(n_18),
.B2(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g33 ( 
.A(n_7),
.B(n_34),
.CON(n_33),
.SN(n_33)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_26),
.B1(n_45),
.B2(n_46),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_23),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_9),
.B(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_27),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_39),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_10),
.A2(n_17),
.B1(n_45),
.B2(n_46),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_57),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_56),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_28),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_15),
.B(n_28),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_19),
.B1(n_25),
.B2(n_27),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_16),
.A2(n_19),
.B1(n_27),
.B2(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_22),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_24),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_51),
.C(n_52),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_29),
.A2(n_30),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.C(n_43),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_31),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_31),
.B(n_71),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_31),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_31),
.A2(n_69),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_31),
.B(n_71),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_31),
.A2(n_69),
.B1(n_186),
.B2(n_187),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_31),
.A2(n_69),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_31),
.A2(n_187),
.B(n_203),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_31),
.A2(n_69),
.B1(n_224),
.B2(n_228),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_31),
.A2(n_69),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_34),
.B(n_44),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_34),
.B(n_81),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_35),
.A2(n_43),
.B1(n_216),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_40),
.B(n_41),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_43),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_43),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_50),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_48),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_44),
.A2(n_48),
.B1(n_68),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_44),
.A2(n_48),
.B1(n_50),
.B2(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_45),
.B(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_51),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_237),
.B(n_243),
.Y(n_57)
);

OAI321xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_211),
.A3(n_230),
.B1(n_235),
.B2(n_236),
.C(n_245),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_197),
.B(n_210),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_178),
.B(n_196),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_106),
.B(n_162),
.C(n_177),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_94),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_63),
.B(n_94),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_85),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_77),
.B2(n_78),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_65),
.B(n_78),
.C(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI211xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_69),
.B(n_70),
.C(n_76),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_75),
.B1(n_79),
.B2(n_84),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_75),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_67),
.A2(n_75),
.B1(n_113),
.B2(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_67),
.B(n_92),
.C(n_117),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_67),
.A2(n_75),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_67),
.B(n_145),
.C(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_75),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_67),
.B(n_79),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_67),
.B(n_168),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_69),
.B(n_216),
.C(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_69),
.B(n_228),
.C(n_229),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_71),
.A2(n_75),
.B(n_139),
.C(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_71),
.A2(n_72),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_92),
.C(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_72),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_72),
.B(n_206),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_74),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_76),
.A2(n_93),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_76),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_169),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_93),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_86),
.A2(n_87),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_86),
.A2(n_87),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_92),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_101),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_101),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_92),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_103),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_96),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_98),
.B1(n_134),
.B2(n_139),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_161),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_154),
.B(n_160),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_141),
.B(n_153),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_131),
.B(n_140),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_120),
.B(n_130),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_115),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_134),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_135),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_144),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_163),
.B(n_164),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_175),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_174),
.C(n_175),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_193),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_185),
.C(n_193),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_183),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_194),
.B(n_195),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_192),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_190),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_199),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_208),
.B2(n_209),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_205),
.C(n_209),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_213),
.C(n_220),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_222),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_221),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_233),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);


endmodule