module fake_jpeg_31447_n_199 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_50),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_22),
.B(n_27),
.C(n_30),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_27),
.B(n_22),
.C(n_33),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_31),
.B1(n_25),
.B2(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_75),
.B1(n_66),
.B2(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_70),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_31),
.B1(n_34),
.B2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_75),
.B1(n_48),
.B2(n_24),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_53),
.B1(n_49),
.B2(n_39),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_42),
.B(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_29),
.B(n_24),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_102),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_74),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_95),
.B(n_64),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_92),
.B1(n_60),
.B2(n_59),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_48),
.B1(n_34),
.B2(n_30),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_83),
.B1(n_81),
.B2(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_94),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_90),
.B1(n_113),
.B2(n_102),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_124),
.B1(n_129),
.B2(n_116),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_81),
.B(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_127),
.B1(n_131),
.B2(n_91),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_71),
.B1(n_80),
.B2(n_88),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_93),
.B1(n_99),
.B2(n_63),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_58),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_79),
.B1(n_57),
.B2(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_32),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_110),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_96),
.B1(n_55),
.B2(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_116),
.B1(n_109),
.B2(n_104),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_134),
.B1(n_140),
.B2(n_106),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_110),
.B1(n_104),
.B2(n_108),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_112),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_97),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_121),
.B(n_127),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_124),
.C(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_150),
.C(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_134),
.C(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_108),
.C(n_112),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_154),
.B1(n_142),
.B2(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_26),
.B1(n_55),
.B2(n_73),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_161),
.Y(n_173)
);

NOR4xp25_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_136),
.C(n_142),
.D(n_137),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_137),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_166),
.Y(n_168)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_141),
.C(n_57),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_156),
.C(n_146),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_57),
.C(n_8),
.Y(n_170)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_5),
.C(n_13),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_9),
.B(n_12),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_12),
.B1(n_15),
.B2(n_3),
.Y(n_180)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_167),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_170),
.C(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_185),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_168),
.C(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_178),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_190),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_193),
.B(n_194),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_188),
.B1(n_181),
.B2(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_195),
.B(n_0),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_2),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_4),
.Y(n_199)
);


endmodule