module fake_jpeg_29641_n_467 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_59),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_72),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_74),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g128 ( 
.A(n_65),
.Y(n_128)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_1),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_83),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_92),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_5),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_30),
.B(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_93),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_87),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_91),
.Y(n_140)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_41),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_47),
.B1(n_45),
.B2(n_32),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_99),
.A2(n_104),
.B1(n_105),
.B2(n_5),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_47),
.B1(n_18),
.B2(n_43),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_34),
.B1(n_44),
.B2(n_43),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_33),
.B1(n_40),
.B2(n_37),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_76),
.B1(n_70),
.B2(n_63),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_45),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_32),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_50),
.A2(n_71),
.B1(n_53),
.B2(n_56),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_73),
.B1(n_61),
.B2(n_51),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_87),
.A2(n_33),
.B1(n_44),
.B2(n_34),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_136),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_22),
.B1(n_31),
.B2(n_27),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_144),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_41),
.Y(n_158)
);

CKINVDCx12_ASAP7_75t_R g142 ( 
.A(n_67),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_79),
.B(n_31),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_37),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_27),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_150),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_153),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_101),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_154),
.B(n_166),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_156),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_161),
.B1(n_165),
.B2(n_173),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_116),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_97),
.A2(n_22),
.B1(n_89),
.B2(n_36),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_85),
.B1(n_82),
.B2(n_57),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_100),
.A2(n_28),
.B1(n_82),
.B2(n_57),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_187),
.B1(n_118),
.B2(n_146),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_116),
.A2(n_40),
.B1(n_37),
.B2(n_24),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_177),
.A2(n_181),
.B(n_131),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_85),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_105),
.B(n_40),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_104),
.A2(n_40),
.B1(n_37),
.B2(n_24),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_98),
.B(n_40),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_195),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_193),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_109),
.A2(n_28),
.B1(n_37),
.B2(n_24),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_120),
.B(n_24),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_143),
.A2(n_149),
.B1(n_110),
.B2(n_109),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_137),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_148),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_17),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_134),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_5),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_SL g196 ( 
.A(n_127),
.B(n_17),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_134),
.B(n_138),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_127),
.B1(n_147),
.B2(n_148),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_150),
.B(n_120),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_217),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_169),
.A2(n_149),
.B1(n_110),
.B2(n_111),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_173),
.B1(n_191),
.B2(n_174),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_118),
.B1(n_96),
.B2(n_146),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_215),
.A2(n_221),
.B(n_233),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_202),
.B1(n_220),
.B2(n_219),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_236),
.B1(n_181),
.B2(n_177),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_114),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_123),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_153),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_125),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_189),
.C(n_188),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_117),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_155),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_155),
.B1(n_179),
.B2(n_161),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_238),
.A2(n_254),
.B1(n_211),
.B2(n_218),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g290 ( 
.A1(n_239),
.A2(n_247),
.B1(n_226),
.B2(n_204),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_257),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_182),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_175),
.B1(n_158),
.B2(n_160),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_246),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_292)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_183),
.B(n_170),
.C(n_152),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_158),
.B1(n_159),
.B2(n_190),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_168),
.B1(n_192),
.B2(n_111),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_117),
.B1(n_103),
.B2(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_191),
.B(n_186),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_256),
.A2(n_260),
.B(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_258),
.B(n_259),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_205),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_214),
.A2(n_156),
.B(n_178),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_213),
.B(n_163),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_261),
.B(n_262),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_167),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_199),
.B(n_167),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_263),
.B(n_267),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_265),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_227),
.B(n_193),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_208),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_180),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_198),
.B(n_180),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_207),
.B(n_180),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_202),
.A2(n_103),
.B1(n_112),
.B2(n_164),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_270),
.A2(n_216),
.B1(n_235),
.B2(n_237),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_210),
.B(n_167),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_226),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_212),
.A2(n_171),
.B(n_134),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_125),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_218),
.C(n_210),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_275),
.B(n_200),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_277),
.A2(n_280),
.B1(n_288),
.B2(n_306),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_278),
.A2(n_295),
.B1(n_299),
.B2(n_303),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_270),
.B1(n_250),
.B2(n_246),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_281),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_225),
.B1(n_172),
.B2(n_206),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_235),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_289),
.A2(n_287),
.B(n_307),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_247),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_254),
.A2(n_172),
.B1(n_206),
.B2(n_204),
.Y(n_295)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_171),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_307),
.C(n_276),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_242),
.B(n_232),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_298),
.B(n_302),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_238),
.A2(n_206),
.B1(n_229),
.B2(n_193),
.Y(n_299)
);

AOI32xp33_ASAP7_75t_L g302 ( 
.A1(n_244),
.A2(n_234),
.A3(n_232),
.B1(n_231),
.B2(n_138),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_229),
.B1(n_231),
.B2(n_156),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_240),
.A2(n_259),
.B1(n_239),
.B2(n_242),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_200),
.C(n_229),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_256),
.B(n_260),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_308),
.A2(n_303),
.B(n_290),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_314),
.C(n_317),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_312),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_265),
.C(n_273),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_286),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_286),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_265),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_261),
.Y(n_318)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_264),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_326),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_292),
.A2(n_253),
.B1(n_243),
.B2(n_252),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_331),
.Y(n_341)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_274),
.Y(n_324)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_241),
.B1(n_244),
.B2(n_253),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_330),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_285),
.B(n_264),
.C(n_267),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_287),
.B(n_258),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_283),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_333),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_278),
.A2(n_268),
.B1(n_269),
.B2(n_248),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_285),
.A2(n_245),
.B1(n_266),
.B2(n_262),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_263),
.Y(n_332)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_247),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_334),
.B(n_336),
.Y(n_344)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_335),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_327),
.A2(n_289),
.B1(n_290),
.B2(n_305),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_343),
.A2(n_363),
.B1(n_330),
.B2(n_323),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_312),
.A2(n_290),
.B(n_296),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_345),
.A2(n_351),
.B(n_313),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_325),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_347),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_332),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_354),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_338),
.A2(n_284),
.B(n_294),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_318),
.B(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_294),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_295),
.B(n_299),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_359),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_279),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_311),
.B(n_284),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_360),
.B(n_335),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_316),
.A2(n_293),
.B1(n_138),
.B2(n_8),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_6),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_364),
.Y(n_372)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_324),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_310),
.C(n_320),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_368),
.C(n_369),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_334),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_349),
.C(n_344),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_326),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_376),
.C(n_379),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_371),
.A2(n_356),
.B1(n_346),
.B2(n_345),
.Y(n_404)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_374),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_385),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_314),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_348),
.B(n_336),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_382),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_317),
.C(n_329),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_331),
.C(n_309),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_389),
.C(n_364),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_386),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_355),
.A2(n_316),
.B1(n_309),
.B2(n_321),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_384),
.A2(n_387),
.B1(n_362),
.B2(n_342),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_350),
.B(n_313),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_343),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_358),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_17),
.C(n_9),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_381),
.A2(n_341),
.B(n_347),
.Y(n_392)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_397),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_390),
.B(n_362),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_395),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_341),
.B1(n_342),
.B2(n_352),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_373),
.Y(n_399)
);

INVx11_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_375),
.A2(n_341),
.B1(n_352),
.B2(n_353),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_406),
.C(n_407),
.Y(n_415)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_404),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g405 ( 
.A1(n_377),
.A2(n_360),
.B(n_359),
.Y(n_405)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_405),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_364),
.C(n_365),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_366),
.C(n_365),
.Y(n_407)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_408),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_369),
.Y(n_410)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_410),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_404),
.A2(n_385),
.B(n_380),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_411),
.A2(n_400),
.B(n_401),
.Y(n_424)
);

AOI322xp5_ASAP7_75t_SL g417 ( 
.A1(n_393),
.A2(n_387),
.A3(n_384),
.B1(n_379),
.B2(n_372),
.C1(n_376),
.C2(n_370),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_420),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_393),
.A2(n_372),
.B1(n_358),
.B2(n_357),
.Y(n_418)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

A2O1A1O1Ixp25_ASAP7_75t_L g423 ( 
.A1(n_392),
.A2(n_357),
.B(n_389),
.C(n_363),
.D(n_12),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_394),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_424),
.A2(n_412),
.B(n_10),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_419),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_425),
.B(n_427),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_416),
.A2(n_413),
.B(n_422),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_426),
.A2(n_432),
.B(n_415),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_407),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_428),
.B(n_418),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_398),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_433),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_416),
.A2(n_406),
.B(n_396),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_398),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_423),
.A2(n_397),
.B1(n_403),
.B2(n_396),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_414),
.B1(n_421),
.B2(n_412),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_17),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_435),
.Y(n_438)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_439),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_440),
.B(n_446),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_SL g441 ( 
.A(n_430),
.B(n_414),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g453 ( 
.A(n_441),
.B(n_445),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_444),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_428),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_433),
.B(n_7),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_431),
.B(n_10),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_447),
.B(n_11),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_437),
.A2(n_429),
.B1(n_436),
.B2(n_434),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_449),
.Y(n_456)
);

INVx6_ASAP7_75t_L g451 ( 
.A(n_445),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_451),
.A2(n_455),
.B(n_11),
.Y(n_459)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_454),
.A2(n_444),
.B(n_12),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_438),
.B(n_424),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_457),
.B(n_459),
.Y(n_461)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_452),
.A2(n_443),
.B(n_13),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_458),
.A2(n_460),
.B(n_14),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_11),
.B(n_13),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_462),
.B(n_463),
.Y(n_465)
);

AOI321xp33_ASAP7_75t_L g463 ( 
.A1(n_456),
.A2(n_453),
.A3(n_451),
.B1(n_448),
.B2(n_450),
.C(n_15),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_461),
.B(n_448),
.C(n_14),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_464),
.B(n_15),
.C(n_465),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_15),
.Y(n_467)
);


endmodule