module fake_jpeg_11265_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_4),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_67),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_75),
.Y(n_80)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_5),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_5),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_66),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_5),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_78),
.Y(n_85)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_74),
.Y(n_82)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_16),
.B1(n_28),
.B2(n_37),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_8),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_38),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_91),
.B(n_100),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_17),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_14),
.B(n_10),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_44),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_104),
.B1(n_116),
.B2(n_41),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_16),
.B1(n_18),
.B2(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_15),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_48),
.A2(n_63),
.B1(n_18),
.B2(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_20),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_49),
.B(n_20),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_128),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_130),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_47),
.A3(n_58),
.B1(n_52),
.B2(n_61),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_30),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_9),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_9),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_84),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_141),
.Y(n_169)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_10),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_132),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_49),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_157),
.C(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_54),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_11),
.B1(n_54),
.B2(n_105),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_156),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_92),
.A2(n_116),
.B1(n_87),
.B2(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_98),
.B1(n_81),
.B2(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_154),
.B1(n_147),
.B2(n_145),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_93),
.B1(n_80),
.B2(n_117),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_84),
.B(n_93),
.C(n_96),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_114),
.A3(n_144),
.B1(n_127),
.B2(n_134),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_83),
.A3(n_91),
.B1(n_82),
.B2(n_90),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_114),
.C(n_119),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_114),
.B(n_119),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_126),
.B(n_150),
.C(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_182),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_168),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_153),
.B1(n_130),
.B2(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_176),
.B1(n_165),
.B2(n_162),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_135),
.B1(n_147),
.B2(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_181),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_184),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_125),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_190),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_201),
.C(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_179),
.C(n_167),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_178),
.C(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_196),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_162),
.B1(n_182),
.B2(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_164),
.B1(n_203),
.B2(n_187),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_178),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_191),
.B1(n_198),
.B2(n_193),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_172),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_185),
.A2(n_176),
.B1(n_168),
.B2(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_169),
.B1(n_175),
.B2(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

AOI221xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_178),
.B1(n_163),
.B2(n_177),
.C(n_161),
.Y(n_208)
);

OAI221xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_189),
.B1(n_200),
.B2(n_186),
.C(n_187),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_197),
.C(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_212),
.B(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_163),
.B1(n_164),
.B2(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_206),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_191),
.B(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_227),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_229),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_187),
.C(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_205),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_215),
.B1(n_206),
.B2(n_214),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_233),
.A2(n_224),
.B1(n_230),
.B2(n_221),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_226),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_219),
.B(n_217),
.C(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_225),
.B1(n_224),
.B2(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_242),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_218),
.B1(n_217),
.B2(n_235),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_240),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_237),
.B1(n_234),
.B2(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_232),
.C(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_250),
.C(n_243),
.Y(n_251)
);

AOI31xp33_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_243),
.A3(n_210),
.B(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_249),
.A2(n_246),
.B(n_245),
.Y(n_252)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_252),
.A2(n_248),
.B(n_232),
.C(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_253),
.Y(n_256)
);


endmodule