module real_jpeg_32920_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_1),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_1),
.A2(n_52),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_1),
.A2(n_52),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_1),
.A2(n_52),
.B1(n_248),
.B2(n_251),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_2),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g401 ( 
.A(n_2),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_3),
.B(n_483),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_6),
.Y(n_199)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g135 ( 
.A1(n_7),
.A2(n_81),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_7),
.A2(n_81),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_7),
.A2(n_81),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_7),
.B(n_324),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_7),
.A2(n_340),
.A3(n_342),
.B1(n_344),
.B2(n_350),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_7),
.B(n_117),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_7),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_7),
.B(n_161),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_8),
.Y(n_355)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_50),
.B1(n_57),
.B2(n_60),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_10),
.A2(n_60),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_60),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_10),
.A2(n_60),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_12),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

AOI22x1_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_47),
.B1(n_73),
.B2(n_76),
.Y(n_72)
);

INVx2_ASAP7_75t_R g76 ( 
.A(n_13),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_76),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_13),
.A2(n_76),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_270),
.B(n_482),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_20),
.B(n_485),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_22),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_24),
.B(n_78),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_25),
.A2(n_34),
.B1(n_46),
.B2(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_25),
.A2(n_72),
.B(n_77),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_25),
.A2(n_34),
.B1(n_72),
.B2(n_232),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_25),
.A2(n_56),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_36),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_26),
.Y(n_324)
);

AO22x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_31),
.Y(n_297)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_32),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_33),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_33),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_33),
.Y(n_142)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_78),
.Y(n_77)
);

AOI22x1_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_50),
.A2(n_82),
.A3(n_291),
.B1(n_295),
.B2(n_298),
.Y(n_290)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_54),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_54),
.B(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_54),
.B(n_486),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_256),
.B(n_266),
.C(n_267),
.D(n_269),
.Y(n_61)
);

OAI21x1_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_238),
.B(n_255),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_205),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_64),
.B(n_205),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_171),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_149),
.B2(n_150),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_67),
.B(n_149),
.C(n_171),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_84),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_68),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_68),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_69),
.Y(n_287)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_70),
.B(n_208),
.C(n_284),
.Y(n_446)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g438 ( 
.A1(n_71),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_71),
.Y(n_441)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_76),
.A2(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_76),
.B(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_77),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g232 ( 
.A(n_78),
.Y(n_232)
);

OAI21x1_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_81),
.B(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_81),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_81),
.B(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_115),
.B2(n_148),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_85),
.B(n_148),
.C(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_86),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_86),
.B(n_229),
.C(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_107),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_87),
.B(n_222),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_99),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

NAND2x1p5_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_99),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_89)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_91),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_91),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_91),
.Y(n_391)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_94),
.Y(n_386)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_98),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_98),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_99),
.B(n_224),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_101),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_104),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_105),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_153),
.B1(n_159),
.B2(n_161),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_109),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22x1_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_119),
.B1(n_122),
.B2(n_126),
.Y(n_118)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_113),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_128),
.B(n_134),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_116),
.A2(n_128),
.B1(n_247),
.B2(n_253),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_R g261 ( 
.A(n_116),
.B(n_253),
.Y(n_261)
);

AOI21x1_ASAP7_75t_L g440 ( 
.A1(n_116),
.A2(n_163),
.B(n_253),
.Y(n_440)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_117),
.B(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_135),
.B(n_139),
.Y(n_210)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_139),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_145),
.Y(n_349)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_151),
.A2(n_152),
.B(n_162),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_162),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_161),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AO22x2_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_161),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_162),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_162),
.A2(n_321),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_162),
.B(n_229),
.C(n_429),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_L g444 ( 
.A1(n_162),
.A2(n_230),
.B1(n_231),
.B2(n_321),
.Y(n_444)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_182),
.B(n_203),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_236),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_181),
.B(n_182),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_173),
.B(n_181),
.Y(n_460)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_175),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_203),
.B1(n_204),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_182),
.A2(n_237),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_190),
.Y(n_306)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_190),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_191),
.B(n_313),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_200),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_193),
.A2(n_304),
.B1(n_310),
.B2(n_313),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_193),
.B(n_313),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_197),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_199),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_199),
.Y(n_394)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_233),
.C(n_234),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_207),
.B(n_233),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_229),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_208),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_208),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_208),
.A2(n_285),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

AOI22x1_ASAP7_75t_L g463 ( 
.A1(n_208),
.A2(n_230),
.B1(n_231),
.B2(n_285),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_211),
.B(n_463),
.Y(n_462)
);

NAND2x1_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_221),
.Y(n_211)
);

OAI22x1_ASAP7_75t_L g431 ( 
.A1(n_212),
.A2(n_337),
.B1(n_416),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_212),
.Y(n_432)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_215),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_216),
.A2(n_330),
.B(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_221),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_221),
.B(n_368),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_221),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_235),
.B(n_465),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_274),
.Y(n_273)
);

NOR2x1_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_254),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_254),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_241),
.C(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_250),
.Y(n_341)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_258),
.Y(n_487)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_262),
.CI(n_264),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_474),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_423),
.B(n_473),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_357),
.B(n_422),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_331),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_281),
.B(n_331),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_282),
.B(n_289),
.C(n_320),
.Y(n_448)
);

XNOR2x1_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_285),
.B(n_410),
.C(n_420),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g454 ( 
.A(n_287),
.B(n_455),
.C(n_456),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_287),
.B(n_455),
.C(n_456),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_320),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_303),
.B1(n_318),
.B2(n_319),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_290),
.B(n_319),
.Y(n_429)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_303),
.B(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_303),
.B(n_403),
.Y(n_404)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx4f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_319),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.C(n_325),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_325),
.B(n_372),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_325),
.B(n_372),
.Y(n_405)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_326),
.B(n_397),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_329),
.B(n_330),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_336),
.C(n_338),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_332),
.A2(n_333),
.B1(n_415),
.B2(n_418),
.Y(n_414)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_367),
.C(n_368),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_337),
.A2(n_338),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_356),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_339),
.B(n_356),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx4f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_413),
.B(n_421),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_369),
.B(n_412),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_366),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_366),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_363),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_373),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_363),
.B(n_435),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_363),
.B(n_435),
.Y(n_445)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_406),
.B(n_411),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_395),
.B(n_405),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_379),
.B1(n_387),
.B2(n_392),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_392),
.B(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_402),
.B(n_404),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

INVx8_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_409),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_419),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_419),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_415),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_451),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_447),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_442),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_442),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_427),
.B(n_471),
.C(n_472),
.Y(n_470)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_444),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_438),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_445),
.C(n_446),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_443),
.B(n_450),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_446),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_448),
.B(n_449),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_466),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_464),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_464),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.C(n_461),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_462),
.Y(n_469)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_470),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_481),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_477),
.B(n_479),
.C(n_480),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_484),
.Y(n_483)
);


endmodule