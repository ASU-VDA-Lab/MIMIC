module fake_jpeg_26398_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_38),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_27),
.C(n_16),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_20),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_44),
.B1(n_45),
.B2(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_22),
.B1(n_43),
.B2(n_23),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_97),
.B(n_56),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_75),
.Y(n_104)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_86),
.Y(n_125)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_74),
.A2(n_98),
.B1(n_100),
.B2(n_48),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_18),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_83),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_95),
.B1(n_45),
.B2(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_19),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_33),
.Y(n_118)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_41),
.B1(n_35),
.B2(n_37),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_23),
.B1(n_17),
.B2(n_31),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_35),
.A3(n_31),
.B1(n_41),
.B2(n_37),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_103),
.B(n_71),
.C(n_100),
.D(n_74),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_41),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_113),
.B1(n_98),
.B2(n_81),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_35),
.B(n_36),
.C(n_45),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_115),
.B1(n_120),
.B2(n_124),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

OA22x2_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_56),
.B1(n_48),
.B2(n_36),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_88),
.B1(n_86),
.B2(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_34),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_77),
.A2(n_60),
.B(n_19),
.C(n_28),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_66),
.A2(n_34),
.B(n_30),
.C(n_28),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_79),
.A2(n_25),
.B(n_29),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_73),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_139),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_118),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_125),
.C(n_115),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_147),
.C(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_143),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_111),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_32),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_145),
.B(n_150),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_81),
.B(n_97),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_91),
.C(n_37),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_16),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_80),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_154),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_18),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_80),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_99),
.B1(n_96),
.B2(n_90),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_28),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_93),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_99),
.B1(n_73),
.B2(n_87),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_126),
.B1(n_116),
.B2(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_33),
.B1(n_25),
.B2(n_29),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_33),
.B1(n_25),
.B2(n_29),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_102),
.B1(n_114),
.B2(n_106),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_164),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_185),
.B1(n_194),
.B2(n_131),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_126),
.B(n_116),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_166),
.A2(n_167),
.B(n_174),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_26),
.B(n_34),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_175),
.B(n_6),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_119),
.B1(n_127),
.B2(n_26),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_183),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_127),
.B(n_121),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_143),
.B1(n_160),
.B2(n_7),
.Y(n_210)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_134),
.A2(n_16),
.B1(n_18),
.B2(n_3),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_9),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_187),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_21),
.B(n_2),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_16),
.C(n_21),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_193),
.C(n_195),
.Y(n_196)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_145),
.A3(n_142),
.B1(n_135),
.B2(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_8),
.C(n_13),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_141),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_7),
.C(n_13),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_136),
.C(n_146),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_164),
.C(n_166),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_150),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_1),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_6),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_6),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_186),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_243),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_171),
.B(n_162),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_235),
.B(n_241),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_169),
.B(n_179),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_201),
.C(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_172),
.C(n_189),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_185),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_172),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_169),
.B(n_187),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_193),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_196),
.B(n_195),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_249),
.Y(n_282)
);

AOI31xp33_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_203),
.A3(n_185),
.B(n_196),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_252),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_238),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_183),
.B1(n_208),
.B2(n_198),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_226),
.B1(n_237),
.B2(n_229),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_223),
.B1(n_218),
.B2(n_197),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_218),
.B1(n_224),
.B2(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_199),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_230),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_205),
.B1(n_224),
.B2(n_185),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_213),
.C(n_207),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_236),
.C(n_243),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_213),
.C(n_215),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_235),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_272),
.B(n_254),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_227),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_279),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_246),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_263),
.B1(n_267),
.B2(n_265),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_237),
.B(n_232),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_251),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_184),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_225),
.C(n_232),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_266),
.C(n_264),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_295),
.C(n_297),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_262),
.B(n_244),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_289),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_292),
.B1(n_284),
.B2(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_263),
.C(n_267),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_291),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_244),
.B(n_251),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_212),
.B1(n_245),
.B2(n_191),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_277),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_174),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_270),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_272),
.B(n_298),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_15),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_289),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_274),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_15),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_282),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_306),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_273),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_276),
.B1(n_281),
.B2(n_274),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_11),
.C(n_10),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_276),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_314),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_11),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_316),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_301),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_309),
.B(n_300),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_311),
.C(n_9),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_314),
.C(n_307),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_319),
.Y(n_325)
);

AOI321xp33_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_318),
.A3(n_321),
.B1(n_9),
.B2(n_4),
.C(n_1),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_2),
.B(n_3),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_4),
.Y(n_329)
);


endmodule