module real_jpeg_16359_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

OAI32xp33_ASAP7_75t_L g17 ( 
.A1(n_0),
.A2(n_18),
.A3(n_21),
.B1(n_27),
.B2(n_31),
.Y(n_17)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_0),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_0),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_0),
.A2(n_30),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_88),
.B1(n_116),
.B2(n_120),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_2),
.A2(n_88),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_2),
.A2(n_88),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_4),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_5),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_6),
.Y(n_210)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_6),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_6),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_8),
.Y(n_113)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_9),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_9),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_215),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_192),
.B(n_214),
.Y(n_12)
);

OAI21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_142),
.B(n_191),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_124),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_15),
.B(n_124),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_58),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_16),
.B(n_91),
.C(n_122),
.Y(n_213)
);

XOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_36),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_17),
.B(n_36),
.Y(n_195)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_19),
.A2(n_102),
.B1(n_104),
.B2(n_106),
.Y(n_101)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_26),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_26),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_30),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_31),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_46),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_37),
.A2(n_128),
.B1(n_129),
.B2(n_136),
.Y(n_127)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_38),
.B(n_47),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_39),
.A2(n_93),
.B(n_97),
.Y(n_92)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_42),
.Y(n_132)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_50),
.A2(n_97),
.A3(n_146),
.B1(n_150),
.B2(n_154),
.Y(n_145)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_109)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_54),
.Y(n_174)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_91),
.B1(n_122),
.B2(n_123),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_59),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_59),
.A2(n_122),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_69),
.B1(n_76),
.B2(n_85),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_60),
.A2(n_69),
.B1(n_76),
.B2(n_85),
.Y(n_199)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_65),
.B(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_67),
.A2(n_206),
.B1(n_208),
.B2(n_210),
.Y(n_205)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

NAND2x1p5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

OA22x2_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_91),
.A2(n_123),
.B1(n_145),
.B2(n_188),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_100),
.B1(n_109),
.B2(n_115),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_100),
.B1(n_109),
.B2(n_115),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_92),
.Y(n_226)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_140),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_125),
.A2(n_126),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_125),
.B(n_195),
.C(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_180),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_127),
.A2(n_161),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_164),
.B(n_190),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_160),
.Y(n_143)
);

NOR2xp67_ASAP7_75t_SL g190 ( 
.A(n_144),
.B(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_185),
.B(n_189),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_179),
.B(n_184),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_186),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_175),
.B(n_199),
.C(n_203),
.Y(n_254)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21x1_ASAP7_75t_SL g223 ( 
.A1(n_183),
.A2(n_224),
.B(n_226),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_213),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_213),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_212),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_211),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_229),
.B1(n_237),
.B2(n_249),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_238),
.B(n_244),
.Y(n_237)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_276),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_219),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_253),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_267),
.B1(n_271),
.B2(n_272),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);


endmodule