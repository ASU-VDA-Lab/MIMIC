module fake_jpeg_1019_n_445 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_45),
.B(n_63),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_55),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_12),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_0),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_26),
.B(n_12),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_73),
.B(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_27),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_79),
.Y(n_127)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_0),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_16),
.Y(n_99)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_32),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g86 ( 
.A(n_42),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_108),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_99),
.B(n_120),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_23),
.B1(n_30),
.B2(n_36),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_45),
.B(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_110),
.B(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_25),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_46),
.A2(n_41),
.B1(n_25),
.B2(n_40),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_35),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_3),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_22),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_86),
.B(n_38),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_16),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_48),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_59),
.B1(n_72),
.B2(n_64),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_138),
.A2(n_140),
.B1(n_145),
.B2(n_149),
.Y(n_219)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_62),
.B1(n_53),
.B2(n_49),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g218 ( 
.A1(n_142),
.A2(n_137),
.B1(n_101),
.B2(n_103),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_57),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_19),
.B1(n_32),
.B2(n_39),
.Y(n_145)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_80),
.B1(n_40),
.B2(n_39),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_51),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_155),
.Y(n_189)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_32),
.B1(n_19),
.B2(n_36),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_38),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_156),
.B(n_164),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_95),
.A2(n_30),
.B1(n_28),
.B2(n_42),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_159),
.B1(n_168),
.B2(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_104),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_11),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_166),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_175),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_8),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_177),
.B1(n_89),
.B2(n_102),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_9),
.B1(n_10),
.B2(n_100),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_96),
.B(n_9),
.C(n_107),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_181),
.Y(n_186)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_119),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_107),
.B(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_90),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_185),
.B(n_207),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_164),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_122),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_123),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_212),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_152),
.A2(n_106),
.B1(n_90),
.B2(n_121),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_123),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_102),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_92),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_150),
.B(n_115),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_115),
.B1(n_101),
.B2(n_103),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_92),
.B1(n_101),
.B2(n_103),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_SL g252 ( 
.A1(n_220),
.A2(n_143),
.B(n_142),
.C(n_151),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_146),
.B(n_121),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_223),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_149),
.A2(n_168),
.B1(n_176),
.B2(n_142),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_222),
.A2(n_177),
.B1(n_154),
.B2(n_140),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_178),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_248),
.Y(n_283)
);

BUFx12_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_244),
.B1(n_253),
.B2(n_185),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_164),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_241),
.Y(n_264)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_156),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_142),
.B1(n_156),
.B2(n_172),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_192),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_245),
.B(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_173),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_257),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_158),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_250),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_217),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_205),
.A2(n_160),
.B1(n_144),
.B2(n_167),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_255),
.B(n_256),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_217),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_180),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_199),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_211),
.A2(n_143),
.B(n_182),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_259),
.A2(n_195),
.B(n_194),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_260),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_261),
.A2(n_262),
.B1(n_281),
.B2(n_290),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_219),
.B1(n_188),
.B2(n_218),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_227),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_289),
.Y(n_300)
);

NOR4xp25_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_184),
.C(n_212),
.D(n_214),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_267),
.A2(n_280),
.B(n_270),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_193),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_234),
.B(n_214),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_291),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_220),
.B1(n_211),
.B2(n_218),
.Y(n_281)
);

CKINVDCx12_ASAP7_75t_R g285 ( 
.A(n_232),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_214),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_242),
.C(n_236),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_231),
.B(n_199),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_235),
.A2(n_218),
.B1(n_191),
.B2(n_190),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_257),
.B(n_191),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_242),
.B(n_224),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_218),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_260),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_295),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_241),
.B(n_213),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_286),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_277),
.Y(n_347)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_235),
.B(n_239),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_322),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_239),
.B(n_259),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_301),
.B(n_316),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_229),
.B(n_247),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_238),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_317),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_313),
.C(n_320),
.Y(n_329)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_274),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_228),
.C(n_225),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_282),
.A2(n_229),
.B(n_252),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_262),
.A2(n_261),
.B1(n_293),
.B2(n_281),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_318),
.B1(n_276),
.B2(n_287),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_253),
.B(n_237),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_233),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_268),
.A2(n_252),
.B1(n_258),
.B2(n_240),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_252),
.B(n_243),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_265),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_182),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_266),
.B(n_213),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_264),
.B(n_203),
.Y(n_324)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_272),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_342),
.Y(n_357)
);

NOR2x1_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_323),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_287),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_328),
.B(n_343),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_311),
.B(n_279),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_336),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_297),
.B1(n_316),
.B2(n_319),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_349),
.B1(n_350),
.B2(n_318),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_272),
.C(n_279),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_339),
.B(n_340),
.C(n_321),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_284),
.C(n_274),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_284),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_288),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_351),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_315),
.B1(n_297),
.B2(n_317),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_277),
.B1(n_294),
.B2(n_278),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_278),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_151),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_303),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_350),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_360),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_354),
.A2(n_345),
.B1(n_314),
.B2(n_321),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_300),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_365),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_333),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_362),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_338),
.A2(n_307),
.B(n_301),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_361),
.B(n_363),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_333),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_341),
.Y(n_363)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_298),
.Y(n_365)
);

XOR2x1_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_338),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_367),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_299),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_299),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_368),
.B(n_369),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_303),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_373),
.C(n_339),
.Y(n_375)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_374),
.A2(n_348),
.B1(n_309),
.B2(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_375),
.B(n_380),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_364),
.A2(n_331),
.B(n_344),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_357),
.B(n_367),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_351),
.C(n_352),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g381 ( 
.A(n_366),
.B(n_302),
.CI(n_331),
.CON(n_381),
.SN(n_381)
);

OAI21xp33_ASAP7_75t_SL g398 ( 
.A1(n_381),
.A2(n_368),
.B(n_372),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_355),
.C(n_358),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_384),
.C(n_273),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_353),
.A2(n_344),
.B(n_349),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_383),
.A2(n_357),
.B(n_356),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_324),
.C(n_297),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_345),
.B1(n_322),
.B2(n_346),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_386),
.A2(n_306),
.B1(n_305),
.B2(n_273),
.Y(n_399)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_387),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_376),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_393),
.B(n_402),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_397),
.Y(n_409)
);

OAI321xp33_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_381),
.A3(n_388),
.B1(n_187),
.B2(n_198),
.C(n_153),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_369),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_401),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_399),
.A2(n_387),
.B1(n_392),
.B2(n_388),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_232),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_389),
.A2(n_162),
.B(n_187),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_403),
.A2(n_394),
.B(n_147),
.Y(n_413)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_203),
.Y(n_406)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_406),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_390),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_408),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_400),
.A2(n_377),
.B1(n_383),
.B2(n_378),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_400),
.A2(n_377),
.B1(n_385),
.B2(n_381),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_413),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_375),
.C(n_382),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_417),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_380),
.C(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_418),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_419),
.A2(n_92),
.B(n_137),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_395),
.C(n_401),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_420),
.B(n_423),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_399),
.C(n_161),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_426),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_148),
.C(n_137),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_427),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_428),
.A2(n_412),
.B1(n_121),
.B2(n_414),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_429),
.B(n_409),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_435),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_421),
.A2(n_410),
.B(n_418),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_432),
.A2(n_434),
.B(n_422),
.Y(n_439)
);

NAND2x1_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_409),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_433),
.B(n_425),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_439),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_436),
.A2(n_424),
.B1(n_427),
.B2(n_414),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_434),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_441),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_443),
.A2(n_437),
.B(n_436),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_430),
.Y(n_445)
);


endmodule