module fake_jpeg_30714_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_12),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_66),
.B1(n_60),
.B2(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_66),
.B1(n_60),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_71),
.B1(n_64),
.B2(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_68),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_65),
.Y(n_104)
);

NAND2x1_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_65),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_65),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_51),
.B1(n_72),
.B2(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_62),
.B1(n_54),
.B2(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_61),
.B1(n_69),
.B2(n_53),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_59),
.B1(n_56),
.B2(n_55),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_115),
.B(n_14),
.Y(n_137)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_114),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_21),
.B1(n_50),
.B2(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_96),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_0),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_5),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_98),
.C(n_95),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_112),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_92),
.A3(n_94),
.B1(n_39),
.B2(n_23),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_1),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_2),
.B(n_3),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_94),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_93),
.A3(n_96),
.B1(n_20),
.B2(n_27),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_129),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_2),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_5),
.B(n_6),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_135),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_9),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_137),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_48),
.B1(n_29),
.B2(n_31),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_46),
.B1(n_36),
.B2(n_38),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_11),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_34),
.B1(n_45),
.B2(n_44),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_15),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_149),
.B1(n_135),
.B2(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_153),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_158),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_122),
.C(n_118),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_122),
.C(n_119),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_127),
.C(n_133),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_140),
.B(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_167),
.A2(n_162),
.B1(n_165),
.B2(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_151),
.C(n_142),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_146),
.C(n_164),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_171),
.B(n_169),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_166),
.B(n_156),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_177),
.Y(n_178)
);


endmodule