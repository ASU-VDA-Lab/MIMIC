module fake_ibex_1613_n_169 (n_7, n_20, n_17, n_25, n_36, n_18, n_3, n_22, n_28, n_32, n_39, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_38, n_15, n_37, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_169);

input n_7;
input n_20;
input n_17;
input n_25;
input n_36;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_38;
input n_15;
input n_37;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_169;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_148;
wire n_76;
wire n_118;
wire n_67;
wire n_164;
wire n_124;
wire n_110;
wire n_47;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_127;
wire n_121;
wire n_109;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_62;
wire n_71;
wire n_153;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_134;
wire n_42;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_44;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_49;
wire n_40;
wire n_66;
wire n_74;
wire n_90;
wire n_58;
wire n_43;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_72;
wire n_166;
wire n_163;
wire n_114;
wire n_97;
wire n_102;
wire n_131;
wire n_123;
wire n_52;
wire n_99;
wire n_135;
wire n_105;
wire n_156;
wire n_126;
wire n_154;
wire n_111;
wire n_104;
wire n_41;
wire n_45;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_149;
wire n_50;
wire n_92;
wire n_144;
wire n_101;
wire n_113;
wire n_138;
wire n_96;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_158;
wire n_132;
wire n_157;
wire n_160;
wire n_56;
wire n_146;
wire n_91;
wire n_54;

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx8_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_10),
.B(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_0),
.B(n_16),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx8_ASAP7_75t_SL g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_3),
.A2(n_4),
.B1(n_12),
.B2(n_21),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_3),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_57),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_60),
.C(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2x1p5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_51),
.Y(n_92)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

NOR2x1p5_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_72),
.Y(n_99)
);

OR2x6_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_66),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_59),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_75),
.C(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_76),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_70),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_76),
.B(n_73),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_73),
.B1(n_101),
.B2(n_107),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_73),
.B(n_97),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_90),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_83),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_94),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_105),
.B(n_102),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_99),
.B(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_103),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_96),
.B(n_97),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_79),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_82),
.A2(n_96),
.B(n_97),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_80),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_92),
.B(n_89),
.C(n_90),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_131),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_110),
.B1(n_125),
.B2(n_124),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_111),
.B1(n_129),
.B2(n_126),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_114),
.B1(n_121),
.B2(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_109),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_116),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_132),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_122),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_123),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_142),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_136),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_156),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_141),
.C(n_144),
.Y(n_163)
);

AOI222xp33_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_152),
.B1(n_154),
.B2(n_157),
.C1(n_160),
.C2(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_161),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_154),
.B1(n_161),
.B2(n_159),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_166),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_159),
.B(n_158),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_150),
.B1(n_158),
.B2(n_155),
.C(n_149),
.Y(n_169)
);


endmodule