module fake_jpeg_6927_n_233 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_17),
.Y(n_27)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_30),
.Y(n_50)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_42),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_45),
.B1(n_14),
.B2(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_14),
.B1(n_16),
.B2(n_22),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_14),
.B1(n_40),
.B2(n_33),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_85),
.B1(n_88),
.B2(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_86),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_33),
.B1(n_30),
.B2(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_28),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_30),
.B1(n_46),
.B2(n_29),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_51),
.C(n_55),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_106),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_72),
.B1(n_88),
.B2(n_85),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_51),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_54),
.B1(n_46),
.B2(n_27),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_70),
.B1(n_71),
.B2(n_87),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_44),
.B1(n_49),
.B2(n_20),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_13),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_122),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_119),
.B1(n_95),
.B2(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_124),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_81),
.B1(n_82),
.B2(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_99),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_69),
.B1(n_84),
.B2(n_44),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_44),
.B(n_43),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_43),
.B(n_48),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_25),
.B(n_1),
.C(n_2),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_89),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_133),
.B(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_135),
.B1(n_137),
.B2(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_102),
.B1(n_95),
.B2(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_84),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_134),
.C(n_120),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_31),
.B(n_28),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_90),
.C(n_49),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_91),
.B1(n_77),
.B2(n_49),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_48),
.B1(n_43),
.B2(n_22),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_19),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_23),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_125),
.Y(n_157)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_25),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_126),
.Y(n_161)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_159),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_108),
.B1(n_125),
.B2(n_126),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_153),
.A2(n_129),
.B1(n_137),
.B2(n_130),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_126),
.C(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_131),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_158),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_31),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_31),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_144),
.B(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_177),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_127),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_174),
.B1(n_153),
.B2(n_149),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_165),
.B1(n_159),
.B2(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_127),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_128),
.B1(n_20),
.B2(n_15),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_15),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_20),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_180),
.Y(n_195)
);

BUFx12f_ASAP7_75t_SL g187 ( 
.A(n_168),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_166),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_164),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.C(n_178),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_148),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_197),
.C(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_171),
.B1(n_170),
.B2(n_173),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_183),
.B1(n_190),
.B2(n_182),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_193),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_172),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_6),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_9),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_24),
.C(n_1),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_0),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_208),
.B(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_5),
.C(n_12),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_210),
.B(n_4),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_0),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_24),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_5),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_6),
.B(n_12),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_197),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_217),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_212),
.B(n_24),
.Y(n_223)
);

AOI21x1_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_5),
.B(n_11),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_223),
.A2(n_4),
.B(n_2),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_4),
.B(n_11),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_224),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_1),
.C(n_2),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_228),
.B(n_2),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_1),
.B(n_3),
.Y(n_232)
);

OAI21x1_ASAP7_75t_SL g233 ( 
.A1(n_232),
.A2(n_3),
.B(n_187),
.Y(n_233)
);


endmodule