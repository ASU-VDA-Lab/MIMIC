module fake_ibex_281_n_7430 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_974, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_854, n_1008, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_7430);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_974;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_7430;

wire n_4557;
wire n_6873;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_7170;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_7029;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_7042;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_7262;
wire n_6616;
wire n_6848;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_7063;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_6744;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_7147;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_7067;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_6842;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_6760;
wire n_7396;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_7082;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_7313;
wire n_7305;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_7332;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_7151;
wire n_2839;
wire n_7013;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_1070;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_6602;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_7397;
wire n_3979;
wire n_7324;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_7105;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_7187;
wire n_4854;
wire n_6732;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_7229;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_7099;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_7251;
wire n_7189;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_6868;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_6724;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_7097;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_7241;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_7264;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_7372;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_6926;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_7358;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_6878;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_7316;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_7207;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_7112;
wire n_7083;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_7026;
wire n_3572;
wire n_6114;
wire n_6996;
wire n_1121;
wire n_4823;
wire n_7366;
wire n_5195;
wire n_5541;
wire n_7033;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_7103;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_6864;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_1042;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_6941;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_6824;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_7169;
wire n_4225;
wire n_7140;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_6912;
wire n_3455;
wire n_6940;
wire n_1591;
wire n_7048;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_7303;
wire n_1409;
wire n_3524;
wire n_2744;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_7192;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_6802;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_7394;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_6855;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_7003;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_7161;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_6958;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_7226;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6711;
wire n_6124;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_7356;
wire n_5199;
wire n_7377;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_7315;
wire n_7360;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_7081;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_7224;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_7131;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_7155;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6971;
wire n_6128;
wire n_2361;
wire n_6804;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_7338;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_7221;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_6714;
wire n_4114;
wire n_6983;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_6857;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_6859;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_7101;
wire n_2954;
wire n_6379;
wire n_6911;
wire n_6766;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_7173;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6893;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_7349;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6850;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_6827;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_7068;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_6699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_6901;
wire n_4115;
wire n_3460;
wire n_2905;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3477;
wire n_3070;
wire n_1575;
wire n_6773;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6765;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_7391;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_7283;
wire n_2884;
wire n_3383;
wire n_7148;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_6704;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_7254;
wire n_2654;
wire n_7199;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_6939;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_6727;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_6883;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_6950;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_7327;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6915;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_7025;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_6922;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6731;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_7090;
wire n_1857;
wire n_1997;
wire n_7174;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_7250;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_6902;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_6837;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_6767;
wire n_7102;
wire n_4858;
wire n_6733;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_6723;
wire n_3339;
wire n_7177;
wire n_6900;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_7233;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_7031;
wire n_1517;
wire n_5973;
wire n_7012;
wire n_7238;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_7030;
wire n_7110;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_6856;
wire n_5770;
wire n_1763;
wire n_6976;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_7121;
wire n_1348;
wire n_7317;
wire n_1191;
wire n_4099;
wire n_7190;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_7429;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_6777;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_7390;
wire n_2410;
wire n_7145;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_6185;
wire n_6706;
wire n_5342;
wire n_6884;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_6745;
wire n_7210;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_1072;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_7191;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_6881;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_7136;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_7213;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_7034;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_6990;
wire n_3650;
wire n_6948;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_6816;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_6712;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_7098;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_7323;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_7149;
wire n_7219;
wire n_4919;
wire n_7320;
wire n_7175;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_1047;
wire n_1878;
wire n_4803;
wire n_1374;
wire n_7357;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_7218;
wire n_6863;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_7292;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_7142;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_7428;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_6805;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_7133;
wire n_2641;
wire n_7306;
wire n_1077;
wire n_7202;
wire n_6771;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_6695;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_7138;
wire n_7370;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_6978;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_6910;
wire n_2394;
wire n_1572;
wire n_7236;
wire n_1245;
wire n_4867;
wire n_7387;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_7122;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6925;
wire n_7024;
wire n_6483;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_6800;
wire n_7410;
wire n_5186;
wire n_7257;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6944;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_6980;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_7282;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_7334;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_7346;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4962;
wire n_1082;
wire n_5397;
wire n_4797;
wire n_2596;
wire n_1488;
wire n_7401;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_7245;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_6946;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_6897;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_7075;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6847;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_7367;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_6737;
wire n_3005;
wire n_4627;
wire n_6936;
wire n_5107;
wire n_6780;
wire n_4309;
wire n_4027;
wire n_7132;
wire n_6758;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_7419;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_7201;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_7265;
wire n_7232;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_1033;
wire n_7023;
wire n_3675;
wire n_7227;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_7273;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_6909;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_7070;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_6989;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_7046;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_7194;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_7290;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_7146;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_6960;
wire n_1226;
wire n_7253;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2682;
wire n_1666;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_6823;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_7414;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_6725;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_7184;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_6914;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_7152;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_6927;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_6916;
wire n_6973;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_7114;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_7354;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_6808;
wire n_7037;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_6747;
wire n_7335;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_6787;
wire n_1970;
wire n_3946;
wire n_7183;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_6784;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_6741;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_5319;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_6807;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_6795;
wire n_6898;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_6785;
wire n_7384;
wire n_6738;
wire n_3030;
wire n_5631;
wire n_6818;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_7393;
wire n_4517;
wire n_6021;
wire n_4511;
wire n_3210;
wire n_3221;
wire n_6966;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_6899;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_6754;
wire n_4067;
wire n_6822;
wire n_6796;
wire n_6849;
wire n_6836;
wire n_4997;
wire n_5906;
wire n_7355;
wire n_6755;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_7084;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_6717;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_6988;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_7256;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_7172;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_7117;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_6790;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_6840;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_7287;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_6748;
wire n_3788;
wire n_3448;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_7301;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_7156;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_6993;
wire n_2390;
wire n_7203;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_1053;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_7408;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_7307;
wire n_2787;
wire n_4540;
wire n_6987;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_7409;
wire n_7087;
wire n_3503;
wire n_2441;
wire n_7280;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_7107;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_6984;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6701;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_7288;
wire n_7248;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_6907;
wire n_4554;
wire n_1260;
wire n_7038;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_6730;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_7153;
wire n_5194;
wire n_7230;
wire n_4579;
wire n_5628;
wire n_6994;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_7308;
wire n_1775;
wire n_6889;
wire n_6361;
wire n_6803;
wire n_2570;
wire n_4025;
wire n_6751;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_7403;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_7369;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_6696;
wire n_2395;
wire n_7089;
wire n_6062;
wire n_4059;
wire n_7258;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_6943;
wire n_1832;
wire n_1128;
wire n_3718;
wire n_2376;
wire n_3398;
wire n_4878;
wire n_6252;
wire n_7080;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_7002;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_6726;
wire n_3238;
wire n_6740;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_6799;
wire n_2463;
wire n_6932;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_7008;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_7049;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_7062;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_6716;
wire n_6797;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_7215;
wire n_7340;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_7154;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_6965;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_7279;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_6846;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_7052;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_6931;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_6700;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_6853;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_7158;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_7299;
wire n_1830;
wire n_6770;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_7095;
wire n_1662;
wire n_7426;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_7076;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_7246;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_6951;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_6949;
wire n_5096;
wire n_6480;
wire n_7380;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_7167;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_6819;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_6937;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_6860;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_6833;
wire n_2159;
wire n_6865;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_7135;
wire n_6794;
wire n_3637;
wire n_7216;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_5900;
wire n_7421;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_7399;
wire n_1956;
wire n_7186;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_6498;
wire n_6720;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_6854;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_7197;
wire n_7015;
wire n_4408;
wire n_1175;
wire n_6832;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_7066;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_6779;
wire n_2567;
wire n_5645;
wire n_7044;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_7329;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_6887;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_6769;
wire n_6903;
wire n_2433;
wire n_7255;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_6861;
wire n_2130;
wire n_4862;
wire n_7270;
wire n_5114;
wire n_7071;
wire n_6697;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_6826;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_7235;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_7129;
wire n_4242;
wire n_7243;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_7342;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_7310;
wire n_2911;
wire n_1828;
wire n_6972;
wire n_1389;
wire n_6380;
wire n_7200;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_6703;
wire n_7116;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6719;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_7208;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_7337;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_7055;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_7073;
wire n_2637;
wire n_7417;
wire n_7159;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_7314;
wire n_3791;
wire n_6904;
wire n_6778;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_7294;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_7016;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_6444;
wire n_7422;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_6749;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_6985;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_7178;
wire n_7330;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_7388;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6692;
wire n_7079;
wire n_6590;
wire n_3036;
wire n_7209;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_7206;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_6702;
wire n_3046;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_7051;
wire n_7278;
wire n_2791;
wire n_1450;
wire n_7416;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_7274;
wire n_1442;
wire n_2168;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_6820;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_6952;
wire n_3261;
wire n_5324;
wire n_6547;
wire n_7065;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_6995;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_7326;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_7423;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_6879;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_7104;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_7106;
wire n_3615;
wire n_7198;
wire n_7381;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_7182;
wire n_6310;
wire n_6852;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_6961;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_7126;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_6956;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_6643;
wire n_6569;
wire n_6814;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_7176;
wire n_4159;
wire n_7056;
wire n_4372;
wire n_5528;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_7368;
wire n_5464;
wire n_6895;
wire n_6548;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_6890;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_6789;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_6867;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_6764;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_6935;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_7382;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_7130;
wire n_6942;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6772;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_6955;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_7427;
wire n_6908;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_6874;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_6736;
wire n_4259;
wire n_1620;
wire n_7376;
wire n_5196;
wire n_5086;
wire n_7018;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_7134;
wire n_3967;
wire n_2373;
wire n_2275;
wire n_1853;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_7348;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_7383;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_7053;
wire n_5483;
wire n_6713;
wire n_6919;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_7240;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_6750;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_6981;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_6828;
wire n_5123;
wire n_6160;
wire n_7043;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_7074;
wire n_7119;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_6875;
wire n_1701;
wire n_5236;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_6870;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_6715;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_7386;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_7007;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_7027;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_7009;
wire n_6140;
wire n_5903;
wire n_7263;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_6663;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_6844;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_6999;
wire n_4571;
wire n_7214;
wire n_6982;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_6843;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_6877;
wire n_2821;
wire n_6892;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_7162;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_7268;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_7398;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_7304;
wire n_7036;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_2490;
wire n_3127;
wire n_7171;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_2300;
wire n_1120;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_5152;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_7293;
wire n_1264;
wire n_6752;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_7363;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_6698;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6977;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_7028;
wire n_1628;
wire n_6810;
wire n_1773;
wire n_7237;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_7039;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_6791;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_6967;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_6768;
wire n_2458;
wire n_7144;
wire n_3032;
wire n_3401;
wire n_7362;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_6947;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6938;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_6906;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_7124;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_6918;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_7143;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_6834;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_6812;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_7123;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_7072;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_6762;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_6992;
wire n_7109;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_7325;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_6759;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_7137;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_7350;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_7311;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_7244;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_7339;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_7247;
wire n_2346;
wire n_4695;
wire n_7331;
wire n_7128;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_7284;
wire n_4163;
wire n_7321;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_7309;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_7163;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_6886;
wire n_4832;
wire n_5229;
wire n_7054;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_2555;
wire n_1587;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_6959;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_7413;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_7185;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_6710;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_6945;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_6776;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_7336;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_6905;
wire n_7120;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_7374;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_6964;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_7001;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_7111;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_6798;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_7165;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_6888;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_7389;
wire n_1501;
wire n_7418;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_7375;
wire n_7096;
wire n_5257;
wire n_7281;
wire n_7300;
wire n_4397;
wire n_6920;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_6781;
wire n_4229;
wire n_4294;
wire n_7085;
wire n_1919;
wire n_4351;
wire n_6811;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_6921;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_7212;
wire n_7285;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_7032;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_7125;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_7160;
wire n_7100;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_7319;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_6722;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_7371;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_7361;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_7010;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_7289;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_7004;
wire n_7021;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_7234;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_6975;
wire n_7266;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6573;
wire n_6786;
wire n_6774;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_6851;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_7211;
wire n_4335;
wire n_7141;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_6729;
wire n_7150;
wire n_6882;
wire n_1168;
wire n_5500;
wire n_7378;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_7420;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_6998;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_6721;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_7271;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_7322;
wire n_7022;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_6885;
wire n_7217;
wire n_7166;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_6806;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_6933;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_7297;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_7179;
wire n_5984;
wire n_6385;
wire n_7415;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_7057;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_6793;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_6746;
wire n_4702;
wire n_1341;
wire n_7411;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_7108;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_7220;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_7223;
wire n_2544;
wire n_7261;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_7092;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_6728;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_7275;
wire n_3768;
wire n_4224;
wire n_7272;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_7249;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_7168;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_7091;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_6858;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_7228;
wire n_3272;
wire n_7353;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_6841;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_6896;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_6954;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_7000;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_7040;
wire n_6132;
wire n_7196;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6872;
wire n_6089;
wire n_5211;
wire n_7205;
wire n_1668;
wire n_7260;
wire n_5861;
wire n_7086;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_7047;
wire n_7412;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_7077;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6831;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6968;
wire n_6415;
wire n_2280;
wire n_1038;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_7402;
wire n_2876;
wire n_6670;
wire n_5321;
wire n_3301;
wire n_2370;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_7405;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_7343;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_6046;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_7252;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_6991;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_6705;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_7188;
wire n_6913;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_7113;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_6734;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_7296;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_6825;
wire n_1036;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_6743;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_7345;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_7157;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_6809;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_7115;
wire n_1884;
wire n_6632;
wire n_1589;
wire n_2717;
wire n_5720;
wire n_7286;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_5561;
wire n_4762;
wire n_1877;
wire n_6871;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_7344;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_6953;
wire n_3145;
wire n_5682;
wire n_6891;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1566;
wire n_1464;
wire n_7127;
wire n_6601;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6565;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_6979;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_7050;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_6930;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_7118;
wire n_7259;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_6821;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_6775;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6815;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_7069;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_7011;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_6763;
wire n_6782;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_6839;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_7164;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_7017;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_6761;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_6974;
wire n_1898;
wire n_1254;
wire n_7312;
wire n_6894;
wire n_2524;
wire n_3927;
wire n_7045;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_7277;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_6997;
wire n_3747;
wire n_1323;
wire n_6753;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_7359;
wire n_3632;
wire n_5200;
wire n_7225;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_7020;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_7392;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_6924;
wire n_5485;
wire n_5737;
wire n_6876;
wire n_7424;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_6962;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_7059;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_6970;
wire n_5185;
wire n_6829;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_6830;
wire n_3290;
wire n_7365;
wire n_3585;
wire n_7094;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_7035;
wire n_5306;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_6838;
wire n_2698;
wire n_6869;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_6735;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_6866;
wire n_4383;
wire n_7395;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_7005;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_6742;
wire n_3063;
wire n_4543;
wire n_6969;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_7180;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_6929;
wire n_2255;
wire n_1820;
wire n_6986;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_6709;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_7385;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_6756;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_6718;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_7078;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_7093;
wire n_1167;
wire n_7333;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_6757;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_6880;
wire n_3824;
wire n_7425;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_7302;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_6934;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_7019;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_7088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_7204;
wire n_7014;
wire n_1165;
wire n_6708;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_7341;
wire n_7407;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_6801;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_7193;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_7373;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_7291;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_6707;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_7239;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_6835;
wire n_7406;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_6792;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_6928;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_7242;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5627;
wire n_5542;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_7181;
wire n_1161;
wire n_1103;
wire n_6739;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_7139;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_7404;
wire n_2870;
wire n_6862;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_7328;
wire n_6783;
wire n_4738;
wire n_7231;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_7058;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_7041;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_6788;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_7364;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_7006;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_6817;
wire n_1661;
wire n_6261;
wire n_7276;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_7269;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_1039;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_6845;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_7222;
wire n_4595;
wire n_4418;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_7347;
wire n_4944;
wire n_7060;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_7064;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_6917;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_7400;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_6813;
wire n_2670;
wire n_7379;
wire n_1745;
wire n_7318;
wire n_7352;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_7295;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_7267;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_6963;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_6923;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_5393;
wire n_4782;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_7061;
wire n_7351;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_7298;
wire n_2497;
wire n_7195;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_6957;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_252),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_1017),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_955),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_784),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_318),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_836),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_929),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_1001),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_140),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1009),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_937),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_364),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_881),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_499),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_154),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_603),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_255),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_639),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_331),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_766),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_727),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_1004),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_863),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1011),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_1002),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_973),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_991),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1021),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_92),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_929),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_286),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_759),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_728),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_875),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_67),
.Y(n_1066)
);

CKINVDCx14_ASAP7_75t_R g1067 ( 
.A(n_710),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_640),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_855),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_529),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_752),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_737),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_72),
.Y(n_1073)
);

BUFx8_ASAP7_75t_SL g1074 ( 
.A(n_175),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_871),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_325),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_658),
.Y(n_1077)
);

BUFx10_ASAP7_75t_L g1078 ( 
.A(n_868),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_757),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_538),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_1019),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_997),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_388),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_712),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_211),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_105),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_872),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_821),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_854),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_363),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_998),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1026),
.Y(n_1092)
);

BUFx10_ASAP7_75t_L g1093 ( 
.A(n_424),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_86),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_847),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_850),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1002),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_450),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_193),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_486),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_660),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_1022),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_282),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_102),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_954),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_926),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_625),
.Y(n_1107)
);

BUFx2_ASAP7_75t_SL g1108 ( 
.A(n_559),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_841),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_219),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_484),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_646),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_622),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_518),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_105),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_764),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_401),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_844),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_468),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_195),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_778),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_674),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_861),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_932),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_437),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_342),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_827),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_132),
.Y(n_1128)
);

BUFx5_ASAP7_75t_L g1129 ( 
.A(n_576),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_921),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_887),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_493),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_112),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_404),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_482),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_911),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_220),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_466),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_67),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_157),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_601),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_788),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_338),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_447),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_547),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_304),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_695),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_542),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_993),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_639),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_414),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_820),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_234),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_121),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_676),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_722),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_242),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_33),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_643),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_129),
.Y(n_1161)
);

BUFx10_ASAP7_75t_L g1162 ( 
.A(n_463),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1014),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_853),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_567),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_571),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_989),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1016),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_285),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_213),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_720),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_271),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_787),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_441),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_790),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_196),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_378),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_219),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_546),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_287),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_432),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_848),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_668),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_920),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_140),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_60),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_983),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_31),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_886),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_140),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_276),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_854),
.Y(n_1192)
);

CKINVDCx14_ASAP7_75t_R g1193 ( 
.A(n_372),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_580),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_509),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_878),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_85),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_614),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_741),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_76),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_870),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_231),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_451),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_259),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_401),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_927),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_733),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_403),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_313),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_570),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_845),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_291),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_241),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1026),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_192),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_715),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_407),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_606),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_887),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_496),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_888),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_386),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_285),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_4),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_381),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_329),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_125),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_185),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_489),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_472),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_325),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_365),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_354),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_493),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_235),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_643),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_602),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_705),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_941),
.Y(n_1239)
);

CKINVDCx16_ASAP7_75t_R g1240 ( 
.A(n_774),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_767),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_31),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_885),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_166),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_350),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_541),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_536),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_382),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_761),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_978),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_262),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_681),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_410),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1014),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_880),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_681),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_208),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_484),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_470),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_126),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_928),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_942),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_182),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_873),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_590),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_846),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_145),
.Y(n_1267)
);

CKINVDCx16_ASAP7_75t_R g1268 ( 
.A(n_895),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_947),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_567),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_108),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_458),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_181),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_365),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_784),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_296),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_758),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_272),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_970),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_722),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_193),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_675),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_442),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_582),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_539),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_1015),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_114),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_232),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_135),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_321),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_27),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_624),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_997),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_549),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_842),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_643),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_332),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_899),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_982),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_620),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_306),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_340),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_815),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1012),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_190),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_869),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_561),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_205),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_21),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_203),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_377),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1027),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_37),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_118),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_281),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_984),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_630),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_366),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_619),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_132),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_640),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_570),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_560),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_745),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_434),
.Y(n_1325)
);

CKINVDCx16_ASAP7_75t_R g1326 ( 
.A(n_349),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_821),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_877),
.Y(n_1328)
);

CKINVDCx16_ASAP7_75t_R g1329 ( 
.A(n_832),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_711),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_160),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_147),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_206),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_825),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_182),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_863),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_15),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_214),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_904),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_962),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_838),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_615),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_973),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_266),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_916),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_701),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1018),
.Y(n_1347)
);

CKINVDCx14_ASAP7_75t_R g1348 ( 
.A(n_995),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_982),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_23),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_320),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_945),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_59),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_82),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_851),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_994),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_678),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_131),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_419),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_144),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_11),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_4),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_101),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_705),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_162),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_322),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_19),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_452),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_462),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_397),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_211),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_215),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_906),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_417),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_833),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_312),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_280),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1000),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_791),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_635),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1003),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_536),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_285),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_992),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_680),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_362),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_366),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_849),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_80),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_107),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_976),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_925),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_324),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_18),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_804),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_501),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_52),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_914),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_636),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1016),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_958),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_836),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_144),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_881),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_742),
.Y(n_1405)
);

BUFx2_ASAP7_75t_SL g1406 ( 
.A(n_514),
.Y(n_1406)
);

CKINVDCx16_ASAP7_75t_R g1407 ( 
.A(n_860),
.Y(n_1407)
);

BUFx5_ASAP7_75t_L g1408 ( 
.A(n_992),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_260),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_119),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_954),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_816),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_332),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_757),
.Y(n_1414)
);

BUFx10_ASAP7_75t_L g1415 ( 
.A(n_518),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_232),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_617),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_395),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_683),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_233),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_19),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_891),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1028),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_130),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_852),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_3),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_532),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_796),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_98),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_868),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_698),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_172),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_246),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_386),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_757),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_751),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_474),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_135),
.Y(n_1438)
);

CKINVDCx16_ASAP7_75t_R g1439 ( 
.A(n_15),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_857),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_879),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_892),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_132),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_286),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_270),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_19),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_631),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_208),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_874),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_13),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_791),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_377),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_57),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_256),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_872),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_356),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_980),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_374),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_68),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_486),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_245),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_546),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_316),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_925),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_105),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_302),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_495),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_536),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_656),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_977),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1010),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_365),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_942),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_834),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_332),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_740),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_286),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_647),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_683),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_678),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_251),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_603),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_722),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_441),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_145),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_638),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_887),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_104),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_377),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_193),
.Y(n_1490)
);

BUFx5_ASAP7_75t_L g1491 ( 
.A(n_560),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_123),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_324),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_215),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_701),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_875),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_866),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_962),
.Y(n_1498)
);

BUFx5_ASAP7_75t_L g1499 ( 
.A(n_171),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_673),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_745),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_760),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_845),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_791),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1007),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_884),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_984),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1030),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_945),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1028),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_795),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_497),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_68),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_763),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_745),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_981),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_856),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1025),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_988),
.Y(n_1519)
);

CKINVDCx14_ASAP7_75t_R g1520 ( 
.A(n_637),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_922),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_318),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_808),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_926),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_707),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_928),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_667),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_491),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_968),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_341),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_578),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_754),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1005),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_224),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_77),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_52),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_485),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1024),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_328),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_45),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_487),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_90),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_740),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_924),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_392),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_120),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_862),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_712),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_227),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_469),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1006),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_961),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_508),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1003),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_23),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_7),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_865),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_503),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_858),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_149),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_641),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_499),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_206),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_252),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_765),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_262),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_761),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_752),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_816),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_169),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_680),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_144),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_312),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_761),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_418),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_930),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1020),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_638),
.Y(n_1578)
);

BUFx5_ASAP7_75t_L g1579 ( 
.A(n_277),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_996),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_464),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_841),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_940),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_330),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_864),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_242),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_490),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_120),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_630),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_847),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1013),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_408),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_828),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_115),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_205),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_883),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_466),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_303),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_600),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_676),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_720),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_278),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_845),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_704),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_34),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_552),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_547),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_859),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_947),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_218),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_510),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_288),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_856),
.Y(n_1613)
);

BUFx8_ASAP7_75t_SL g1614 ( 
.A(n_409),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_662),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_372),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_990),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_730),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_391),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_683),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_80),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_235),
.Y(n_1622)
);

CKINVDCx16_ASAP7_75t_R g1623 ( 
.A(n_1008),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_986),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_821),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1023),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_369),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_290),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1022),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_979),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_766),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_975),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_328),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_217),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_561),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_345),
.Y(n_1636)
);

INVx4_ASAP7_75t_R g1637 ( 
.A(n_21),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1029),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_378),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_882),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_575),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_764),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_876),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_677),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_284),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_623),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_245),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_407),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_505),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_843),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_227),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_657),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_641),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_16),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_278),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_910),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_572),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_389),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_532),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_336),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_858),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_250),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_987),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_161),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_985),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_999),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_827),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_867),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1457),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1047),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1125),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1167),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1127),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1044),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1456),
.Y(n_1676)
);

CKINVDCx16_ASAP7_75t_R g1677 ( 
.A(n_1240),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1485),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1408),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1408),
.Y(n_1680)
);

CKINVDCx16_ASAP7_75t_R g1681 ( 
.A(n_1326),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1545),
.Y(n_1682)
);

INVxp67_ASAP7_75t_SL g1683 ( 
.A(n_1177),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1634),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1408),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1237),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1067),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1381),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1276),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1067),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1342),
.Y(n_1691)
);

CKINVDCx14_ASAP7_75t_R g1692 ( 
.A(n_1193),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1193),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1074),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1581),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1207),
.Y(n_1696)
);

BUFx2_ASAP7_75t_SL g1697 ( 
.A(n_1078),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1520),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1329),
.B(n_1),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1231),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1408),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1311),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1520),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1351),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1078),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1421),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1074),
.Y(n_1707)
);

INVxp67_ASAP7_75t_SL g1708 ( 
.A(n_1177),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1035),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1037),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1408),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1040),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1408),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1045),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1046),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1208),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1614),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1614),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1054),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1348),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1060),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1408),
.Y(n_1722)
);

CKINVDCx16_ASAP7_75t_R g1723 ( 
.A(n_1407),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1439),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1062),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1063),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1072),
.Y(n_1727)
);

INVxp33_ASAP7_75t_L g1728 ( 
.A(n_1261),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1079),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1080),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1084),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1094),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1098),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1348),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1099),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1208),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1107),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1522),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1571),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1110),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1111),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1078),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1112),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1121),
.Y(n_1744)
);

INVx4_ASAP7_75t_R g1745 ( 
.A(n_1229),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1032),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1093),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1093),
.B(n_0),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1131),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1138),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1036),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1140),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1146),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1129),
.Y(n_1754)
);

INVxp33_ASAP7_75t_SL g1755 ( 
.A(n_1043),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1154),
.Y(n_1756)
);

CKINVDCx16_ASAP7_75t_R g1757 ( 
.A(n_1093),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1229),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1457),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1050),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1129),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1052),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1315),
.Y(n_1763)
);

CKINVDCx16_ASAP7_75t_R g1764 ( 
.A(n_1101),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1160),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1166),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1357),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1172),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1176),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1188),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1129),
.Y(n_1771)
);

CKINVDCx20_ASAP7_75t_R g1772 ( 
.A(n_1357),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1442),
.Y(n_1773)
);

CKINVDCx14_ASAP7_75t_R g1774 ( 
.A(n_1101),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1189),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1201),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1210),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1211),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1224),
.Y(n_1779)
);

INVxp33_ASAP7_75t_L g1780 ( 
.A(n_1041),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1225),
.Y(n_1781)
);

CKINVDCx14_ASAP7_75t_R g1782 ( 
.A(n_1101),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1228),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1315),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1233),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1238),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1243),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1380),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1247),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1251),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1252),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1257),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1263),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1380),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1268),
.B(n_2),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1266),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1129),
.B(n_0),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1272),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1274),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1275),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1283),
.Y(n_1801)
);

CKINVDCx16_ASAP7_75t_R g1802 ( 
.A(n_1153),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1129),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1457),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_1767),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1774),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1784),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1782),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1757),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1703),
.B(n_1064),
.Y(n_1810)
);

CKINVDCx20_ASAP7_75t_R g1811 ( 
.A(n_1772),
.Y(n_1811)
);

BUFx2_ASAP7_75t_SL g1812 ( 
.A(n_1742),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1688),
.Y(n_1813)
);

CKINVDCx20_ASAP7_75t_R g1814 ( 
.A(n_1764),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1794),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1705),
.B(n_1373),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1802),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1763),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1707),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1717),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1763),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1718),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1755),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1683),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1677),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1708),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1681),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1716),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1723),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1736),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1694),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1692),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1746),
.Y(n_1833)
);

CKINVDCx20_ASAP7_75t_R g1834 ( 
.A(n_1724),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1758),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1751),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1705),
.B(n_1042),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1788),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1671),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1760),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1672),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1674),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1696),
.B(n_1065),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1676),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1739),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1738),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1678),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1682),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1670),
.Y(n_1849)
);

CKINVDCx16_ASAP7_75t_R g1850 ( 
.A(n_1742),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1762),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1684),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1704),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1687),
.Y(n_1854)
);

INVxp67_ASAP7_75t_SL g1855 ( 
.A(n_1696),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1690),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1704),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1693),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1698),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1747),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1797),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_1747),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1675),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1720),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1734),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1797),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1697),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1773),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1709),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1675),
.B(n_1068),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1699),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1673),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1700),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1702),
.Y(n_1874)
);

INVxp67_ASAP7_75t_SL g1875 ( 
.A(n_1706),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1748),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1710),
.Y(n_1877)
);

CKINVDCx20_ASAP7_75t_R g1878 ( 
.A(n_1795),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1754),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1712),
.B(n_1075),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1686),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1689),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1691),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1695),
.Y(n_1884)
);

CKINVDCx16_ASAP7_75t_R g1885 ( 
.A(n_1728),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1714),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1715),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1719),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1721),
.Y(n_1889)
);

INVxp33_ASAP7_75t_SL g1890 ( 
.A(n_1745),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1725),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1726),
.Y(n_1892)
);

CKINVDCx16_ASAP7_75t_R g1893 ( 
.A(n_1727),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1729),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1730),
.B(n_1400),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1731),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1732),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1733),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1780),
.Y(n_1899)
);

INVxp67_ASAP7_75t_SL g1900 ( 
.A(n_1735),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1737),
.B(n_1519),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1740),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1741),
.B(n_1743),
.Y(n_1903)
);

CKINVDCx16_ASAP7_75t_R g1904 ( 
.A(n_1744),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1749),
.B(n_1623),
.Y(n_1905)
);

INVxp67_ASAP7_75t_L g1906 ( 
.A(n_1750),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1752),
.Y(n_1907)
);

CKINVDCx20_ASAP7_75t_R g1908 ( 
.A(n_1753),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1761),
.Y(n_1909)
);

INVxp67_ASAP7_75t_L g1910 ( 
.A(n_1756),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1765),
.Y(n_1911)
);

INVxp67_ASAP7_75t_L g1912 ( 
.A(n_1766),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1768),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1769),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1770),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1775),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1776),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1777),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1778),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1779),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1781),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1783),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1785),
.Y(n_1923)
);

INVxp67_ASAP7_75t_SL g1924 ( 
.A(n_1786),
.Y(n_1924)
);

NOR2xp67_ASAP7_75t_L g1925 ( 
.A(n_1787),
.B(n_1389),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1789),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_L g1927 ( 
.A(n_1790),
.B(n_1412),
.Y(n_1927)
);

INVxp67_ASAP7_75t_SL g1928 ( 
.A(n_1791),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1792),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1793),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1796),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1798),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1799),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1800),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1801),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1679),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1680),
.Y(n_1937)
);

INVxp33_ASAP7_75t_L g1938 ( 
.A(n_1685),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1701),
.Y(n_1939)
);

CKINVDCx20_ASAP7_75t_R g1940 ( 
.A(n_1711),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1713),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1722),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1771),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1803),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1670),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1670),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1759),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1759),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1759),
.B(n_1076),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1804),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1804),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1804),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1774),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1784),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1774),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1774),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1784),
.Y(n_1957)
);

BUFx2_ASAP7_75t_L g1958 ( 
.A(n_1774),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1724),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1784),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1784),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_R g1962 ( 
.A(n_1774),
.B(n_1077),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1774),
.Y(n_1963)
);

CKINVDCx20_ASAP7_75t_R g1964 ( 
.A(n_1767),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1705),
.B(n_1083),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1774),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1696),
.B(n_1153),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1774),
.Y(n_1968)
);

BUFx2_ASAP7_75t_L g1969 ( 
.A(n_1774),
.Y(n_1969)
);

INVxp67_ASAP7_75t_SL g1970 ( 
.A(n_1696),
.Y(n_1970)
);

CKINVDCx16_ASAP7_75t_R g1971 ( 
.A(n_1757),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1724),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1774),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1784),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1767),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1767),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1784),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_R g1978 ( 
.A(n_1774),
.B(n_1085),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1784),
.Y(n_1979)
);

CKINVDCx14_ASAP7_75t_R g1980 ( 
.A(n_1774),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1705),
.B(n_1087),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1774),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1767),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1784),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1774),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1705),
.B(n_1088),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1784),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1784),
.Y(n_1988)
);

INVxp33_ASAP7_75t_SL g1989 ( 
.A(n_1724),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1774),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1784),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1784),
.Y(n_1992)
);

CKINVDCx16_ASAP7_75t_R g1993 ( 
.A(n_1757),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1784),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1670),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1774),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1784),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1784),
.Y(n_1998)
);

CKINVDCx20_ASAP7_75t_R g1999 ( 
.A(n_1767),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1774),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1784),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1705),
.B(n_1089),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1774),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1784),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1784),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1767),
.Y(n_2006)
);

CKINVDCx20_ASAP7_75t_R g2007 ( 
.A(n_1767),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1784),
.Y(n_2008)
);

INVxp67_ASAP7_75t_SL g2009 ( 
.A(n_1696),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1784),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1784),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1784),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1784),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1774),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1784),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1784),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1774),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1784),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1705),
.B(n_1090),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1784),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1784),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1774),
.Y(n_2022)
);

BUFx2_ASAP7_75t_L g2023 ( 
.A(n_1774),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1784),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1774),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1774),
.Y(n_2026)
);

CKINVDCx20_ASAP7_75t_R g2027 ( 
.A(n_1767),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1774),
.Y(n_2028)
);

INVxp33_ASAP7_75t_SL g2029 ( 
.A(n_1724),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1774),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1784),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1724),
.B(n_1108),
.Y(n_2032)
);

CKINVDCx16_ASAP7_75t_R g2033 ( 
.A(n_1757),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1774),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1899),
.B(n_1855),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1861),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1866),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1813),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1850),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1924),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1815),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1924),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1928),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1928),
.B(n_1129),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1926),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1862),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1949),
.Y(n_2047)
);

OA21x2_ASAP7_75t_L g2048 ( 
.A1(n_1943),
.A2(n_1288),
.B(n_1284),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1839),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1841),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1869),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_1958),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1877),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1984),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1842),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1969),
.Y(n_2056)
);

AND2x6_ASAP7_75t_L g2057 ( 
.A(n_1967),
.B(n_1452),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1855),
.B(n_1153),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1886),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1844),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1847),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1848),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1888),
.B(n_1129),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1852),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1962),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1978),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1916),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1980),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1906),
.B(n_1910),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1970),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1970),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1912),
.B(n_1491),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1900),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_2023),
.B(n_1363),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1887),
.Y(n_2075)
);

AND2x6_ASAP7_75t_L g2076 ( 
.A(n_1853),
.B(n_1452),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1824),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1826),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1860),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_2018),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2009),
.B(n_1818),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1863),
.B(n_1893),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1806),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1889),
.A2(n_1894),
.B1(n_1902),
.B2(n_1892),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1891),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1828),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1896),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1812),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1821),
.B(n_1491),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1830),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1897),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1904),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_SL g2093 ( 
.A1(n_1805),
.A2(n_1964),
.B1(n_1975),
.B2(n_1811),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1835),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1843),
.B(n_1491),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_1885),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1908),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1838),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1875),
.A2(n_1100),
.B1(n_1103),
.B2(n_1096),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1898),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1903),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1880),
.B(n_1491),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1911),
.Y(n_2103)
);

BUFx2_ASAP7_75t_L g2104 ( 
.A(n_1919),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1959),
.B(n_1162),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_R g2106 ( 
.A(n_1808),
.B(n_1363),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1907),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1966),
.B(n_1370),
.Y(n_2108)
);

AND2x6_ASAP7_75t_L g2109 ( 
.A(n_1857),
.B(n_1455),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1971),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1917),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1965),
.B(n_1491),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_2034),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1923),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1953),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1972),
.B(n_1370),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1932),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1993),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1913),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_1955),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1914),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1915),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1918),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_SL g2124 ( 
.A(n_1823),
.B(n_1404),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1868),
.B(n_1162),
.Y(n_2125)
);

BUFx3_ASAP7_75t_L g2126 ( 
.A(n_1956),
.Y(n_2126)
);

AND2x4_ASAP7_75t_L g2127 ( 
.A(n_1963),
.B(n_1968),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1920),
.Y(n_2128)
);

AND2x6_ASAP7_75t_L g2129 ( 
.A(n_1922),
.B(n_1929),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1873),
.B(n_1162),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1973),
.Y(n_2131)
);

BUFx2_ASAP7_75t_L g2132 ( 
.A(n_1921),
.Y(n_2132)
);

OAI22xp5_ASAP7_75t_SL g2133 ( 
.A1(n_1976),
.A2(n_1418),
.B1(n_1459),
.B2(n_1404),
.Y(n_2133)
);

CKINVDCx20_ASAP7_75t_R g2134 ( 
.A(n_2033),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1874),
.B(n_1200),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_1933),
.Y(n_2136)
);

CKINVDCx11_ASAP7_75t_R g2137 ( 
.A(n_1814),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1930),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1931),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_1875),
.B(n_1200),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1982),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_1810),
.B(n_1981),
.Y(n_2142)
);

CKINVDCx11_ASAP7_75t_R g2143 ( 
.A(n_1983),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1935),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1925),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1986),
.B(n_1491),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1985),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1927),
.B(n_1381),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1945),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1990),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2002),
.B(n_2019),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_1870),
.Y(n_2152)
);

AND2x4_ASAP7_75t_L g2153 ( 
.A(n_1807),
.B(n_1470),
.Y(n_2153)
);

OA21x2_ASAP7_75t_L g2154 ( 
.A1(n_1944),
.A2(n_1291),
.B(n_1290),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1954),
.B(n_1470),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1946),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1996),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_2000),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1895),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_2003),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1901),
.Y(n_2161)
);

OA21x2_ASAP7_75t_L g2162 ( 
.A1(n_1936),
.A2(n_1294),
.B(n_1292),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_2014),
.Y(n_2163)
);

NOR2x1_ASAP7_75t_L g2164 ( 
.A(n_2032),
.B(n_1455),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_2017),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1957),
.B(n_1082),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1952),
.Y(n_2167)
);

INVx3_ASAP7_75t_L g2168 ( 
.A(n_2022),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_1960),
.B(n_1092),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1961),
.B(n_1097),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1837),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1816),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1876),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1905),
.B(n_1491),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1974),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_1977),
.B(n_1124),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1939),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1934),
.B(n_1200),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1941),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1979),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1879),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1987),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_2025),
.Y(n_2183)
);

NOR2xp67_ASAP7_75t_L g2184 ( 
.A(n_1809),
.B(n_1817),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1988),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_2026),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1991),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1992),
.Y(n_2188)
);

BUFx3_ASAP7_75t_L g2189 ( 
.A(n_2028),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1994),
.B(n_1150),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1997),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1938),
.B(n_1499),
.Y(n_2192)
);

CKINVDCx20_ASAP7_75t_R g2193 ( 
.A(n_1834),
.Y(n_2193)
);

AND2x2_ASAP7_75t_SL g2194 ( 
.A(n_1989),
.B(n_2029),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1937),
.B(n_1499),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1909),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1942),
.B(n_1998),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2001),
.B(n_1499),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1947),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1948),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_2030),
.Y(n_2201)
);

AND2x6_ASAP7_75t_L g2202 ( 
.A(n_2004),
.B(n_1488),
.Y(n_2202)
);

INVx3_ASAP7_75t_L g2203 ( 
.A(n_1867),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2005),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2008),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2010),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2011),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_1845),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_1950),
.A2(n_1137),
.B(n_1069),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1882),
.B(n_1220),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_2012),
.B(n_1104),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1872),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1999),
.Y(n_2213)
);

BUFx2_ASAP7_75t_L g2214 ( 
.A(n_1833),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2013),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2015),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_2006),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2016),
.B(n_1499),
.Y(n_2218)
);

AND2x4_ASAP7_75t_L g2219 ( 
.A(n_2020),
.B(n_1168),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2021),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2024),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2031),
.B(n_1418),
.Y(n_2222)
);

OA21x2_ASAP7_75t_L g2223 ( 
.A1(n_1951),
.A2(n_1303),
.B(n_1296),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1883),
.B(n_1220),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1836),
.Y(n_2225)
);

CKINVDCx20_ASAP7_75t_R g2226 ( 
.A(n_2007),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1940),
.B(n_1499),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1840),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_1851),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1881),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1884),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1890),
.B(n_1499),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_2027),
.Y(n_2233)
);

AND2x4_ASAP7_75t_SL g2234 ( 
.A(n_1846),
.B(n_1871),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1854),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1825),
.B(n_1459),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_1827),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1829),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1831),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1849),
.Y(n_2240)
);

CKINVDCx20_ASAP7_75t_R g2241 ( 
.A(n_1878),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_1856),
.Y(n_2242)
);

CKINVDCx20_ASAP7_75t_R g2243 ( 
.A(n_1859),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1832),
.B(n_1462),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_SL g2245 ( 
.A(n_1858),
.B(n_1462),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1819),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1864),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1865),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1820),
.B(n_1220),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1822),
.B(n_1109),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_1849),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_L g2252 ( 
.A(n_1849),
.B(n_1113),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1849),
.B(n_1499),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1995),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1995),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1995),
.Y(n_2256)
);

INVx4_ASAP7_75t_L g2257 ( 
.A(n_1995),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_1810),
.B(n_1114),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1861),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1813),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1861),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1813),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1813),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_1899),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1861),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1850),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1861),
.Y(n_2267)
);

CKINVDCx20_ASAP7_75t_R g2268 ( 
.A(n_1850),
.Y(n_2268)
);

BUFx2_ASAP7_75t_L g2269 ( 
.A(n_1899),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1855),
.B(n_1184),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_1850),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_1899),
.B(n_1242),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_1810),
.B(n_1115),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1861),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1813),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1813),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1861),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1813),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1861),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_1899),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_1861),
.B(n_1579),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1899),
.B(n_1242),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1861),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1813),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1813),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1813),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1850),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1850),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1889),
.B(n_1242),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1861),
.Y(n_2290)
);

BUFx3_ASAP7_75t_L g2291 ( 
.A(n_1958),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_1850),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_1850),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_1855),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_1958),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_1861),
.B(n_1579),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1813),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1958),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_1850),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_1899),
.B(n_1324),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1861),
.Y(n_2301)
);

INVx4_ASAP7_75t_L g2302 ( 
.A(n_1958),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_1855),
.B(n_1206),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1861),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1861),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_1861),
.Y(n_2306)
);

INVx3_ASAP7_75t_L g2307 ( 
.A(n_1850),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_1958),
.Y(n_2308)
);

CKINVDCx20_ASAP7_75t_R g2309 ( 
.A(n_1850),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_1850),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1813),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1861),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1958),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1958),
.Y(n_2314)
);

CKINVDCx20_ASAP7_75t_R g2315 ( 
.A(n_1850),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1813),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1861),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_1958),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1813),
.Y(n_2319)
);

INVx3_ASAP7_75t_L g2320 ( 
.A(n_1850),
.Y(n_2320)
);

OA21x2_ASAP7_75t_L g2321 ( 
.A1(n_1861),
.A2(n_1309),
.B(n_1306),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_1958),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_1810),
.B(n_1119),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_1850),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1861),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1889),
.B(n_1324),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_1958),
.Y(n_2327)
);

INVxp67_ASAP7_75t_L g2328 ( 
.A(n_1899),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1861),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1861),
.Y(n_2330)
);

OAI21x1_ASAP7_75t_L g2331 ( 
.A1(n_1861),
.A2(n_1137),
.B(n_1069),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_1861),
.A2(n_1123),
.B1(n_1128),
.B2(n_1122),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1861),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1861),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_1889),
.B(n_1324),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1861),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1813),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1861),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1850),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1861),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_1850),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_1899),
.B(n_1358),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2036),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2331),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2088),
.B(n_1132),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2037),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2259),
.B(n_2261),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2269),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2265),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2328),
.B(n_1066),
.Y(n_2350)
);

INVx5_ASAP7_75t_L g2351 ( 
.A(n_2129),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2267),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2274),
.B(n_1133),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2277),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2279),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2283),
.B(n_1134),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2290),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2301),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2304),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2305),
.Y(n_2360)
);

NAND3xp33_ASAP7_75t_L g2361 ( 
.A(n_2084),
.B(n_1139),
.C(n_1135),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2306),
.B(n_1141),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2269),
.B(n_1049),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2312),
.B(n_1142),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2317),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2325),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_SL g2367 ( 
.A(n_2329),
.B(n_2330),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_SL g2368 ( 
.A(n_2126),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2035),
.B(n_1477),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2056),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2333),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2334),
.Y(n_2372)
);

INVx1_ASAP7_75t_SL g2373 ( 
.A(n_2193),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2336),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2338),
.Y(n_2375)
);

AO21x2_ASAP7_75t_L g2376 ( 
.A1(n_2209),
.A2(n_1336),
.B(n_1321),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_2129),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2340),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2101),
.B(n_1143),
.Y(n_2379)
);

INVx8_ASAP7_75t_L g2380 ( 
.A(n_2052),
.Y(n_2380)
);

BUFx2_ASAP7_75t_L g2381 ( 
.A(n_2264),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_2152),
.B(n_1145),
.Y(n_2382)
);

INVx3_ASAP7_75t_L g2383 ( 
.A(n_2129),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2051),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2077),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2177),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2053),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2280),
.B(n_1073),
.Y(n_2388)
);

CKINVDCx6p67_ASAP7_75t_R g2389 ( 
.A(n_2137),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2082),
.B(n_1477),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_SL g2391 ( 
.A(n_2147),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2078),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2140),
.B(n_1148),
.Y(n_2393)
);

AOI21x1_ASAP7_75t_L g2394 ( 
.A1(n_2112),
.A2(n_1354),
.B(n_1337),
.Y(n_2394)
);

INVx4_ASAP7_75t_L g2395 ( 
.A(n_2080),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2058),
.B(n_1151),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2086),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2059),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2142),
.B(n_1152),
.Y(n_2399)
);

INVx8_ASAP7_75t_L g2400 ( 
.A(n_2052),
.Y(n_2400)
);

AO22x2_ASAP7_75t_L g2401 ( 
.A1(n_2116),
.A2(n_1406),
.B1(n_1149),
.B2(n_1157),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2090),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2069),
.B(n_1155),
.Y(n_2403)
);

AOI21x1_ASAP7_75t_L g2404 ( 
.A1(n_2146),
.A2(n_1367),
.B(n_1362),
.Y(n_2404)
);

INVx3_ASAP7_75t_L g2405 ( 
.A(n_2179),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2075),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2085),
.Y(n_2407)
);

AND3x2_ASAP7_75t_L g2408 ( 
.A(n_2124),
.B(n_1392),
.C(n_1057),
.Y(n_2408)
);

INVx1_ASAP7_75t_SL g2409 ( 
.A(n_2268),
.Y(n_2409)
);

INVx4_ASAP7_75t_L g2410 ( 
.A(n_2080),
.Y(n_2410)
);

CKINVDCx6p67_ASAP7_75t_R g2411 ( 
.A(n_2291),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2091),
.Y(n_2412)
);

BUFx6f_ASAP7_75t_SL g2413 ( 
.A(n_2189),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_2038),
.Y(n_2414)
);

INVx5_ASAP7_75t_L g2415 ( 
.A(n_2076),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2130),
.B(n_1156),
.Y(n_2416)
);

BUFx6f_ASAP7_75t_L g2417 ( 
.A(n_2321),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2094),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2295),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2100),
.Y(n_2420)
);

AND2x2_ASAP7_75t_SL g2421 ( 
.A(n_2194),
.B(n_1057),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2135),
.B(n_1161),
.Y(n_2422)
);

BUFx6f_ASAP7_75t_L g2423 ( 
.A(n_2321),
.Y(n_2423)
);

BUFx2_ASAP7_75t_L g2424 ( 
.A(n_2309),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2103),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2119),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2123),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2098),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_2210),
.B(n_1164),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2121),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2070),
.B(n_1165),
.Y(n_2431)
);

CKINVDCx6p67_ASAP7_75t_R g2432 ( 
.A(n_2143),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2128),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2122),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_2224),
.B(n_2105),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2178),
.B(n_1070),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_2107),
.B(n_1169),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2125),
.B(n_1086),
.Y(n_2438)
);

BUFx10_ASAP7_75t_L g2439 ( 
.A(n_2127),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2111),
.B(n_1170),
.Y(n_2440)
);

AO21x2_ASAP7_75t_L g2441 ( 
.A1(n_2151),
.A2(n_1371),
.B(n_1368),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2039),
.B(n_2287),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2138),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2139),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2144),
.Y(n_2445)
);

INVx1_ASAP7_75t_SL g2446 ( 
.A(n_2315),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2281),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2114),
.B(n_1171),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_SL g2449 ( 
.A(n_2117),
.B(n_1173),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2296),
.Y(n_2450)
);

INVx4_ASAP7_75t_L g2451 ( 
.A(n_2295),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2049),
.Y(n_2452)
);

OAI22xp5_ASAP7_75t_L g2453 ( 
.A1(n_2071),
.A2(n_1126),
.B1(n_1178),
.B2(n_1095),
.Y(n_2453)
);

BUFx10_ASAP7_75t_L g2454 ( 
.A(n_2225),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2292),
.B(n_1183),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2067),
.B(n_1202),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2260),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2262),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2050),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2045),
.B(n_1216),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2055),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2263),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2040),
.B(n_1174),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2299),
.B(n_1218),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2275),
.Y(n_2465)
);

NAND2xp33_ASAP7_75t_L g2466 ( 
.A(n_2076),
.B(n_1579),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2060),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2276),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2061),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2062),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2064),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2307),
.B(n_2310),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2044),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2266),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2042),
.B(n_1175),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2278),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2284),
.Y(n_2477)
);

INVx1_ASAP7_75t_SL g2478 ( 
.A(n_2208),
.Y(n_2478)
);

NAND2xp33_ASAP7_75t_SL g2479 ( 
.A(n_2079),
.B(n_1392),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2285),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2048),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2048),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2271),
.Y(n_2483)
);

AOI21x1_ASAP7_75t_L g2484 ( 
.A1(n_2102),
.A2(n_2095),
.B(n_2253),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2154),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2154),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2286),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_2162),
.Y(n_2488)
);

NOR2x1p5_ASAP7_75t_L g2489 ( 
.A(n_2320),
.B(n_1179),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2272),
.B(n_2282),
.Y(n_2490)
);

NOR2x1p5_ASAP7_75t_L g2491 ( 
.A(n_2324),
.B(n_1180),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2162),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2043),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2341),
.B(n_1219),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2073),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_2332),
.B(n_1181),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2300),
.B(n_1267),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2047),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2342),
.B(n_1273),
.Y(n_2499)
);

INVxp67_ASAP7_75t_SL g2500 ( 
.A(n_2092),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2214),
.B(n_1297),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_2298),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2172),
.B(n_1182),
.Y(n_2503)
);

INVx3_ASAP7_75t_L g2504 ( 
.A(n_2297),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2270),
.B(n_1185),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2046),
.B(n_1120),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2311),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2316),
.Y(n_2508)
);

INVx5_ASAP7_75t_L g2509 ( 
.A(n_2076),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2319),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2159),
.B(n_1186),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2161),
.B(n_1190),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_2337),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2181),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2214),
.B(n_1341),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2196),
.Y(n_2516)
);

NAND2xp33_ASAP7_75t_SL g2517 ( 
.A(n_2288),
.B(n_2293),
.Y(n_2517)
);

INVx3_ASAP7_75t_L g2518 ( 
.A(n_2109),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2089),
.Y(n_2519)
);

INVx3_ASAP7_75t_L g2520 ( 
.A(n_2109),
.Y(n_2520)
);

NOR2xp33_ASAP7_75t_L g2521 ( 
.A(n_2173),
.B(n_1478),
.Y(n_2521)
);

NAND2xp33_ASAP7_75t_L g2522 ( 
.A(n_2109),
.B(n_1579),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2223),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2223),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2270),
.B(n_1192),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2255),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2175),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2257),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2198),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2099),
.B(n_1194),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2218),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2199),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2200),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2171),
.B(n_1195),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2192),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2303),
.B(n_1196),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2303),
.B(n_1197),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2063),
.Y(n_2538)
);

AND3x2_ASAP7_75t_L g2539 ( 
.A(n_2245),
.B(n_1501),
.C(n_1493),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2212),
.B(n_1198),
.Y(n_2540)
);

AO21x2_ASAP7_75t_L g2541 ( 
.A1(n_2195),
.A2(n_1375),
.B(n_1374),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2072),
.Y(n_2542)
);

BUFx6f_ASAP7_75t_L g2543 ( 
.A(n_2298),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2208),
.B(n_1159),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2180),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2057),
.B(n_1199),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2182),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2251),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2057),
.B(n_1204),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2339),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2197),
.B(n_1503),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2185),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2148),
.Y(n_2553)
);

BUFx10_ASAP7_75t_L g2554 ( 
.A(n_2225),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2148),
.Y(n_2555)
);

BUFx6f_ASAP7_75t_L g2556 ( 
.A(n_2308),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2294),
.B(n_1205),
.Y(n_2557)
);

NAND2xp33_ASAP7_75t_L g2558 ( 
.A(n_2057),
.B(n_1579),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2187),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2258),
.B(n_1209),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2188),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2191),
.Y(n_2562)
);

AO21x2_ASAP7_75t_L g2563 ( 
.A1(n_2174),
.A2(n_2227),
.B(n_2252),
.Y(n_2563)
);

CKINVDCx6p67_ASAP7_75t_R g2564 ( 
.A(n_2302),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2145),
.Y(n_2565)
);

NAND3xp33_ASAP7_75t_L g2566 ( 
.A(n_2273),
.B(n_1215),
.C(n_1212),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_2308),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2164),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2203),
.B(n_1217),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2204),
.Y(n_2570)
);

INVx4_ASAP7_75t_L g2571 ( 
.A(n_2313),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2041),
.B(n_2054),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2136),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2205),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2206),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2106),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2243),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2207),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2215),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2216),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2289),
.B(n_1532),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2220),
.Y(n_2582)
);

BUFx10_ASAP7_75t_L g2583 ( 
.A(n_2229),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2221),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2149),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2081),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2153),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2153),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2241),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2155),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2155),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2323),
.B(n_1221),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2166),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2166),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2169),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2169),
.B(n_1222),
.Y(n_2596)
);

INVx2_ASAP7_75t_SL g2597 ( 
.A(n_2313),
.Y(n_2597)
);

AND3x2_ASAP7_75t_L g2598 ( 
.A(n_2087),
.B(n_1564),
.C(n_1553),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2170),
.Y(n_2599)
);

CKINVDCx6p67_ASAP7_75t_R g2600 ( 
.A(n_2134),
.Y(n_2600)
);

INVxp33_ASAP7_75t_L g2601 ( 
.A(n_2096),
.Y(n_2601)
);

NAND3xp33_ASAP7_75t_L g2602 ( 
.A(n_2250),
.B(n_1226),
.C(n_1223),
.Y(n_2602)
);

INVxp67_ASAP7_75t_SL g2603 ( 
.A(n_2314),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2314),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2170),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2176),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2087),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2156),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2176),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2190),
.Y(n_2610)
);

CKINVDCx6p67_ASAP7_75t_R g2611 ( 
.A(n_2226),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2190),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2219),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2219),
.Y(n_2614)
);

BUFx10_ASAP7_75t_L g2615 ( 
.A(n_2229),
.Y(n_2615)
);

INVx8_ASAP7_75t_L g2616 ( 
.A(n_2318),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2202),
.B(n_1227),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2167),
.Y(n_2618)
);

INVx3_ASAP7_75t_L g2619 ( 
.A(n_2202),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2097),
.Y(n_2620)
);

NAND2xp33_ASAP7_75t_L g2621 ( 
.A(n_2202),
.B(n_1579),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2254),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2240),
.Y(n_2623)
);

NAND3xp33_ASAP7_75t_L g2624 ( 
.A(n_2211),
.B(n_1232),
.C(n_1230),
.Y(n_2624)
);

INVx4_ASAP7_75t_L g2625 ( 
.A(n_2318),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2222),
.B(n_1568),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2256),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2249),
.B(n_1574),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2232),
.Y(n_2629)
);

BUFx2_ASAP7_75t_L g2630 ( 
.A(n_2097),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2326),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2335),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2322),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2322),
.B(n_1234),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2327),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2327),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2248),
.Y(n_2637)
);

NOR2x1p5_ASAP7_75t_L g2638 ( 
.A(n_2246),
.B(n_1236),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_SL g2639 ( 
.A(n_2083),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2235),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2228),
.B(n_1241),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2104),
.Y(n_2642)
);

INVxp67_ASAP7_75t_L g2643 ( 
.A(n_2104),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2150),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2242),
.B(n_1608),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2132),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_2074),
.B(n_1615),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2108),
.B(n_2132),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2163),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2247),
.B(n_1244),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2230),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2231),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2213),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2165),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2247),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2237),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2238),
.Y(n_2657)
);

NAND2xp33_ASAP7_75t_L g2658 ( 
.A(n_2065),
.B(n_1579),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2168),
.B(n_1245),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2184),
.B(n_1246),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2083),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2113),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2113),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2115),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2115),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_SL g2666 ( 
.A(n_2066),
.B(n_1249),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2120),
.Y(n_2667)
);

AOI21x1_ASAP7_75t_L g2668 ( 
.A1(n_2236),
.A2(n_1386),
.B(n_1382),
.Y(n_2668)
);

INVxp33_ASAP7_75t_L g2669 ( 
.A(n_2093),
.Y(n_2669)
);

INVxp67_ASAP7_75t_L g2670 ( 
.A(n_2133),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2120),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2131),
.Y(n_2672)
);

INVx3_ASAP7_75t_SL g2673 ( 
.A(n_2068),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2131),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2141),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2234),
.B(n_1668),
.Y(n_2676)
);

AND3x2_ASAP7_75t_L g2677 ( 
.A(n_2244),
.B(n_1081),
.C(n_1033),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2141),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2157),
.B(n_1253),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2157),
.Y(n_2680)
);

OR2x2_ASAP7_75t_L g2681 ( 
.A(n_2217),
.B(n_1203),
.Y(n_2681)
);

AO21x2_ASAP7_75t_L g2682 ( 
.A1(n_2158),
.A2(n_1417),
.B(n_1414),
.Y(n_2682)
);

INVx5_ASAP7_75t_L g2683 ( 
.A(n_2158),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2186),
.B(n_1256),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2186),
.Y(n_2685)
);

INVxp33_ASAP7_75t_L g2686 ( 
.A(n_2233),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2110),
.Y(n_2687)
);

INVx2_ASAP7_75t_SL g2688 ( 
.A(n_2118),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2160),
.B(n_1258),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2183),
.B(n_1259),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2201),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2239),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2331),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2088),
.B(n_1260),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2331),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2331),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2088),
.B(n_1264),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2129),
.Y(n_2698)
);

AND2x4_ASAP7_75t_L g2699 ( 
.A(n_2101),
.B(n_1279),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2331),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2193),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2331),
.Y(n_2702)
);

INVx3_ASAP7_75t_L g2703 ( 
.A(n_2129),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2036),
.Y(n_2704)
);

AND2x2_ASAP7_75t_SL g2705 ( 
.A(n_2194),
.B(n_1102),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2331),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2331),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2036),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2331),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_SL g2710 ( 
.A(n_2126),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2088),
.B(n_1270),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2328),
.B(n_1271),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2036),
.Y(n_2713)
);

BUFx3_ASAP7_75t_L g2714 ( 
.A(n_2056),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2036),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2036),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2331),
.Y(n_2717)
);

INVx3_ASAP7_75t_L g2718 ( 
.A(n_2129),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2331),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2036),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_2129),
.Y(n_2721)
);

NAND3x1_ASAP7_75t_L g2722 ( 
.A(n_2039),
.B(n_1591),
.C(n_1340),
.Y(n_2722)
);

INVx2_ASAP7_75t_SL g2723 ( 
.A(n_2269),
.Y(n_2723)
);

BUFx3_ASAP7_75t_L g2724 ( 
.A(n_2056),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2036),
.Y(n_2725)
);

INVxp33_ASAP7_75t_L g2726 ( 
.A(n_2264),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2328),
.B(n_1278),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2036),
.B(n_1281),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2331),
.Y(n_2729)
);

BUFx10_ASAP7_75t_L g2730 ( 
.A(n_2088),
.Y(n_2730)
);

NOR3xp33_ASAP7_75t_L g2731 ( 
.A(n_2133),
.B(n_1280),
.C(n_1235),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2331),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2331),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2036),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_2088),
.B(n_1282),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2343),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2734),
.Y(n_2737)
);

INVxp67_ASAP7_75t_SL g2738 ( 
.A(n_2698),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2352),
.Y(n_2739)
);

INVxp33_ASAP7_75t_SL g2740 ( 
.A(n_2453),
.Y(n_2740)
);

BUFx6f_ASAP7_75t_L g2741 ( 
.A(n_2543),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2543),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2355),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2380),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_2381),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2357),
.Y(n_2746)
);

INVx2_ASAP7_75t_SL g2747 ( 
.A(n_2380),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2586),
.B(n_1289),
.Y(n_2748)
);

OR2x6_ASAP7_75t_L g2749 ( 
.A(n_2400),
.B(n_1059),
.Y(n_2749)
);

BUFx10_ASAP7_75t_L g2750 ( 
.A(n_2639),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2360),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2346),
.B(n_1295),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2365),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2348),
.B(n_1300),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2372),
.Y(n_2755)
);

BUFx3_ASAP7_75t_L g2756 ( 
.A(n_2400),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2369),
.B(n_1358),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2723),
.B(n_1358),
.Y(n_2758)
);

INVx5_ASAP7_75t_L g2759 ( 
.A(n_2616),
.Y(n_2759)
);

INVx2_ASAP7_75t_SL g2760 ( 
.A(n_2616),
.Y(n_2760)
);

INVx4_ASAP7_75t_L g2761 ( 
.A(n_2564),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2346),
.B(n_1301),
.Y(n_2762)
);

BUFx6f_ASAP7_75t_L g2763 ( 
.A(n_2543),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2556),
.B(n_1488),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2350),
.A2(n_1302),
.B1(n_1307),
.B2(n_1305),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2375),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2349),
.B(n_2354),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2556),
.B(n_1589),
.Y(n_2768)
);

NOR2xp33_ASAP7_75t_L g2769 ( 
.A(n_2438),
.B(n_2551),
.Y(n_2769)
);

BUFx6f_ASAP7_75t_L g2770 ( 
.A(n_2556),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2349),
.B(n_1310),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2452),
.Y(n_2772)
);

NAND2xp33_ASAP7_75t_L g2773 ( 
.A(n_2698),
.B(n_1313),
.Y(n_2773)
);

INVx4_ASAP7_75t_L g2774 ( 
.A(n_2567),
.Y(n_2774)
);

AND2x4_ASAP7_75t_L g2775 ( 
.A(n_2567),
.B(n_2604),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2698),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2452),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2459),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2497),
.B(n_1314),
.Y(n_2779)
);

INVx4_ASAP7_75t_L g2780 ( 
.A(n_2567),
.Y(n_2780)
);

AND2x6_ASAP7_75t_L g2781 ( 
.A(n_2721),
.B(n_1589),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2604),
.B(n_1590),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2370),
.Y(n_2783)
);

INVxp67_ASAP7_75t_L g2784 ( 
.A(n_2363),
.Y(n_2784)
);

BUFx6f_ASAP7_75t_L g2785 ( 
.A(n_2604),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2721),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_2721),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2447),
.A2(n_1319),
.B1(n_1320),
.B2(n_1318),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2378),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2390),
.B(n_1415),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_2683),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2354),
.Y(n_2792)
);

INVx6_ASAP7_75t_L g2793 ( 
.A(n_2454),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_SL g2794 ( 
.A(n_2388),
.B(n_1323),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2460),
.A2(n_1415),
.B1(n_1655),
.B2(n_1590),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2358),
.B(n_1325),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2358),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2359),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2359),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2351),
.B(n_1327),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2366),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2366),
.B(n_1328),
.Y(n_2802)
);

INVx4_ASAP7_75t_L g2803 ( 
.A(n_2683),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2371),
.B(n_1331),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_L g2805 ( 
.A(n_2351),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2371),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2374),
.B(n_1332),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2374),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2704),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2704),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2708),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2708),
.B(n_1333),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2713),
.B(n_1334),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2713),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2715),
.B(n_1338),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2499),
.B(n_1344),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2351),
.B(n_1346),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2715),
.Y(n_2818)
);

INVx3_ASAP7_75t_L g2819 ( 
.A(n_2377),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2417),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2716),
.B(n_1350),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2716),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2720),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2720),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2725),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2459),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2725),
.B(n_1353),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2574),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2377),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2714),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2527),
.B(n_1355),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2417),
.Y(n_2832)
);

INVx1_ASAP7_75t_SL g2833 ( 
.A(n_2411),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2575),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2495),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2578),
.Y(n_2836)
);

AOI21x1_ASAP7_75t_L g2837 ( 
.A1(n_2481),
.A2(n_1213),
.B(n_1158),
.Y(n_2837)
);

BUFx10_ASAP7_75t_L g2838 ( 
.A(n_2639),
.Y(n_2838)
);

CKINVDCx20_ASAP7_75t_R g2839 ( 
.A(n_2389),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2579),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2501),
.B(n_1285),
.Y(n_2841)
);

AND2x2_ASAP7_75t_SL g2842 ( 
.A(n_2421),
.B(n_1158),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2545),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2547),
.B(n_2552),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2383),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2515),
.B(n_1415),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2559),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2561),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_SL g2849 ( 
.A(n_2726),
.B(n_1359),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_2417),
.Y(n_2850)
);

INVx2_ASAP7_75t_SL g2851 ( 
.A(n_2454),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2562),
.B(n_1361),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_2415),
.B(n_2509),
.Y(n_2853)
);

INVx3_ASAP7_75t_L g2854 ( 
.A(n_2383),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2570),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2584),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2435),
.B(n_2628),
.Y(n_2857)
);

INVx2_ASAP7_75t_SL g2858 ( 
.A(n_2554),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2580),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2582),
.B(n_1655),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2385),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2415),
.B(n_2509),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2461),
.B(n_1364),
.Y(n_2863)
);

INVxp67_ASAP7_75t_SL g2864 ( 
.A(n_2548),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2461),
.Y(n_2865)
);

AO21x2_ASAP7_75t_L g2866 ( 
.A1(n_2481),
.A2(n_1438),
.B(n_1430),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2469),
.B(n_2470),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2469),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_2640),
.B(n_1293),
.Y(n_2869)
);

BUFx6f_ASAP7_75t_L g2870 ( 
.A(n_2423),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2415),
.B(n_1365),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2470),
.B(n_1366),
.Y(n_2872)
);

BUFx3_ASAP7_75t_L g2873 ( 
.A(n_2683),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2471),
.B(n_1369),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2392),
.Y(n_2875)
);

INVx4_ASAP7_75t_L g2876 ( 
.A(n_2554),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2471),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2493),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2436),
.B(n_1167),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2637),
.B(n_1339),
.Y(n_2880)
);

OAI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2670),
.A2(n_1376),
.B1(n_1379),
.B2(n_1372),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2478),
.B(n_1383),
.Y(n_2882)
);

NAND2x1p5_ASAP7_75t_L g2883 ( 
.A(n_2724),
.B(n_2451),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2397),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2402),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2699),
.B(n_1387),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2418),
.Y(n_2887)
);

OAI21xp33_ASAP7_75t_L g2888 ( 
.A1(n_2399),
.A2(n_1390),
.B(n_1388),
.Y(n_2888)
);

INVx2_ASAP7_75t_SL g2889 ( 
.A(n_2583),
.Y(n_2889)
);

INVx4_ASAP7_75t_L g2890 ( 
.A(n_2583),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2509),
.B(n_1393),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_2432),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2447),
.A2(n_1396),
.B1(n_1397),
.B2(n_1394),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_2611),
.Y(n_2894)
);

INVx1_ASAP7_75t_SL g2895 ( 
.A(n_2506),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2428),
.Y(n_2896)
);

INVx4_ASAP7_75t_L g2897 ( 
.A(n_2615),
.Y(n_2897)
);

AOI22xp33_ASAP7_75t_SL g2898 ( 
.A1(n_2401),
.A2(n_1167),
.B1(n_1286),
.B2(n_1399),
.Y(n_2898)
);

INVx3_ASAP7_75t_L g2899 ( 
.A(n_2703),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2699),
.B(n_1402),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2430),
.Y(n_2901)
);

INVx4_ASAP7_75t_L g2902 ( 
.A(n_2615),
.Y(n_2902)
);

INVx5_ASAP7_75t_L g2903 ( 
.A(n_2451),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2434),
.Y(n_2904)
);

INVx2_ASAP7_75t_SL g2905 ( 
.A(n_2730),
.Y(n_2905)
);

HB1xp67_ASAP7_75t_L g2906 ( 
.A(n_2607),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2467),
.Y(n_2907)
);

INVxp67_ASAP7_75t_L g2908 ( 
.A(n_2681),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2703),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2498),
.Y(n_2910)
);

INVx5_ASAP7_75t_L g2911 ( 
.A(n_2571),
.Y(n_2911)
);

INVx4_ASAP7_75t_L g2912 ( 
.A(n_2571),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2384),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2456),
.A2(n_1405),
.B1(n_1410),
.B2(n_1409),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2595),
.Y(n_2915)
);

AND2x2_ASAP7_75t_SL g2916 ( 
.A(n_2705),
.B(n_1213),
.Y(n_2916)
);

INVx4_ASAP7_75t_L g2917 ( 
.A(n_2625),
.Y(n_2917)
);

INVx1_ASAP7_75t_SL g2918 ( 
.A(n_2620),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2479),
.B(n_1413),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2387),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2398),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2599),
.Y(n_2922)
);

NAND3xp33_ASAP7_75t_L g2923 ( 
.A(n_2566),
.B(n_1669),
.C(n_1419),
.Y(n_2923)
);

AND2x6_ASAP7_75t_L g2924 ( 
.A(n_2718),
.B(n_1048),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2605),
.Y(n_2925)
);

NAND2x1p5_ASAP7_75t_L g2926 ( 
.A(n_2625),
.B(n_1308),
.Y(n_2926)
);

BUFx6f_ASAP7_75t_L g2927 ( 
.A(n_2423),
.Y(n_2927)
);

INVx4_ASAP7_75t_L g2928 ( 
.A(n_2539),
.Y(n_2928)
);

INVx3_ASAP7_75t_L g2929 ( 
.A(n_2718),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2606),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2423),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2613),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2614),
.Y(n_2933)
);

INVx1_ASAP7_75t_SL g2934 ( 
.A(n_2630),
.Y(n_2934)
);

INVx3_ASAP7_75t_L g2935 ( 
.A(n_2518),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2408),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2379),
.B(n_1416),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2406),
.Y(n_2938)
);

BUFx4f_ASAP7_75t_L g2939 ( 
.A(n_2600),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2593),
.Y(n_2940)
);

NOR3xp33_ASAP7_75t_L g2941 ( 
.A(n_2490),
.B(n_2361),
.C(n_2416),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_R g2942 ( 
.A(n_2577),
.B(n_1424),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2730),
.B(n_2712),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2594),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2601),
.B(n_1426),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2609),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2401),
.B(n_1286),
.Y(n_2947)
);

AND2x4_ASAP7_75t_L g2948 ( 
.A(n_2610),
.B(n_2612),
.Y(n_2948)
);

OAI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2450),
.A2(n_1428),
.B1(n_1431),
.B2(n_1427),
.Y(n_2949)
);

BUFx6f_ASAP7_75t_L g2950 ( 
.A(n_2486),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2407),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2450),
.A2(n_1435),
.B1(n_1436),
.B2(n_1433),
.Y(n_2952)
);

OR2x6_ASAP7_75t_L g2953 ( 
.A(n_2701),
.B(n_1059),
.Y(n_2953)
);

INVx4_ASAP7_75t_L g2954 ( 
.A(n_2419),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2412),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2645),
.B(n_1286),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_L g2957 ( 
.A(n_2486),
.Y(n_2957)
);

INVxp33_ASAP7_75t_L g2958 ( 
.A(n_2676),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2420),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_L g2960 ( 
.A(n_2486),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2425),
.Y(n_2961)
);

INVx5_ASAP7_75t_L g2962 ( 
.A(n_2395),
.Y(n_2962)
);

AND2x6_ASAP7_75t_L g2963 ( 
.A(n_2518),
.B(n_1048),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2426),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_2520),
.Y(n_2965)
);

INVxp67_ASAP7_75t_SL g2966 ( 
.A(n_2573),
.Y(n_2966)
);

INVx4_ASAP7_75t_SL g2967 ( 
.A(n_2368),
.Y(n_2967)
);

NAND2xp33_ASAP7_75t_L g2968 ( 
.A(n_2488),
.B(n_1445),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2427),
.Y(n_2969)
);

NOR2xp33_ASAP7_75t_L g2970 ( 
.A(n_2643),
.B(n_2647),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2433),
.Y(n_2971)
);

BUFx2_ASAP7_75t_L g2972 ( 
.A(n_2455),
.Y(n_2972)
);

BUFx6f_ASAP7_75t_L g2973 ( 
.A(n_2488),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2347),
.B(n_1437),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2443),
.Y(n_2975)
);

AO22x2_ASAP7_75t_L g2976 ( 
.A1(n_2482),
.A2(n_1330),
.B1(n_1335),
.B2(n_1322),
.Y(n_2976)
);

AND2x4_ASAP7_75t_L g2977 ( 
.A(n_2395),
.B(n_1343),
.Y(n_2977)
);

BUFx3_ASAP7_75t_L g2978 ( 
.A(n_2662),
.Y(n_2978)
);

OR2x6_ASAP7_75t_L g2979 ( 
.A(n_2589),
.B(n_1136),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2444),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2410),
.B(n_1471),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2445),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2727),
.B(n_1440),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2410),
.B(n_1505),
.Y(n_2984)
);

OR2x2_ASAP7_75t_L g2985 ( 
.A(n_2373),
.B(n_1517),
.Y(n_2985)
);

INVx1_ASAP7_75t_SL g2986 ( 
.A(n_2544),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2353),
.B(n_1441),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2626),
.B(n_1443),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2728),
.B(n_2393),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2396),
.B(n_1444),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2463),
.B(n_1446),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2386),
.Y(n_2992)
);

INVx3_ASAP7_75t_L g2993 ( 
.A(n_2520),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2651),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2652),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2386),
.Y(n_2996)
);

NAND2x1p5_ASAP7_75t_L g2997 ( 
.A(n_2662),
.B(n_1403),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2588),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2587),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2590),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2405),
.Y(n_3001)
);

INVx4_ASAP7_75t_L g3002 ( 
.A(n_2368),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2521),
.B(n_1447),
.Y(n_3003)
);

NOR2xp33_ASAP7_75t_SL g3004 ( 
.A(n_2576),
.B(n_1448),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2475),
.B(n_1449),
.Y(n_3005)
);

INVx1_ASAP7_75t_SL g3006 ( 
.A(n_2472),
.Y(n_3006)
);

CKINVDCx5p33_ASAP7_75t_R g3007 ( 
.A(n_2653),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2591),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2431),
.B(n_1450),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2405),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2441),
.B(n_1451),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2514),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_2488),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2464),
.B(n_1458),
.Y(n_3014)
);

INVx3_ASAP7_75t_L g3015 ( 
.A(n_2619),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2516),
.Y(n_3016)
);

OAI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2669),
.A2(n_1461),
.B1(n_1463),
.B2(n_1460),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2581),
.B(n_1465),
.Y(n_3018)
);

AO22x2_ASAP7_75t_L g3019 ( 
.A1(n_2482),
.A2(n_1432),
.B1(n_1489),
.B2(n_1425),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2494),
.Y(n_3020)
);

BUFx2_ASAP7_75t_L g3021 ( 
.A(n_2598),
.Y(n_3021)
);

BUFx2_ASAP7_75t_L g3022 ( 
.A(n_2474),
.Y(n_3022)
);

NAND2x1p5_ASAP7_75t_L g3023 ( 
.A(n_2665),
.B(n_1494),
.Y(n_3023)
);

INVx3_ASAP7_75t_L g3024 ( 
.A(n_2619),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2505),
.B(n_2525),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2483),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2532),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2533),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2629),
.B(n_1466),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2422),
.B(n_1467),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2553),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2555),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2668),
.Y(n_3033)
);

INVx2_ASAP7_75t_SL g3034 ( 
.A(n_2439),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2409),
.B(n_1556),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2457),
.Y(n_3036)
);

AND2x6_ASAP7_75t_L g3037 ( 
.A(n_2473),
.B(n_1048),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_2429),
.B(n_2642),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2458),
.Y(n_3039)
);

AO22x2_ASAP7_75t_L g3040 ( 
.A1(n_2485),
.A2(n_1665),
.B1(n_1633),
.B2(n_1250),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2462),
.Y(n_3041)
);

AND3x4_ASAP7_75t_L g3042 ( 
.A(n_2731),
.B(n_1239),
.C(n_1136),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_2446),
.B(n_1469),
.Y(n_3043)
);

BUFx3_ASAP7_75t_L g3044 ( 
.A(n_2665),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2536),
.B(n_1474),
.Y(n_3045)
);

AND2x4_ASAP7_75t_L g3046 ( 
.A(n_2585),
.B(n_1507),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2523),
.Y(n_3047)
);

CKINVDCx5p33_ASAP7_75t_R g3048 ( 
.A(n_2673),
.Y(n_3048)
);

BUFx4f_ASAP7_75t_L g3049 ( 
.A(n_2692),
.Y(n_3049)
);

OR2x2_ASAP7_75t_L g3050 ( 
.A(n_2596),
.B(n_1476),
.Y(n_3050)
);

INVx4_ASAP7_75t_L g3051 ( 
.A(n_2391),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2465),
.Y(n_3052)
);

NOR2x1p5_ASAP7_75t_L g3053 ( 
.A(n_2692),
.B(n_1480),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2468),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2537),
.B(n_1481),
.Y(n_3055)
);

AOI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2648),
.A2(n_1495),
.B1(n_1496),
.B2(n_1490),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2476),
.Y(n_3057)
);

OAI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2473),
.A2(n_1502),
.B1(n_1504),
.B2(n_1497),
.Y(n_3058)
);

INVx1_ASAP7_75t_SL g3059 ( 
.A(n_2442),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_L g3060 ( 
.A(n_2524),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2656),
.B(n_2657),
.Y(n_3061)
);

BUFx6f_ASAP7_75t_L g3062 ( 
.A(n_2344),
.Y(n_3062)
);

OR2x2_ASAP7_75t_L g3063 ( 
.A(n_2550),
.B(n_1506),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2477),
.Y(n_3064)
);

INVx3_ASAP7_75t_L g3065 ( 
.A(n_2585),
.Y(n_3065)
);

AND2x4_ASAP7_75t_L g3066 ( 
.A(n_2608),
.B(n_1509),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2693),
.Y(n_3067)
);

BUFx6f_ASAP7_75t_L g3068 ( 
.A(n_2695),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2391),
.Y(n_3069)
);

INVx2_ASAP7_75t_SL g3070 ( 
.A(n_2439),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2480),
.Y(n_3071)
);

CKINVDCx8_ASAP7_75t_R g3072 ( 
.A(n_2424),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2659),
.B(n_1511),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2487),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2507),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2646),
.B(n_2382),
.Y(n_3076)
);

BUFx6f_ASAP7_75t_L g3077 ( 
.A(n_2696),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2508),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_SL g3079 ( 
.A(n_2617),
.B(n_1513),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2510),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2565),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2367),
.Y(n_3082)
);

AND2x4_ASAP7_75t_L g3083 ( 
.A(n_2608),
.B(n_1516),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2650),
.B(n_1514),
.Y(n_3084)
);

BUFx3_ASAP7_75t_L g3085 ( 
.A(n_2502),
.Y(n_3085)
);

OR2x6_ASAP7_75t_L g3086 ( 
.A(n_2722),
.B(n_1239),
.Y(n_3086)
);

INVx4_ASAP7_75t_L g3087 ( 
.A(n_2413),
.Y(n_3087)
);

NOR2x1p5_ASAP7_75t_L g3088 ( 
.A(n_2691),
.B(n_1515),
.Y(n_3088)
);

BUFx2_ASAP7_75t_L g3089 ( 
.A(n_2677),
.Y(n_3089)
);

OAI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_2686),
.A2(n_1525),
.B1(n_1528),
.B2(n_1523),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_2489),
.B(n_1530),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_2546),
.B(n_1531),
.Y(n_3092)
);

INVx4_ASAP7_75t_SL g3093 ( 
.A(n_2413),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_L g3094 ( 
.A(n_2700),
.Y(n_3094)
);

AND2x4_ASAP7_75t_L g3095 ( 
.A(n_2618),
.B(n_1518),
.Y(n_3095)
);

AND2x6_ASAP7_75t_L g3096 ( 
.A(n_2519),
.B(n_1048),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2702),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2414),
.Y(n_3098)
);

INVx3_ASAP7_75t_L g3099 ( 
.A(n_2618),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_2528),
.Y(n_3100)
);

BUFx6f_ASAP7_75t_L g3101 ( 
.A(n_2706),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_SL g3102 ( 
.A(n_2549),
.B(n_2597),
.Y(n_3102)
);

INVx3_ASAP7_75t_L g3103 ( 
.A(n_2414),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2504),
.Y(n_3104)
);

INVx5_ASAP7_75t_L g3105 ( 
.A(n_2661),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2504),
.Y(n_3106)
);

OR2x6_ASAP7_75t_L g3107 ( 
.A(n_2688),
.B(n_2638),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2513),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2513),
.Y(n_3109)
);

AND2x6_ASAP7_75t_L g3110 ( 
.A(n_2529),
.B(n_1051),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2560),
.B(n_1535),
.Y(n_3111)
);

BUFx4f_ASAP7_75t_L g3112 ( 
.A(n_2687),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2568),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2557),
.A2(n_1537),
.B1(n_1540),
.B2(n_1536),
.Y(n_3114)
);

BUFx3_ASAP7_75t_L g3115 ( 
.A(n_2633),
.Y(n_3115)
);

INVx4_ASAP7_75t_SL g3116 ( 
.A(n_2710),
.Y(n_3116)
);

NOR2xp33_ASAP7_75t_L g3117 ( 
.A(n_2689),
.B(n_1542),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2592),
.B(n_1543),
.Y(n_3118)
);

OR2x6_ASAP7_75t_L g3119 ( 
.A(n_2491),
.B(n_2663),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2635),
.Y(n_3120)
);

OR2x2_ASAP7_75t_L g3121 ( 
.A(n_2690),
.B(n_1546),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2707),
.Y(n_3122)
);

INVx3_ASAP7_75t_L g3123 ( 
.A(n_2636),
.Y(n_3123)
);

BUFx6f_ASAP7_75t_L g3124 ( 
.A(n_2709),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2500),
.B(n_1547),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2717),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2356),
.Y(n_3127)
);

BUFx3_ASAP7_75t_L g3128 ( 
.A(n_2667),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2362),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2719),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2526),
.B(n_1548),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2364),
.Y(n_3132)
);

BUFx6f_ASAP7_75t_L g3133 ( 
.A(n_2729),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_2679),
.B(n_1549),
.Y(n_3134)
);

AND2x4_ASAP7_75t_L g3135 ( 
.A(n_2631),
.B(n_1526),
.Y(n_3135)
);

BUFx6f_ASAP7_75t_L g3136 ( 
.A(n_2732),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2682),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2664),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2485),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2632),
.B(n_1550),
.Y(n_3140)
);

INVx4_ASAP7_75t_L g3141 ( 
.A(n_2710),
.Y(n_3141)
);

HB1xp67_ASAP7_75t_L g3142 ( 
.A(n_2603),
.Y(n_3142)
);

OAI21xp33_ASAP7_75t_L g3143 ( 
.A1(n_2641),
.A2(n_1557),
.B(n_1555),
.Y(n_3143)
);

INVx8_ASAP7_75t_L g3144 ( 
.A(n_2517),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2733),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2492),
.Y(n_3146)
);

CKINVDCx5p33_ASAP7_75t_R g3147 ( 
.A(n_2671),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2492),
.Y(n_3148)
);

BUFx6f_ASAP7_75t_L g3149 ( 
.A(n_2672),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2531),
.Y(n_3150)
);

XOR2xp5_ASAP7_75t_L g3151 ( 
.A(n_2602),
.B(n_1559),
.Y(n_3151)
);

AND2x6_ASAP7_75t_L g3152 ( 
.A(n_2538),
.B(n_1051),
.Y(n_3152)
);

INVx6_ASAP7_75t_L g3153 ( 
.A(n_2675),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2542),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2394),
.Y(n_3155)
);

INVx3_ASAP7_75t_L g3156 ( 
.A(n_2680),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2403),
.B(n_1561),
.Y(n_3157)
);

AOI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_2530),
.A2(n_1565),
.B1(n_1566),
.B2(n_1562),
.Y(n_3158)
);

OAI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_2684),
.A2(n_1573),
.B1(n_1578),
.B2(n_1567),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2404),
.Y(n_3160)
);

BUFx2_ASAP7_75t_L g3161 ( 
.A(n_2664),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2376),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_2511),
.B(n_1582),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2535),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2503),
.B(n_1584),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_2512),
.B(n_1585),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2622),
.Y(n_3167)
);

NAND2x1p5_ASAP7_75t_L g3168 ( 
.A(n_2674),
.B(n_1105),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2541),
.Y(n_3169)
);

INVx2_ASAP7_75t_L g3170 ( 
.A(n_2623),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2572),
.B(n_1586),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2627),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2484),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2674),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_SL g3175 ( 
.A(n_2660),
.B(n_1587),
.Y(n_3175)
);

NAND2x1p5_ASAP7_75t_L g3176 ( 
.A(n_2678),
.B(n_1051),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_2496),
.A2(n_2624),
.B1(n_2534),
.B2(n_2678),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2644),
.Y(n_3178)
);

INVx1_ASAP7_75t_SL g3179 ( 
.A(n_2634),
.Y(n_3179)
);

INVx3_ASAP7_75t_L g3180 ( 
.A(n_2685),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2649),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2654),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2655),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2563),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2437),
.B(n_1588),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2440),
.Y(n_3186)
);

OR2x2_ASAP7_75t_L g3187 ( 
.A(n_2540),
.B(n_1592),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2448),
.Y(n_3188)
);

AND2x6_ASAP7_75t_L g3189 ( 
.A(n_2558),
.B(n_1051),
.Y(n_3189)
);

INVx4_ASAP7_75t_L g3190 ( 
.A(n_2621),
.Y(n_3190)
);

OR2x2_ASAP7_75t_L g3191 ( 
.A(n_2735),
.B(n_1593),
.Y(n_3191)
);

INVx3_ASAP7_75t_L g3192 ( 
.A(n_2466),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2449),
.B(n_1594),
.Y(n_3193)
);

BUFx6f_ASAP7_75t_L g3194 ( 
.A(n_2569),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2345),
.B(n_1596),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2694),
.Y(n_3196)
);

BUFx4f_ASAP7_75t_L g3197 ( 
.A(n_2522),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2697),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2711),
.B(n_1597),
.Y(n_3199)
);

AOI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2666),
.A2(n_1599),
.B1(n_1600),
.B2(n_1598),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2658),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2343),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2352),
.Y(n_3203)
);

HB1xp67_ASAP7_75t_L g3204 ( 
.A(n_2381),
.Y(n_3204)
);

INVxp67_ASAP7_75t_SL g3205 ( 
.A(n_2698),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_2389),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2352),
.Y(n_3207)
);

AND2x4_ASAP7_75t_L g3208 ( 
.A(n_2586),
.B(n_1533),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_2348),
.B(n_1602),
.Y(n_3209)
);

INVx4_ASAP7_75t_L g3210 ( 
.A(n_2380),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2343),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_2453),
.B(n_1603),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_2698),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2343),
.Y(n_3214)
);

INVx2_ASAP7_75t_SL g3215 ( 
.A(n_2380),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2343),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_2586),
.B(n_1544),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_2369),
.B(n_1604),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2343),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2586),
.B(n_1605),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2586),
.B(n_1607),
.Y(n_3221)
);

OR2x6_ASAP7_75t_L g3222 ( 
.A(n_2380),
.B(n_1262),
.Y(n_3222)
);

BUFx4f_ASAP7_75t_L g3223 ( 
.A(n_2389),
.Y(n_3223)
);

OR2x2_ASAP7_75t_L g3224 ( 
.A(n_2453),
.B(n_1611),
.Y(n_3224)
);

INVx1_ASAP7_75t_SL g3225 ( 
.A(n_2381),
.Y(n_3225)
);

BUFx10_ASAP7_75t_L g3226 ( 
.A(n_2639),
.Y(n_3226)
);

HB1xp67_ASAP7_75t_L g3227 ( 
.A(n_2381),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2343),
.Y(n_3228)
);

INVx1_ASAP7_75t_SL g3229 ( 
.A(n_2381),
.Y(n_3229)
);

NOR2xp33_ASAP7_75t_L g3230 ( 
.A(n_2438),
.B(n_1612),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2348),
.B(n_1613),
.Y(n_3231)
);

INVx4_ASAP7_75t_L g3232 ( 
.A(n_2380),
.Y(n_3232)
);

BUFx4f_ASAP7_75t_L g3233 ( 
.A(n_2389),
.Y(n_3233)
);

OR2x2_ASAP7_75t_L g3234 ( 
.A(n_2453),
.B(n_1616),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_2438),
.B(n_1618),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2352),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2343),
.Y(n_3237)
);

OR2x2_ASAP7_75t_L g3238 ( 
.A(n_2453),
.B(n_1621),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2586),
.B(n_1622),
.Y(n_3239)
);

INVx2_ASAP7_75t_SL g3240 ( 
.A(n_2380),
.Y(n_3240)
);

AND2x2_ASAP7_75t_L g3241 ( 
.A(n_2369),
.B(n_1625),
.Y(n_3241)
);

AND2x6_ASAP7_75t_L g3242 ( 
.A(n_2698),
.B(n_1071),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_2543),
.Y(n_3243)
);

OR2x2_ASAP7_75t_L g3244 ( 
.A(n_2453),
.B(n_1628),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2586),
.B(n_1639),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2343),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2343),
.Y(n_3247)
);

INVx4_ASAP7_75t_L g3248 ( 
.A(n_2380),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_2586),
.B(n_1552),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2352),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2586),
.B(n_1642),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2586),
.B(n_1643),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2369),
.B(n_1644),
.Y(n_3253)
);

OR2x2_ASAP7_75t_L g3254 ( 
.A(n_2453),
.B(n_1649),
.Y(n_3254)
);

BUFx2_ASAP7_75t_L g3255 ( 
.A(n_2381),
.Y(n_3255)
);

INVx1_ASAP7_75t_SL g3256 ( 
.A(n_2381),
.Y(n_3256)
);

HB1xp67_ASAP7_75t_L g3257 ( 
.A(n_2381),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2343),
.Y(n_3258)
);

INVx4_ASAP7_75t_SL g3259 ( 
.A(n_2368),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_2543),
.Y(n_3260)
);

BUFx10_ASAP7_75t_L g3261 ( 
.A(n_2639),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2369),
.B(n_1650),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2369),
.B(n_1651),
.Y(n_3263)
);

INVx4_ASAP7_75t_L g3264 ( 
.A(n_2380),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2352),
.Y(n_3265)
);

INVx4_ASAP7_75t_L g3266 ( 
.A(n_2380),
.Y(n_3266)
);

BUFx8_ASAP7_75t_SL g3267 ( 
.A(n_2701),
.Y(n_3267)
);

INVx4_ASAP7_75t_L g3268 ( 
.A(n_2380),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_2352),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_2586),
.B(n_1554),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2452),
.Y(n_3271)
);

BUFx3_ASAP7_75t_L g3272 ( 
.A(n_2380),
.Y(n_3272)
);

AND2x6_ASAP7_75t_L g3273 ( 
.A(n_2698),
.B(n_1071),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_2453),
.B(n_1652),
.Y(n_3274)
);

INVx3_ASAP7_75t_L g3275 ( 
.A(n_2698),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_2381),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2352),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_2389),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_2389),
.Y(n_3279)
);

CKINVDCx16_ASAP7_75t_R g3280 ( 
.A(n_2479),
.Y(n_3280)
);

INVx4_ASAP7_75t_L g3281 ( 
.A(n_2380),
.Y(n_3281)
);

INVx6_ASAP7_75t_L g3282 ( 
.A(n_2454),
.Y(n_3282)
);

OR2x2_ASAP7_75t_L g3283 ( 
.A(n_2453),
.B(n_1654),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_2352),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2352),
.Y(n_3285)
);

CKINVDCx20_ASAP7_75t_R g3286 ( 
.A(n_2564),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_2438),
.B(n_1656),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2438),
.B(n_1658),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_2369),
.B(n_1660),
.Y(n_3289)
);

AND2x6_ASAP7_75t_L g3290 ( 
.A(n_2698),
.B(n_1071),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_SL g3291 ( 
.A(n_2348),
.B(n_1662),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_2460),
.A2(n_1663),
.B1(n_1038),
.B2(n_1039),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2343),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2343),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_2348),
.B(n_1034),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_2352),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2343),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2343),
.Y(n_3298)
);

NOR2xp33_ASAP7_75t_L g3299 ( 
.A(n_2438),
.B(n_1053),
.Y(n_3299)
);

BUFx6f_ASAP7_75t_L g3300 ( 
.A(n_2543),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_2352),
.Y(n_3301)
);

INVx4_ASAP7_75t_L g3302 ( 
.A(n_2380),
.Y(n_3302)
);

OR2x6_ASAP7_75t_L g3303 ( 
.A(n_2380),
.B(n_1262),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2343),
.Y(n_3304)
);

AND2x4_ASAP7_75t_SL g3305 ( 
.A(n_2564),
.B(n_1071),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2343),
.Y(n_3306)
);

HB1xp67_ASAP7_75t_L g3307 ( 
.A(n_2381),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2586),
.B(n_1453),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2343),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_2369),
.B(n_1055),
.Y(n_3310)
);

INVx3_ASAP7_75t_L g3311 ( 
.A(n_2698),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_2438),
.B(n_1056),
.Y(n_3312)
);

BUFx3_ASAP7_75t_L g3313 ( 
.A(n_2380),
.Y(n_3313)
);

HB1xp67_ASAP7_75t_L g3314 ( 
.A(n_2381),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2343),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2352),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_2460),
.A2(n_1061),
.B1(n_1091),
.B2(n_1058),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2586),
.B(n_1454),
.Y(n_3318)
);

BUFx3_ASAP7_75t_L g3319 ( 
.A(n_2380),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_2352),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_2460),
.A2(n_1130),
.B1(n_1163),
.B2(n_1106),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2343),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_2438),
.B(n_1187),
.Y(n_3323)
);

NOR2x1p5_ASAP7_75t_L g3324 ( 
.A(n_2389),
.B(n_1214),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_2438),
.B(n_1254),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_2352),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2352),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2586),
.B(n_1468),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_2369),
.B(n_1269),
.Y(n_3329)
);

OAI21xp33_ASAP7_75t_SL g3330 ( 
.A1(n_2481),
.A2(n_1653),
.B(n_1647),
.Y(n_3330)
);

AND2x6_ASAP7_75t_L g3331 ( 
.A(n_2698),
.B(n_1144),
.Y(n_3331)
);

INVx2_ASAP7_75t_SL g3332 ( 
.A(n_2380),
.Y(n_3332)
);

BUFx2_ASAP7_75t_L g3333 ( 
.A(n_2381),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_2343),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2586),
.B(n_1472),
.Y(n_3335)
);

AOI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_2350),
.A2(n_1299),
.B1(n_1304),
.B2(n_1298),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_2438),
.B(n_1312),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2343),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_2698),
.Y(n_3339)
);

CKINVDCx5p33_ASAP7_75t_R g3340 ( 
.A(n_2389),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2352),
.Y(n_3341)
);

AND2x4_ASAP7_75t_L g3342 ( 
.A(n_2586),
.B(n_1576),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2452),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_2352),
.Y(n_3344)
);

BUFx10_ASAP7_75t_L g3345 ( 
.A(n_2639),
.Y(n_3345)
);

CKINVDCx20_ASAP7_75t_R g3346 ( 
.A(n_2564),
.Y(n_3346)
);

BUFx3_ASAP7_75t_L g3347 ( 
.A(n_2380),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2352),
.Y(n_3348)
);

INVx4_ASAP7_75t_L g3349 ( 
.A(n_2380),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_2352),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_2343),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2586),
.B(n_1475),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_2438),
.B(n_1316),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2352),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2343),
.Y(n_3355)
);

BUFx6f_ASAP7_75t_L g3356 ( 
.A(n_2543),
.Y(n_3356)
);

AND2x4_ASAP7_75t_L g3357 ( 
.A(n_2586),
.B(n_1632),
.Y(n_3357)
);

INVx4_ASAP7_75t_L g3358 ( 
.A(n_2380),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_2348),
.B(n_1657),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_2698),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2343),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_2460),
.A2(n_1347),
.B1(n_1349),
.B2(n_1345),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2343),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_2389),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_2348),
.B(n_1666),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_2586),
.B(n_1664),
.Y(n_3366)
);

BUFx2_ASAP7_75t_L g3367 ( 
.A(n_2381),
.Y(n_3367)
);

AND2x4_ASAP7_75t_L g3368 ( 
.A(n_2586),
.B(n_1479),
.Y(n_3368)
);

INVx4_ASAP7_75t_L g3369 ( 
.A(n_2380),
.Y(n_3369)
);

BUFx4f_ASAP7_75t_L g3370 ( 
.A(n_2389),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2352),
.Y(n_3371)
);

NAND3x1_ASAP7_75t_L g3372 ( 
.A(n_2731),
.B(n_1483),
.C(n_1482),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2352),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2352),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2452),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_2369),
.B(n_1352),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_2352),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_2348),
.B(n_1378),
.Y(n_3378)
);

INVx4_ASAP7_75t_SL g3379 ( 
.A(n_2368),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2452),
.Y(n_3380)
);

INVx4_ASAP7_75t_L g3381 ( 
.A(n_2380),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_2380),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2452),
.Y(n_3383)
);

NAND2x1p5_ASAP7_75t_L g3384 ( 
.A(n_2683),
.B(n_1144),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_L g3385 ( 
.A(n_2438),
.B(n_1384),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_2586),
.B(n_1486),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2343),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2586),
.B(n_1487),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_2586),
.B(n_1492),
.Y(n_3389)
);

INVx3_ASAP7_75t_L g3390 ( 
.A(n_2698),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2586),
.B(n_1500),
.Y(n_3391)
);

INVxp67_ASAP7_75t_L g3392 ( 
.A(n_2381),
.Y(n_3392)
);

INVx2_ASAP7_75t_SL g3393 ( 
.A(n_2380),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_2352),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_2369),
.B(n_1391),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_2740),
.B(n_1398),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3218),
.B(n_1401),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3280),
.B(n_1638),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3368),
.B(n_3386),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_SL g3400 ( 
.A(n_2928),
.B(n_1667),
.Y(n_3400)
);

OAI221xp5_ASAP7_75t_L g3401 ( 
.A1(n_2769),
.A2(n_1422),
.B1(n_1473),
.B2(n_1423),
.C(n_1411),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_SL g3402 ( 
.A(n_2928),
.B(n_1498),
.Y(n_3402)
);

O2A1O1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_2989),
.A2(n_1534),
.B(n_1541),
.C(n_1527),
.Y(n_3403)
);

AND2x6_ASAP7_75t_L g3404 ( 
.A(n_2805),
.B(n_1144),
.Y(n_3404)
);

NOR3xp33_ASAP7_75t_L g3405 ( 
.A(n_2898),
.B(n_1560),
.C(n_1558),
.Y(n_3405)
);

BUFx5_ASAP7_75t_L g3406 ( 
.A(n_3242),
.Y(n_3406)
);

OR2x2_ASAP7_75t_L g3407 ( 
.A(n_2986),
.B(n_1508),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3368),
.B(n_1570),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3386),
.B(n_3389),
.Y(n_3409)
);

INVx2_ASAP7_75t_SL g3410 ( 
.A(n_2759),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_2797),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3241),
.B(n_1510),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3389),
.B(n_1572),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3253),
.B(n_1521),
.Y(n_3414)
);

BUFx12f_ASAP7_75t_L g3415 ( 
.A(n_2892),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_2808),
.Y(n_3416)
);

AOI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_2970),
.A2(n_2842),
.B1(n_2895),
.B2(n_2916),
.Y(n_3417)
);

NAND2x1_ASAP7_75t_L g3418 ( 
.A(n_3242),
.B(n_1637),
.Y(n_3418)
);

NOR3xp33_ASAP7_75t_L g3419 ( 
.A(n_2779),
.B(n_1595),
.C(n_1575),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3208),
.B(n_1601),
.Y(n_3420)
);

NAND2xp33_ASAP7_75t_L g3421 ( 
.A(n_3152),
.B(n_1524),
.Y(n_3421)
);

INVx2_ASAP7_75t_SL g3422 ( 
.A(n_2759),
.Y(n_3422)
);

O2A1O1Ixp33_ASAP7_75t_L g3423 ( 
.A1(n_3025),
.A2(n_2947),
.B(n_2794),
.C(n_2908),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_2811),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_2745),
.B(n_1529),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_3330),
.A2(n_1255),
.B(n_1265),
.C(n_1248),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3061),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3208),
.B(n_1606),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2835),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3217),
.B(n_1610),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_2958),
.B(n_1538),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_2857),
.A2(n_1577),
.B1(n_1580),
.B2(n_1551),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2865),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_2884),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_SL g3435 ( 
.A(n_3225),
.B(n_1626),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2868),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3229),
.B(n_1629),
.Y(n_3437)
);

OR2x6_ASAP7_75t_L g3438 ( 
.A(n_2761),
.B(n_1356),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2877),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3146),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3217),
.B(n_1620),
.Y(n_3441)
);

NAND2xp33_ASAP7_75t_L g3442 ( 
.A(n_3152),
.B(n_1583),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3249),
.B(n_1627),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3249),
.B(n_1635),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_2887),
.Y(n_3445)
);

INVx5_ASAP7_75t_L g3446 ( 
.A(n_2761),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3148),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3270),
.B(n_1636),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3270),
.B(n_1640),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3342),
.B(n_1641),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_2784),
.B(n_1609),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_2976),
.A2(n_1624),
.B1(n_1630),
.B2(n_1617),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_3256),
.B(n_1144),
.Y(n_3453)
);

NAND2xp33_ASAP7_75t_SL g3454 ( 
.A(n_3053),
.B(n_3088),
.Y(n_3454)
);

INVx3_ASAP7_75t_L g3455 ( 
.A(n_2805),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_2907),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_2736),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3262),
.B(n_1645),
.Y(n_3458)
);

AND2x6_ASAP7_75t_SL g3459 ( 
.A(n_3086),
.B(n_1661),
.Y(n_3459)
);

AOI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_2976),
.A2(n_1255),
.B1(n_1265),
.B2(n_1248),
.Y(n_3460)
);

NAND2xp33_ASAP7_75t_L g3461 ( 
.A(n_3152),
.B(n_1147),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3342),
.B(n_1356),
.Y(n_3462)
);

O2A1O1Ixp33_ASAP7_75t_L g3463 ( 
.A1(n_2816),
.A2(n_1464),
.B(n_1287),
.C(n_1317),
.Y(n_3463)
);

INVx2_ASAP7_75t_SL g3464 ( 
.A(n_2759),
.Y(n_3464)
);

NOR2xp67_ASAP7_75t_L g3465 ( 
.A(n_3154),
.B(n_2),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_2926),
.B(n_1147),
.Y(n_3466)
);

NAND3xp33_ASAP7_75t_L g3467 ( 
.A(n_2941),
.B(n_3235),
.C(n_3230),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3357),
.B(n_1464),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3357),
.B(n_1277),
.Y(n_3469)
);

NOR2xp33_ASAP7_75t_L g3470 ( 
.A(n_3018),
.B(n_1277),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3255),
.B(n_1147),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3366),
.B(n_1287),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3366),
.B(n_1317),
.Y(n_3473)
);

INVx3_ASAP7_75t_L g3474 ( 
.A(n_2805),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_2772),
.B(n_1360),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3154),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3150),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_2772),
.B(n_1360),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3150),
.Y(n_3479)
);

INVxp67_ASAP7_75t_SL g3480 ( 
.A(n_3204),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2737),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3263),
.B(n_1377),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3164),
.Y(n_3483)
);

OAI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2937),
.A2(n_1385),
.B(n_1377),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3164),
.Y(n_3485)
);

O2A1O1Ixp5_ASAP7_75t_L g3486 ( 
.A1(n_3190),
.A2(n_3197),
.B(n_3184),
.C(n_3155),
.Y(n_3486)
);

AND2x4_ASAP7_75t_L g3487 ( 
.A(n_2903),
.B(n_1385),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_2777),
.B(n_2778),
.Y(n_3488)
);

NAND2xp33_ASAP7_75t_SL g3489 ( 
.A(n_2791),
.B(n_1395),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2777),
.B(n_1395),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_2778),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_SL g3492 ( 
.A(n_3333),
.B(n_3367),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_2972),
.A2(n_1191),
.B1(n_1429),
.B2(n_1147),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_2843),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_2826),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_2826),
.B(n_1420),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_L g3497 ( 
.A(n_2841),
.B(n_1420),
.Y(n_3497)
);

INVx2_ASAP7_75t_L g3498 ( 
.A(n_3271),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3271),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3343),
.Y(n_3500)
);

INVxp67_ASAP7_75t_L g3501 ( 
.A(n_3227),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3343),
.B(n_1539),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_2936),
.B(n_2942),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3287),
.B(n_1539),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3375),
.B(n_3380),
.Y(n_3505)
);

AOI22xp33_ASAP7_75t_L g3506 ( 
.A1(n_3042),
.A2(n_1429),
.B1(n_1434),
.B2(n_1191),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3375),
.Y(n_3507)
);

INVx3_ASAP7_75t_L g3508 ( 
.A(n_2774),
.Y(n_3508)
);

INVx5_ASAP7_75t_L g3509 ( 
.A(n_3242),
.Y(n_3509)
);

INVxp67_ASAP7_75t_L g3510 ( 
.A(n_3257),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3380),
.B(n_1563),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_2847),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3383),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_SL g3514 ( 
.A(n_3090),
.B(n_1191),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_2848),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3288),
.B(n_1563),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3383),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_2918),
.B(n_1569),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_2855),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_2878),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_2994),
.B(n_1569),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2995),
.B(n_1619),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_2934),
.B(n_1619),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_3212),
.B(n_1631),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3224),
.B(n_1631),
.Y(n_3525)
);

INVx2_ASAP7_75t_SL g3526 ( 
.A(n_3305),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_2792),
.B(n_1648),
.Y(n_3527)
);

INVxp67_ASAP7_75t_SL g3528 ( 
.A(n_3276),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_L g3529 ( 
.A(n_3234),
.B(n_1648),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2856),
.Y(n_3530)
);

AOI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3019),
.A2(n_1659),
.B1(n_1429),
.B2(n_1434),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2798),
.B(n_1659),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_L g3533 ( 
.A(n_3238),
.B(n_0),
.Y(n_3533)
);

NAND2x1p5_ASAP7_75t_L g3534 ( 
.A(n_3210),
.B(n_3232),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_3244),
.B(n_3254),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_L g3536 ( 
.A(n_3274),
.B(n_2),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_2741),
.B(n_1191),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_2741),
.B(n_1429),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_2799),
.B(n_3),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2861),
.Y(n_3540)
);

INVx1_ASAP7_75t_SL g3541 ( 
.A(n_3286),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_2801),
.B(n_2806),
.Y(n_3542)
);

AOI22xp33_ASAP7_75t_L g3543 ( 
.A1(n_3003),
.A2(n_1484),
.B1(n_1512),
.B2(n_1434),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_2809),
.B(n_3),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_2746),
.Y(n_3545)
);

AND2x4_ASAP7_75t_L g3546 ( 
.A(n_2903),
.B(n_4),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_2753),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3289),
.A2(n_1484),
.B1(n_1512),
.B2(n_1434),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_SL g3549 ( 
.A(n_2741),
.B(n_1484),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2810),
.B(n_5),
.Y(n_3550)
);

AOI22x1_ASAP7_75t_L g3551 ( 
.A1(n_3019),
.A2(n_1484),
.B1(n_1646),
.B2(n_1512),
.Y(n_3551)
);

OAI21xp33_ASAP7_75t_L g3552 ( 
.A1(n_3040),
.A2(n_1646),
.B(n_1512),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_2814),
.B(n_5),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_2742),
.B(n_1646),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_2875),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_2818),
.B(n_5),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_2766),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_2822),
.B(n_6),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_2828),
.Y(n_3559)
);

AND2x2_ASAP7_75t_SL g3560 ( 
.A(n_3223),
.B(n_1457),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_2834),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_2823),
.B(n_6),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_2757),
.B(n_6),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_2824),
.B(n_7),
.Y(n_3564)
);

INVx5_ASAP7_75t_L g3565 ( 
.A(n_3242),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2885),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_2836),
.Y(n_3567)
);

BUFx3_ASAP7_75t_L g3568 ( 
.A(n_3346),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_2896),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_2825),
.B(n_7),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_2901),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2904),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3202),
.B(n_8),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3211),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3214),
.B(n_8),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3216),
.B(n_3219),
.Y(n_3576)
);

OR2x6_ASAP7_75t_L g3577 ( 
.A(n_3144),
.B(n_1646),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_L g3578 ( 
.A(n_3283),
.B(n_8),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_2742),
.B(n_2763),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3228),
.B(n_9),
.Y(n_3580)
);

NOR2xp67_ASAP7_75t_L g3581 ( 
.A(n_2774),
.B(n_10),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_L g3582 ( 
.A(n_3392),
.B(n_9),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3237),
.B(n_9),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_SL g3584 ( 
.A(n_2742),
.B(n_889),
.Y(n_3584)
);

AOI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3020),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3246),
.B(n_10),
.Y(n_3586)
);

AOI22xp33_ASAP7_75t_L g3587 ( 
.A1(n_3086),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_3587)
);

OAI22xp5_ASAP7_75t_SL g3588 ( 
.A1(n_2839),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_3588)
);

AND2x4_ASAP7_75t_L g3589 ( 
.A(n_2903),
.B(n_14),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3247),
.B(n_14),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_SL g3591 ( 
.A(n_2750),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3258),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3293),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3294),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3299),
.B(n_15),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2840),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3297),
.B(n_16),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3298),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3304),
.B(n_16),
.Y(n_3599)
);

NOR2xp67_ASAP7_75t_L g3600 ( 
.A(n_2780),
.B(n_18),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_3312),
.B(n_17),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3306),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3309),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3315),
.B(n_17),
.Y(n_3604)
);

INVx8_ASAP7_75t_L g3605 ( 
.A(n_3144),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3322),
.B(n_3334),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_SL g3607 ( 
.A(n_2763),
.B(n_889),
.Y(n_3607)
);

BUFx4f_ASAP7_75t_L g3608 ( 
.A(n_3107),
.Y(n_3608)
);

AOI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_2882),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3338),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3351),
.B(n_20),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3355),
.B(n_3361),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3363),
.B(n_20),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3387),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_SL g3615 ( 
.A(n_2763),
.B(n_890),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_2859),
.Y(n_3616)
);

INVx3_ASAP7_75t_L g3617 ( 
.A(n_2780),
.Y(n_3617)
);

INVx2_ASAP7_75t_SL g3618 ( 
.A(n_2793),
.Y(n_3618)
);

AOI22xp5_ASAP7_75t_L g3619 ( 
.A1(n_3040),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3323),
.B(n_22),
.Y(n_3620)
);

BUFx2_ASAP7_75t_L g3621 ( 
.A(n_3307),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_SL g3622 ( 
.A(n_2770),
.B(n_890),
.Y(n_3622)
);

NAND2xp33_ASAP7_75t_L g3623 ( 
.A(n_3152),
.B(n_22),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3203),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_L g3625 ( 
.A(n_3325),
.B(n_24),
.Y(n_3625)
);

INVxp67_ASAP7_75t_L g3626 ( 
.A(n_3314),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_2739),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_L g3628 ( 
.A(n_3337),
.B(n_3353),
.Y(n_3628)
);

O2A1O1Ixp33_ASAP7_75t_L g3629 ( 
.A1(n_3017),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_2770),
.B(n_891),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_SL g3631 ( 
.A(n_2770),
.B(n_892),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_2743),
.Y(n_3632)
);

BUFx3_ASAP7_75t_L g3633 ( 
.A(n_2756),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3207),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3236),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_2751),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_2785),
.B(n_893),
.Y(n_3637)
);

AOI22xp5_ASAP7_75t_L g3638 ( 
.A1(n_3372),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_SL g3639 ( 
.A(n_2785),
.B(n_893),
.Y(n_3639)
);

BUFx6f_ASAP7_75t_L g3640 ( 
.A(n_2785),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_2844),
.B(n_25),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3250),
.Y(n_3642)
);

NOR2xp33_ASAP7_75t_L g3643 ( 
.A(n_3385),
.B(n_2919),
.Y(n_3643)
);

OAI21xp33_ASAP7_75t_L g3644 ( 
.A1(n_2795),
.A2(n_26),
.B(n_27),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_L g3645 ( 
.A1(n_2790),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_3645)
);

BUFx6f_ASAP7_75t_L g3646 ( 
.A(n_3243),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3243),
.B(n_894),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_2879),
.B(n_28),
.Y(n_3648)
);

NAND2xp33_ASAP7_75t_L g3649 ( 
.A(n_3110),
.B(n_28),
.Y(n_3649)
);

O2A1O1Ixp5_ASAP7_75t_L g3650 ( 
.A1(n_3190),
.A2(n_3197),
.B(n_3155),
.C(n_3160),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_2767),
.B(n_29),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_2867),
.B(n_29),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_L g3653 ( 
.A(n_3006),
.B(n_30),
.Y(n_3653)
);

INVx3_ASAP7_75t_L g3654 ( 
.A(n_2775),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_2846),
.B(n_30),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3310),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_3656)
);

INVx8_ASAP7_75t_L g3657 ( 
.A(n_2911),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_2775),
.Y(n_3658)
);

NOR2xp33_ASAP7_75t_L g3659 ( 
.A(n_3179),
.B(n_2983),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_2755),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3058),
.B(n_32),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3076),
.B(n_32),
.Y(n_3662)
);

OR2x6_ASAP7_75t_L g3663 ( 
.A(n_2749),
.B(n_33),
.Y(n_3663)
);

AOI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_3038),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3014),
.B(n_34),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3265),
.Y(n_3666)
);

A2O1A1Ixp33_ASAP7_75t_L g3667 ( 
.A1(n_3082),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3329),
.B(n_35),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_2789),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3376),
.B(n_36),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3395),
.B(n_36),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3269),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3277),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3043),
.B(n_37),
.Y(n_3674)
);

BUFx3_ASAP7_75t_L g3675 ( 
.A(n_3272),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3284),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3243),
.B(n_894),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_SL g3678 ( 
.A(n_3260),
.B(n_895),
.Y(n_3678)
);

NAND2xp33_ASAP7_75t_L g3679 ( 
.A(n_3110),
.B(n_38),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_2988),
.B(n_3125),
.Y(n_3680)
);

BUFx6f_ASAP7_75t_L g3681 ( 
.A(n_3260),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_2997),
.B(n_38),
.Y(n_3682)
);

O2A1O1Ixp33_ASAP7_75t_L g3683 ( 
.A1(n_3011),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_2788),
.B(n_39),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3059),
.B(n_39),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_2893),
.B(n_40),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3023),
.B(n_40),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_2910),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_2881),
.B(n_41),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_2949),
.B(n_41),
.Y(n_3690)
);

NAND3xp33_ASAP7_75t_L g3691 ( 
.A(n_3177),
.B(n_41),
.C(n_42),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3285),
.Y(n_3692)
);

NOR2xp67_ASAP7_75t_L g3693 ( 
.A(n_2962),
.B(n_43),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_2966),
.B(n_42),
.Y(n_3694)
);

A2O1A1Ixp33_ASAP7_75t_L g3695 ( 
.A1(n_2888),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_3695)
);

INVx2_ASAP7_75t_SL g3696 ( 
.A(n_2793),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_2952),
.B(n_43),
.Y(n_3697)
);

OAI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_2953),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_SL g3699 ( 
.A(n_3260),
.B(n_896),
.Y(n_3699)
);

O2A1O1Ixp33_ASAP7_75t_L g3700 ( 
.A1(n_3111),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3296),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_2849),
.B(n_46),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_2869),
.B(n_47),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3301),
.Y(n_3704)
);

OR2x2_ASAP7_75t_L g3705 ( 
.A(n_2985),
.B(n_47),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3316),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_SL g3707 ( 
.A(n_3300),
.B(n_896),
.Y(n_3707)
);

INVx2_ASAP7_75t_SL g3708 ( 
.A(n_3282),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_3300),
.B(n_897),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_3300),
.B(n_897),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_2869),
.B(n_47),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3320),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_2880),
.B(n_48),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3326),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_2758),
.B(n_2956),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_2880),
.B(n_48),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3327),
.Y(n_3717)
);

AOI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3135),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3056),
.B(n_49),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_SL g3720 ( 
.A(n_3356),
.B(n_2911),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3135),
.B(n_3117),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3341),
.Y(n_3722)
);

BUFx3_ASAP7_75t_L g3723 ( 
.A(n_3313),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_L g3724 ( 
.A(n_3063),
.B(n_49),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3344),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_L g3726 ( 
.A(n_2906),
.B(n_50),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3356),
.B(n_898),
.Y(n_3727)
);

INVx2_ASAP7_75t_SL g3728 ( 
.A(n_3282),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_2886),
.B(n_50),
.Y(n_3729)
);

INVx2_ASAP7_75t_SL g3730 ( 
.A(n_2750),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3356),
.B(n_898),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_2860),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3348),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3308),
.B(n_3318),
.Y(n_3734)
);

INVx2_ASAP7_75t_SL g3735 ( 
.A(n_2838),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3328),
.B(n_51),
.Y(n_3736)
);

OAI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3335),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_3737)
);

AOI22xp5_ASAP7_75t_L g3738 ( 
.A1(n_2860),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3352),
.B(n_54),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_2754),
.B(n_3209),
.Y(n_3740)
);

NAND3xp33_ASAP7_75t_L g3741 ( 
.A(n_2923),
.B(n_55),
.C(n_56),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3388),
.B(n_55),
.Y(n_3742)
);

NOR2xp33_ASAP7_75t_L g3743 ( 
.A(n_3231),
.B(n_56),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3350),
.Y(n_3744)
);

OR2x2_ASAP7_75t_L g3745 ( 
.A(n_3035),
.B(n_56),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3354),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3371),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3373),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_2953),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3374),
.Y(n_3750)
);

NOR2xp33_ASAP7_75t_L g3751 ( 
.A(n_3291),
.B(n_57),
.Y(n_3751)
);

INVx2_ASAP7_75t_SL g3752 ( 
.A(n_2838),
.Y(n_3752)
);

OR2x6_ASAP7_75t_L g3753 ( 
.A(n_2749),
.B(n_3222),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3377),
.Y(n_3754)
);

INVx2_ASAP7_75t_SL g3755 ( 
.A(n_3226),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3391),
.B(n_58),
.Y(n_3756)
);

AOI22xp33_ASAP7_75t_L g3757 ( 
.A1(n_2979),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_2864),
.B(n_60),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_2911),
.B(n_899),
.Y(n_3759)
);

OAI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_2914),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3394),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_2955),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_2940),
.B(n_61),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_R g3764 ( 
.A(n_3048),
.B(n_3206),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_2959),
.Y(n_3765)
);

NOR2x1p5_ASAP7_75t_L g3766 ( 
.A(n_3278),
.B(n_3279),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_2900),
.B(n_61),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3139),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_2944),
.B(n_62),
.Y(n_3769)
);

NOR2xp33_ASAP7_75t_L g3770 ( 
.A(n_3121),
.B(n_62),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3168),
.B(n_63),
.Y(n_3771)
);

O2A1O1Ixp33_ASAP7_75t_L g3772 ( 
.A1(n_3118),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_2964),
.Y(n_3773)
);

INVxp33_ASAP7_75t_L g3774 ( 
.A(n_2830),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_2946),
.B(n_64),
.Y(n_3775)
);

NOR2xp33_ASAP7_75t_L g3776 ( 
.A(n_3091),
.B(n_64),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_2748),
.B(n_65),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3139),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3220),
.B(n_65),
.Y(n_3779)
);

NAND3xp33_ASAP7_75t_L g3780 ( 
.A(n_3033),
.B(n_66),
.C(n_67),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_2913),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3221),
.B(n_66),
.Y(n_3782)
);

XNOR2xp5_ASAP7_75t_L g3783 ( 
.A(n_3324),
.B(n_66),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_SL g3784 ( 
.A(n_3049),
.B(n_900),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_2979),
.B(n_68),
.Y(n_3785)
);

NAND2x1p5_ASAP7_75t_L g3786 ( 
.A(n_3210),
.B(n_69),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_2969),
.Y(n_3787)
);

OR2x6_ASAP7_75t_L g3788 ( 
.A(n_3222),
.B(n_3303),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_2765),
.B(n_69),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_2920),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_2921),
.Y(n_3791)
);

INVx4_ASAP7_75t_L g3792 ( 
.A(n_3232),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3239),
.B(n_69),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_2975),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_2980),
.Y(n_3795)
);

AOI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_2945),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3796)
);

INVxp67_ASAP7_75t_L g3797 ( 
.A(n_3004),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3081),
.Y(n_3798)
);

BUFx6f_ASAP7_75t_L g3799 ( 
.A(n_2820),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3245),
.B(n_70),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_SL g3801 ( 
.A(n_3049),
.B(n_900),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_2915),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3072),
.B(n_70),
.Y(n_3803)
);

AOI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3151),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3804)
);

NAND2xp33_ASAP7_75t_L g3805 ( 
.A(n_3110),
.B(n_71),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_2922),
.Y(n_3806)
);

INVx2_ASAP7_75t_L g3807 ( 
.A(n_2938),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3251),
.B(n_73),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3252),
.B(n_73),
.Y(n_3809)
);

OR2x2_ASAP7_75t_L g3810 ( 
.A(n_3050),
.B(n_74),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_3112),
.B(n_901),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_2990),
.B(n_74),
.Y(n_3812)
);

BUFx6f_ASAP7_75t_L g3813 ( 
.A(n_2820),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_2925),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_2951),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_SL g3816 ( 
.A(n_3112),
.B(n_901),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_2961),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_2930),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_L g3819 ( 
.A(n_3191),
.B(n_74),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3292),
.B(n_75),
.Y(n_3820)
);

AOI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_3089),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_3187),
.B(n_75),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_2948),
.B(n_2752),
.Y(n_3823)
);

AOI22xp33_ASAP7_75t_L g3824 ( 
.A1(n_3021),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_2948),
.B(n_78),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_2932),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_2762),
.B(n_78),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_3073),
.B(n_79),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_2962),
.B(n_902),
.Y(n_3829)
);

AOI22xp5_ASAP7_75t_L g3830 ( 
.A1(n_3143),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3830)
);

NOR2xp67_ASAP7_75t_SL g3831 ( 
.A(n_3340),
.B(n_79),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_SL g3832 ( 
.A(n_2962),
.B(n_902),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_2933),
.Y(n_3833)
);

NOR2xp67_ASAP7_75t_L g3834 ( 
.A(n_2776),
.B(n_82),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_2771),
.B(n_81),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3046),
.B(n_81),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_2796),
.B(n_82),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_2971),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_2791),
.B(n_2803),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_2802),
.B(n_83),
.Y(n_3840)
);

OR2x2_ASAP7_75t_L g3841 ( 
.A(n_3022),
.B(n_83),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_2982),
.Y(n_3842)
);

NOR2xp33_ASAP7_75t_L g3843 ( 
.A(n_3030),
.B(n_83),
.Y(n_3843)
);

HB1xp67_ASAP7_75t_L g3844 ( 
.A(n_3303),
.Y(n_3844)
);

NOR2xp33_ASAP7_75t_SL g3845 ( 
.A(n_3223),
.B(n_84),
.Y(n_3845)
);

OR2x2_ASAP7_75t_L g3846 ( 
.A(n_3026),
.B(n_2783),
.Y(n_3846)
);

NAND2xp33_ASAP7_75t_SL g3847 ( 
.A(n_2803),
.B(n_84),
.Y(n_3847)
);

INVx2_ASAP7_75t_SL g3848 ( 
.A(n_3226),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3027),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3039),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_2939),
.B(n_903),
.Y(n_3851)
);

NOR2xp67_ASAP7_75t_SL g3852 ( 
.A(n_3364),
.B(n_84),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3195),
.B(n_85),
.Y(n_3853)
);

AOI22xp33_ASAP7_75t_L g3854 ( 
.A1(n_2977),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_2804),
.B(n_86),
.Y(n_3855)
);

BUFx2_ASAP7_75t_L g3856 ( 
.A(n_3319),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_SL g3857 ( 
.A1(n_3107),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3857)
);

INVx8_ASAP7_75t_L g3858 ( 
.A(n_2781),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_SL g3859 ( 
.A(n_2939),
.B(n_903),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_2876),
.B(n_904),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3028),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3041),
.Y(n_3862)
);

OAI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3119),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_2807),
.B(n_88),
.Y(n_3864)
);

INVx1_ASAP7_75t_SL g3865 ( 
.A(n_3347),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_SL g3866 ( 
.A(n_2876),
.B(n_905),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3054),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_SL g3868 ( 
.A(n_2890),
.B(n_905),
.Y(n_3868)
);

INVx2_ASAP7_75t_SL g3869 ( 
.A(n_3261),
.Y(n_3869)
);

OAI21xp33_ASAP7_75t_L g3870 ( 
.A1(n_2987),
.A2(n_89),
.B(n_90),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3012),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_SL g3872 ( 
.A(n_2890),
.B(n_906),
.Y(n_3872)
);

INVx2_ASAP7_75t_SL g3873 ( 
.A(n_3261),
.Y(n_3873)
);

INVx8_ASAP7_75t_L g3874 ( 
.A(n_2781),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_2812),
.B(n_90),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_2813),
.B(n_91),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3016),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_2897),
.B(n_907),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3057),
.Y(n_3879)
);

INVx2_ASAP7_75t_SL g3880 ( 
.A(n_3345),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_2815),
.B(n_91),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_2897),
.B(n_907),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_2821),
.B(n_91),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_2827),
.B(n_92),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_2902),
.B(n_2833),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_2863),
.B(n_92),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_2902),
.B(n_908),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3163),
.B(n_93),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3064),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3074),
.Y(n_3890)
);

AOI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3037),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3891)
);

NOR2xp33_ASAP7_75t_L g3892 ( 
.A(n_3166),
.B(n_93),
.Y(n_3892)
);

INVxp67_ASAP7_75t_L g3893 ( 
.A(n_3142),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3036),
.Y(n_3894)
);

NAND2xp33_ASAP7_75t_L g3895 ( 
.A(n_3110),
.B(n_94),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3075),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_2764),
.B(n_908),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_SL g3898 ( 
.A(n_2764),
.B(n_909),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3052),
.Y(n_3899)
);

CKINVDCx5p33_ASAP7_75t_R g3900 ( 
.A(n_3233),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_L g3901 ( 
.A(n_3185),
.B(n_3193),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_2768),
.B(n_2782),
.Y(n_3902)
);

NOR2xp33_ASAP7_75t_L g3903 ( 
.A(n_3157),
.B(n_94),
.Y(n_3903)
);

NOR2xp67_ASAP7_75t_SL g3904 ( 
.A(n_3007),
.B(n_95),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_2872),
.B(n_95),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_2874),
.B(n_96),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3045),
.B(n_96),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3078),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_2977),
.A2(n_2981),
.B1(n_2984),
.B2(n_3046),
.Y(n_3909)
);

AOI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3037),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_3910)
);

NOR2xp33_ASAP7_75t_L g3911 ( 
.A(n_3295),
.B(n_97),
.Y(n_3911)
);

NOR2xp33_ASAP7_75t_L g3912 ( 
.A(n_3359),
.B(n_97),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3055),
.B(n_98),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_2991),
.B(n_99),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3365),
.B(n_99),
.Y(n_3915)
);

NOR2xp67_ASAP7_75t_L g3916 ( 
.A(n_2776),
.B(n_100),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_2768),
.B(n_909),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3005),
.B(n_99),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3009),
.B(n_100),
.Y(n_3919)
);

INVxp67_ASAP7_75t_L g3920 ( 
.A(n_2782),
.Y(n_3920)
);

AOI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3037),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_3921)
);

OR2x2_ASAP7_75t_L g3922 ( 
.A(n_3248),
.B(n_101),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3071),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3159),
.B(n_102),
.Y(n_3924)
);

INVx4_ASAP7_75t_L g3925 ( 
.A(n_3248),
.Y(n_3925)
);

NOR2xp67_ASAP7_75t_L g3926 ( 
.A(n_2786),
.B(n_104),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_SL g3927 ( 
.A(n_2912),
.B(n_910),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3066),
.B(n_103),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_2912),
.B(n_911),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_2917),
.B(n_912),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_SL g3931 ( 
.A(n_2917),
.B(n_912),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3066),
.B(n_103),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3378),
.B(n_3084),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3080),
.Y(n_3934)
);

A2O1A1Ixp33_ASAP7_75t_L g3935 ( 
.A1(n_3137),
.A2(n_106),
.B(n_103),
.C(n_104),
.Y(n_3935)
);

CKINVDCx5p33_ASAP7_75t_R g3936 ( 
.A(n_3233),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_L g3937 ( 
.A(n_2831),
.B(n_106),
.Y(n_3937)
);

OR2x2_ASAP7_75t_L g3938 ( 
.A(n_3264),
.B(n_106),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3031),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3032),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_SL g3941 ( 
.A(n_3047),
.B(n_913),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3047),
.B(n_913),
.Y(n_3942)
);

NOR2xp33_ASAP7_75t_L g3943 ( 
.A(n_3134),
.B(n_107),
.Y(n_3943)
);

NOR2xp33_ASAP7_75t_L g3944 ( 
.A(n_3198),
.B(n_107),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3047),
.B(n_914),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_2852),
.B(n_108),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_2998),
.B(n_108),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3167),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3127),
.B(n_109),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3129),
.B(n_109),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3132),
.B(n_109),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_2943),
.B(n_110),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3188),
.B(n_110),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3083),
.B(n_110),
.Y(n_3954)
);

INVx3_ASAP7_75t_L g3955 ( 
.A(n_3384),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3083),
.B(n_111),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_3196),
.B(n_111),
.Y(n_3957)
);

OAI22xp5_ASAP7_75t_L g3958 ( 
.A1(n_3160),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3095),
.B(n_112),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3095),
.B(n_113),
.Y(n_3960)
);

OAI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3119),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_3961)
);

NOR2x1_ASAP7_75t_L g3962 ( 
.A(n_3264),
.B(n_114),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3060),
.B(n_915),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_3186),
.B(n_115),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3097),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3114),
.B(n_116),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_2999),
.B(n_116),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3126),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3000),
.B(n_116),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3680),
.B(n_2981),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3460),
.B(n_3173),
.Y(n_3971)
);

INVx3_ASAP7_75t_L g3972 ( 
.A(n_3792),
.Y(n_3972)
);

AND2x2_ASAP7_75t_SL g3973 ( 
.A(n_3560),
.B(n_3370),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3476),
.Y(n_3974)
);

BUFx12f_ASAP7_75t_L g3975 ( 
.A(n_3900),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_L g3976 ( 
.A1(n_3535),
.A2(n_2984),
.B1(n_3194),
.B2(n_3037),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3460),
.B(n_3169),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3427),
.B(n_3008),
.Y(n_3978)
);

NOR2x2_ASAP7_75t_L g3979 ( 
.A(n_3663),
.B(n_3370),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3477),
.Y(n_3980)
);

INVx2_ASAP7_75t_SL g3981 ( 
.A(n_3446),
.Y(n_3981)
);

AND2x4_ASAP7_75t_L g3982 ( 
.A(n_3577),
.B(n_3138),
.Y(n_3982)
);

CKINVDCx8_ASAP7_75t_R g3983 ( 
.A(n_3459),
.Y(n_3983)
);

OAI22xp33_ASAP7_75t_L g3984 ( 
.A1(n_3663),
.A2(n_3051),
.B1(n_3087),
.B2(n_3002),
.Y(n_3984)
);

INVx2_ASAP7_75t_L g3985 ( 
.A(n_3479),
.Y(n_3985)
);

AOI21x1_ASAP7_75t_L g3986 ( 
.A1(n_3579),
.A2(n_2837),
.B(n_3162),
.Y(n_3986)
);

BUFx2_ASAP7_75t_L g3987 ( 
.A(n_3657),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3429),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_3577),
.B(n_3174),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3577),
.B(n_2786),
.Y(n_3990)
);

INVx2_ASAP7_75t_L g3991 ( 
.A(n_3483),
.Y(n_3991)
);

INVx2_ASAP7_75t_SL g3992 ( 
.A(n_3446),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3457),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3552),
.B(n_3060),
.Y(n_3994)
);

AND2x4_ASAP7_75t_L g3995 ( 
.A(n_3509),
.B(n_2787),
.Y(n_3995)
);

NOR3xp33_ASAP7_75t_L g3996 ( 
.A(n_3467),
.B(n_3131),
.C(n_3175),
.Y(n_3996)
);

INVx4_ASAP7_75t_L g3997 ( 
.A(n_3446),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3458),
.B(n_3317),
.Y(n_3998)
);

NOR2x2_ASAP7_75t_L g3999 ( 
.A(n_3663),
.B(n_3267),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3481),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_L g4001 ( 
.A(n_3901),
.B(n_3194),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3497),
.B(n_3482),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3494),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3512),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3531),
.B(n_3509),
.Y(n_4005)
);

INVx5_ASAP7_75t_L g4006 ( 
.A(n_3657),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3515),
.Y(n_4007)
);

CKINVDCx5p33_ASAP7_75t_R g4008 ( 
.A(n_3415),
.Y(n_4008)
);

INVxp67_ASAP7_75t_L g4009 ( 
.A(n_3480),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3524),
.B(n_3321),
.Y(n_4010)
);

OR2x6_ASAP7_75t_L g4011 ( 
.A(n_3605),
.B(n_3266),
.Y(n_4011)
);

AND2x2_ASAP7_75t_SL g4012 ( 
.A(n_3608),
.B(n_3002),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3485),
.Y(n_4013)
);

INVx3_ASAP7_75t_L g4014 ( 
.A(n_3792),
.Y(n_4014)
);

BUFx3_ASAP7_75t_L g4015 ( 
.A(n_3633),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3519),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3531),
.B(n_3060),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3509),
.B(n_2873),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3520),
.Y(n_4019)
);

CKINVDCx5p33_ASAP7_75t_R g4020 ( 
.A(n_3764),
.Y(n_4020)
);

AND2x4_ASAP7_75t_L g4021 ( 
.A(n_3565),
.B(n_2787),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3525),
.B(n_3362),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3411),
.Y(n_4023)
);

INVx3_ASAP7_75t_L g4024 ( 
.A(n_3925),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3416),
.Y(n_4025)
);

BUFx6f_ASAP7_75t_L g4026 ( 
.A(n_3657),
.Y(n_4026)
);

INVxp67_ASAP7_75t_L g4027 ( 
.A(n_3528),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_SL g4028 ( 
.A(n_3565),
.B(n_2954),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3424),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_SL g4030 ( 
.A(n_3565),
.B(n_3551),
.Y(n_4030)
);

A2O1A1Ixp33_ASAP7_75t_L g4031 ( 
.A1(n_3847),
.A2(n_2968),
.B(n_3099),
.C(n_3065),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3529),
.B(n_3147),
.Y(n_4032)
);

AND2x4_ASAP7_75t_L g4033 ( 
.A(n_3491),
.B(n_3495),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3530),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3665),
.B(n_2883),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3433),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3715),
.B(n_3178),
.Y(n_4037)
);

CKINVDCx5p33_ASAP7_75t_R g4038 ( 
.A(n_3936),
.Y(n_4038)
);

CKINVDCx20_ASAP7_75t_R g4039 ( 
.A(n_3568),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3836),
.B(n_3158),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3417),
.B(n_3181),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3498),
.B(n_3213),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_L g4043 ( 
.A1(n_3628),
.A2(n_3194),
.B1(n_3096),
.B2(n_3161),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3452),
.B(n_2954),
.Y(n_4044)
);

AOI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_3405),
.A2(n_3096),
.B1(n_2781),
.B2(n_3029),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3540),
.Y(n_4046)
);

NOR2x1p5_ASAP7_75t_L g4047 ( 
.A(n_3925),
.B(n_2894),
.Y(n_4047)
);

AND2x4_ASAP7_75t_L g4048 ( 
.A(n_3499),
.B(n_3213),
.Y(n_4048)
);

OAI21xp33_ASAP7_75t_SL g4049 ( 
.A1(n_3619),
.A2(n_2862),
.B(n_2853),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_3591),
.Y(n_4050)
);

AND2x4_ASAP7_75t_L g4051 ( 
.A(n_3500),
.B(n_3507),
.Y(n_4051)
);

AND2x4_ASAP7_75t_SL g4052 ( 
.A(n_3753),
.B(n_3345),
.Y(n_4052)
);

INVx4_ASAP7_75t_L g4053 ( 
.A(n_3605),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3555),
.Y(n_4054)
);

INVx1_ASAP7_75t_SL g4055 ( 
.A(n_3865),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3566),
.Y(n_4056)
);

BUFx6f_ASAP7_75t_L g4057 ( 
.A(n_3799),
.Y(n_4057)
);

INVx3_ASAP7_75t_L g4058 ( 
.A(n_3534),
.Y(n_4058)
);

NOR2xp67_ASAP7_75t_L g4059 ( 
.A(n_3410),
.B(n_3266),
.Y(n_4059)
);

CKINVDCx5p33_ASAP7_75t_R g4060 ( 
.A(n_3591),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3569),
.Y(n_4061)
);

NAND2x1p5_ASAP7_75t_L g4062 ( 
.A(n_3608),
.B(n_3268),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3571),
.B(n_3182),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3436),
.Y(n_4064)
);

O2A1O1Ixp5_ASAP7_75t_L g4065 ( 
.A1(n_3489),
.A2(n_3192),
.B(n_2891),
.C(n_2871),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3572),
.B(n_3140),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3574),
.Y(n_4067)
);

BUFx6f_ASAP7_75t_L g4068 ( 
.A(n_3799),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3592),
.Y(n_4069)
);

INVx1_ASAP7_75t_SL g4070 ( 
.A(n_3856),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3593),
.Y(n_4071)
);

BUFx6f_ASAP7_75t_L g4072 ( 
.A(n_3799),
.Y(n_4072)
);

INVx3_ASAP7_75t_L g4073 ( 
.A(n_3605),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_SL g4074 ( 
.A(n_3581),
.B(n_2820),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3594),
.B(n_2851),
.Y(n_4075)
);

BUFx6f_ASAP7_75t_L g4076 ( 
.A(n_3813),
.Y(n_4076)
);

INVx3_ASAP7_75t_L g4077 ( 
.A(n_3675),
.Y(n_4077)
);

AOI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_3396),
.A2(n_3336),
.B1(n_3171),
.B2(n_3165),
.Y(n_4078)
);

OAI21x1_ASAP7_75t_L g4079 ( 
.A1(n_3650),
.A2(n_3145),
.B(n_3130),
.Y(n_4079)
);

CKINVDCx5p33_ASAP7_75t_R g4080 ( 
.A(n_3766),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3581),
.B(n_2832),
.Y(n_4081)
);

CKINVDCx6p67_ASAP7_75t_R g4082 ( 
.A(n_3723),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3439),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3598),
.Y(n_4084)
);

BUFx2_ASAP7_75t_L g4085 ( 
.A(n_3753),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3600),
.B(n_3693),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_3928),
.B(n_3200),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3934),
.Y(n_4088)
);

AND2x6_ASAP7_75t_L g4089 ( 
.A(n_3955),
.B(n_2832),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3602),
.Y(n_4090)
);

BUFx6f_ASAP7_75t_L g4091 ( 
.A(n_3813),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_3461),
.A2(n_2850),
.B(n_2832),
.Y(n_4092)
);

NOR2xp33_ASAP7_75t_L g4093 ( 
.A(n_3846),
.B(n_3721),
.Y(n_4093)
);

INVx4_ASAP7_75t_L g4094 ( 
.A(n_3753),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3603),
.B(n_2858),
.Y(n_4095)
);

INVx5_ASAP7_75t_L g4096 ( 
.A(n_3404),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3932),
.B(n_2978),
.Y(n_4097)
);

NOR2xp33_ASAP7_75t_R g4098 ( 
.A(n_3454),
.B(n_3069),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_3513),
.B(n_3275),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3610),
.B(n_2889),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_SL g4101 ( 
.A(n_3600),
.B(n_2850),
.Y(n_4101)
);

CKINVDCx16_ASAP7_75t_R g4102 ( 
.A(n_3845),
.Y(n_4102)
);

AND2x4_ASAP7_75t_L g4103 ( 
.A(n_3517),
.B(n_3275),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3440),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3614),
.B(n_3034),
.Y(n_4105)
);

AOI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_3533),
.A2(n_3092),
.B1(n_2905),
.B2(n_3079),
.Y(n_4106)
);

AND2x4_ASAP7_75t_SL g4107 ( 
.A(n_3788),
.B(n_3268),
.Y(n_4107)
);

INVx5_ASAP7_75t_L g4108 ( 
.A(n_3404),
.Y(n_4108)
);

INVx3_ASAP7_75t_L g4109 ( 
.A(n_3788),
.Y(n_4109)
);

AND2x4_ASAP7_75t_L g4110 ( 
.A(n_3508),
.B(n_3311),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3688),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3399),
.B(n_3070),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_SL g4113 ( 
.A(n_3693),
.B(n_2850),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3576),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3409),
.B(n_3183),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3606),
.Y(n_4116)
);

CKINVDCx5p33_ASAP7_75t_R g4117 ( 
.A(n_3541),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3536),
.B(n_2974),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3612),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3447),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_3578),
.B(n_3085),
.Y(n_4121)
);

AND2x4_ASAP7_75t_L g4122 ( 
.A(n_3508),
.B(n_3311),
.Y(n_4122)
);

INVx4_ASAP7_75t_L g4123 ( 
.A(n_3788),
.Y(n_4123)
);

AOI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3776),
.A2(n_3096),
.B1(n_3199),
.B2(n_2781),
.Y(n_4124)
);

AOI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_3595),
.A2(n_3096),
.B1(n_3102),
.B2(n_3051),
.Y(n_4125)
);

AND2x4_ASAP7_75t_L g4126 ( 
.A(n_3617),
.B(n_3339),
.Y(n_4126)
);

INVxp67_ASAP7_75t_L g4127 ( 
.A(n_3621),
.Y(n_4127)
);

AOI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_3623),
.A2(n_2927),
.B(n_2870),
.Y(n_4128)
);

CKINVDCx5p33_ASAP7_75t_R g4129 ( 
.A(n_3783),
.Y(n_4129)
);

INVx3_ASAP7_75t_L g4130 ( 
.A(n_3526),
.Y(n_4130)
);

INVx2_ASAP7_75t_L g4131 ( 
.A(n_3434),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3445),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_SL g4133 ( 
.A(n_3619),
.B(n_2870),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3770),
.B(n_3113),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_3719),
.B(n_2744),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3456),
.Y(n_4136)
);

NOR3xp33_ASAP7_75t_SL g4137 ( 
.A(n_3588),
.B(n_3857),
.C(n_3503),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3627),
.Y(n_4138)
);

INVx3_ASAP7_75t_L g4139 ( 
.A(n_3422),
.Y(n_4139)
);

BUFx6f_ASAP7_75t_L g4140 ( 
.A(n_3813),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_SL g4141 ( 
.A(n_3406),
.B(n_2870),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3397),
.B(n_2747),
.Y(n_4142)
);

O2A1O1Ixp33_ASAP7_75t_L g4143 ( 
.A1(n_3403),
.A2(n_3423),
.B(n_3734),
.C(n_3698),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3768),
.Y(n_4144)
);

AND2x4_ASAP7_75t_L g4145 ( 
.A(n_3617),
.B(n_3339),
.Y(n_4145)
);

AND2x6_ASAP7_75t_L g4146 ( 
.A(n_3955),
.B(n_2927),
.Y(n_4146)
);

NOR2xp33_ASAP7_75t_L g4147 ( 
.A(n_3643),
.B(n_3281),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3412),
.B(n_2760),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3632),
.Y(n_4149)
);

BUFx3_ASAP7_75t_L g4150 ( 
.A(n_3464),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3414),
.B(n_3215),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_3778),
.Y(n_4152)
);

AND2x4_ASAP7_75t_L g4153 ( 
.A(n_3654),
.B(n_3360),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_SL g4154 ( 
.A(n_3406),
.B(n_2927),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_3909),
.B(n_3240),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3636),
.Y(n_4156)
);

OR2x2_ASAP7_75t_L g4157 ( 
.A(n_3705),
.B(n_3332),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_3545),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3660),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3789),
.B(n_3382),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3729),
.B(n_3393),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_SL g4162 ( 
.A(n_3406),
.B(n_2931),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_SL g4163 ( 
.A(n_3406),
.B(n_2931),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_SL g4164 ( 
.A(n_3406),
.B(n_2931),
.Y(n_4164)
);

AND2x4_ASAP7_75t_L g4165 ( 
.A(n_3654),
.B(n_3360),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_R g4166 ( 
.A(n_3858),
.B(n_3281),
.Y(n_4166)
);

BUFx4f_ASAP7_75t_L g4167 ( 
.A(n_3786),
.Y(n_4167)
);

BUFx3_ASAP7_75t_L g4168 ( 
.A(n_3618),
.Y(n_4168)
);

BUFx6f_ASAP7_75t_L g4169 ( 
.A(n_3640),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_3547),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_L g4171 ( 
.A1(n_3601),
.A2(n_3189),
.B1(n_3099),
.B2(n_3065),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3669),
.Y(n_4172)
);

INVx5_ASAP7_75t_L g4173 ( 
.A(n_3404),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3798),
.Y(n_4174)
);

BUFx3_ASAP7_75t_L g4175 ( 
.A(n_3696),
.Y(n_4175)
);

INVx3_ASAP7_75t_L g4176 ( 
.A(n_3730),
.Y(n_4176)
);

AND2x4_ASAP7_75t_L g4177 ( 
.A(n_3658),
.B(n_3390),
.Y(n_4177)
);

NAND2x1p5_ASAP7_75t_L g4178 ( 
.A(n_3546),
.B(n_3302),
.Y(n_4178)
);

OAI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_3891),
.A2(n_3176),
.B1(n_3192),
.B2(n_3103),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3762),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3765),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3767),
.B(n_3128),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_3557),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3620),
.B(n_3010),
.Y(n_4184)
);

AOI22xp33_ASAP7_75t_L g4185 ( 
.A1(n_3625),
.A2(n_3189),
.B1(n_3100),
.B2(n_2992),
.Y(n_4185)
);

AOI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_3853),
.A2(n_3141),
.B1(n_3087),
.B2(n_2773),
.Y(n_4186)
);

NOR2xp33_ASAP7_75t_L g4187 ( 
.A(n_3774),
.B(n_3302),
.Y(n_4187)
);

AOI22xp5_ASAP7_75t_L g4188 ( 
.A1(n_3843),
.A2(n_3141),
.B1(n_2800),
.B2(n_2817),
.Y(n_4188)
);

OR2x6_ASAP7_75t_L g4189 ( 
.A(n_3858),
.B(n_3349),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3559),
.Y(n_4190)
);

OR2x2_ASAP7_75t_L g4191 ( 
.A(n_3745),
.B(n_3349),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_3542),
.B(n_3358),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_SL g4193 ( 
.A(n_3891),
.B(n_2950),
.Y(n_4193)
);

AND2x4_ASAP7_75t_L g4194 ( 
.A(n_3658),
.B(n_3390),
.Y(n_4194)
);

AOI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_3819),
.A2(n_3369),
.B1(n_3381),
.B2(n_3358),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_3419),
.B(n_3369),
.Y(n_4196)
);

BUFx8_ASAP7_75t_L g4197 ( 
.A(n_3735),
.Y(n_4197)
);

INVx5_ASAP7_75t_L g4198 ( 
.A(n_3404),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_SL g4199 ( 
.A(n_3910),
.B(n_2950),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_3682),
.B(n_3044),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3820),
.B(n_3381),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_3844),
.B(n_3105),
.Y(n_4202)
);

OR2x6_ASAP7_75t_L g4203 ( 
.A(n_3858),
.B(n_2967),
.Y(n_4203)
);

O2A1O1Ixp33_ASAP7_75t_L g4204 ( 
.A1(n_3470),
.A2(n_3104),
.B(n_3108),
.C(n_3098),
.Y(n_4204)
);

INVx2_ASAP7_75t_SL g4205 ( 
.A(n_3752),
.Y(n_4205)
);

NOR2xp33_ASAP7_75t_L g4206 ( 
.A(n_3797),
.B(n_3740),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3822),
.B(n_3100),
.Y(n_4207)
);

BUFx4f_ASAP7_75t_L g4208 ( 
.A(n_3438),
.Y(n_4208)
);

NAND2x1p5_ASAP7_75t_L g4209 ( 
.A(n_3546),
.B(n_3105),
.Y(n_4209)
);

AND2x4_ASAP7_75t_SL g4210 ( 
.A(n_3438),
.B(n_3103),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_SL g4211 ( 
.A(n_3910),
.B(n_2950),
.Y(n_4211)
);

AOI22xp5_ASAP7_75t_L g4212 ( 
.A1(n_3888),
.A2(n_3109),
.B1(n_3001),
.B2(n_2996),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_3921),
.B(n_2957),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_SL g4214 ( 
.A(n_3921),
.B(n_2957),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_3561),
.Y(n_4215)
);

HB1xp67_ASAP7_75t_L g4216 ( 
.A(n_3893),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3773),
.Y(n_4217)
);

AND2x4_ASAP7_75t_L g4218 ( 
.A(n_3834),
.B(n_2819),
.Y(n_4218)
);

AND2x6_ASAP7_75t_L g4219 ( 
.A(n_3589),
.B(n_2957),
.Y(n_4219)
);

INVx3_ASAP7_75t_L g4220 ( 
.A(n_3755),
.Y(n_4220)
);

INVx5_ASAP7_75t_L g4221 ( 
.A(n_3874),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3648),
.B(n_3105),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3787),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_3810),
.B(n_3115),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_3501),
.B(n_3153),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_3687),
.B(n_117),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_3834),
.B(n_2819),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3794),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_3510),
.B(n_3626),
.Y(n_4229)
);

NOR3xp33_ASAP7_75t_SL g4230 ( 
.A(n_3863),
.B(n_3961),
.C(n_3402),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_SL g4231 ( 
.A(n_3465),
.B(n_2960),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_3795),
.Y(n_4232)
);

AOI21xp33_ASAP7_75t_L g4233 ( 
.A1(n_3504),
.A2(n_3201),
.B(n_2866),
.Y(n_4233)
);

BUFx3_ASAP7_75t_L g4234 ( 
.A(n_3708),
.Y(n_4234)
);

A2O1A1Ixp33_ASAP7_75t_L g4235 ( 
.A1(n_3649),
.A2(n_3106),
.B(n_3180),
.C(n_3156),
.Y(n_4235)
);

NOR2xp33_ASAP7_75t_L g4236 ( 
.A(n_3492),
.B(n_3153),
.Y(n_4236)
);

CKINVDCx5p33_ASAP7_75t_R g4237 ( 
.A(n_3438),
.Y(n_4237)
);

INVx2_ASAP7_75t_SL g4238 ( 
.A(n_3848),
.Y(n_4238)
);

INVx5_ASAP7_75t_L g4239 ( 
.A(n_3874),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_3408),
.B(n_3156),
.Y(n_4240)
);

INVx2_ASAP7_75t_SL g4241 ( 
.A(n_3869),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_3850),
.Y(n_4242)
);

CKINVDCx20_ASAP7_75t_R g4243 ( 
.A(n_3885),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_3567),
.Y(n_4244)
);

INVx2_ASAP7_75t_SL g4245 ( 
.A(n_3873),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3596),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3413),
.B(n_3180),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_SL g4248 ( 
.A(n_3465),
.B(n_2960),
.Y(n_4248)
);

OR2x6_ASAP7_75t_L g4249 ( 
.A(n_3874),
.B(n_2967),
.Y(n_4249)
);

INVx5_ASAP7_75t_L g4250 ( 
.A(n_3640),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_3616),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_3624),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_3563),
.B(n_3516),
.Y(n_4253)
);

CKINVDCx5p33_ASAP7_75t_R g4254 ( 
.A(n_3880),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_3916),
.B(n_2960),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_3862),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_3634),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_SL g4258 ( 
.A(n_3916),
.B(n_3926),
.Y(n_4258)
);

AOI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_3892),
.A2(n_3189),
.B1(n_3106),
.B2(n_2924),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_3420),
.B(n_3120),
.Y(n_4260)
);

AND2x4_ASAP7_75t_L g4261 ( 
.A(n_3926),
.B(n_2829),
.Y(n_4261)
);

BUFx2_ASAP7_75t_L g4262 ( 
.A(n_3728),
.Y(n_4262)
);

OAI21xp33_ASAP7_75t_SL g4263 ( 
.A1(n_3732),
.A2(n_3738),
.B(n_3718),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3867),
.Y(n_4264)
);

INVx3_ASAP7_75t_L g4265 ( 
.A(n_3589),
.Y(n_4265)
);

INVx3_ASAP7_75t_L g4266 ( 
.A(n_3487),
.Y(n_4266)
);

AOI22xp5_ASAP7_75t_SL g4267 ( 
.A1(n_3785),
.A2(n_3093),
.B1(n_3259),
.B2(n_3116),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3428),
.B(n_3120),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3879),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3430),
.B(n_3123),
.Y(n_4270)
);

OAI21xp33_ASAP7_75t_L g4271 ( 
.A1(n_3903),
.A2(n_3172),
.B(n_3170),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_SL g4272 ( 
.A(n_3487),
.B(n_2973),
.Y(n_4272)
);

BUFx6f_ASAP7_75t_L g4273 ( 
.A(n_3640),
.Y(n_4273)
);

INVx2_ASAP7_75t_SL g4274 ( 
.A(n_3922),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3441),
.B(n_3123),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_3679),
.A2(n_3013),
.B(n_2973),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_3694),
.B(n_117),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_3635),
.Y(n_4278)
);

INVx3_ASAP7_75t_L g4279 ( 
.A(n_3938),
.Y(n_4279)
);

OAI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_3484),
.A2(n_3189),
.B(n_2924),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_3889),
.Y(n_4281)
);

BUFx12f_ASAP7_75t_L g4282 ( 
.A(n_3841),
.Y(n_4282)
);

BUFx3_ASAP7_75t_L g4283 ( 
.A(n_3455),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_3443),
.B(n_3149),
.Y(n_4284)
);

BUFx5_ASAP7_75t_L g4285 ( 
.A(n_3692),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_3444),
.B(n_3149),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_SL g4287 ( 
.A(n_3732),
.B(n_2973),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_L g4288 ( 
.A(n_3659),
.B(n_3149),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_L g4289 ( 
.A(n_3724),
.B(n_3093),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_3642),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_3448),
.B(n_3116),
.Y(n_4291)
);

NOR2xp33_ASAP7_75t_L g4292 ( 
.A(n_3674),
.B(n_3259),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_3488),
.B(n_2829),
.Y(n_4293)
);

BUFx2_ASAP7_75t_L g4294 ( 
.A(n_3455),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_SL g4295 ( 
.A(n_3738),
.B(n_3013),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3449),
.B(n_3379),
.Y(n_4296)
);

BUFx2_ASAP7_75t_L g4297 ( 
.A(n_3474),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_3666),
.Y(n_4298)
);

BUFx6f_ASAP7_75t_SL g4299 ( 
.A(n_3890),
.Y(n_4299)
);

CKINVDCx16_ASAP7_75t_R g4300 ( 
.A(n_3771),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3450),
.B(n_3379),
.Y(n_4301)
);

NOR2xp33_ASAP7_75t_L g4302 ( 
.A(n_3425),
.B(n_2845),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_3896),
.Y(n_4303)
);

BUFx6f_ASAP7_75t_L g4304 ( 
.A(n_3646),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_3641),
.B(n_2845),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3908),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_3802),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3672),
.Y(n_4308)
);

INVxp67_ASAP7_75t_L g4309 ( 
.A(n_3582),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_3673),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_3823),
.B(n_2854),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_3676),
.Y(n_4312)
);

NAND2xp33_ASAP7_75t_L g4313 ( 
.A(n_3644),
.B(n_3331),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_3806),
.B(n_2854),
.Y(n_4314)
);

A2O1A1Ixp33_ASAP7_75t_L g4315 ( 
.A1(n_3805),
.A2(n_2899),
.B(n_2929),
.C(n_2909),
.Y(n_4315)
);

INVx4_ASAP7_75t_L g4316 ( 
.A(n_3474),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_3704),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_3814),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3818),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_3706),
.Y(n_4320)
);

BUFx3_ASAP7_75t_L g4321 ( 
.A(n_3701),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_SL g4322 ( 
.A(n_3718),
.B(n_3013),
.Y(n_4322)
);

AOI22xp33_ASAP7_75t_L g4323 ( 
.A1(n_3506),
.A2(n_3689),
.B1(n_3943),
.B2(n_3828),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_3826),
.B(n_3833),
.Y(n_4324)
);

OR2x6_ASAP7_75t_L g4325 ( 
.A(n_3962),
.B(n_2899),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_3714),
.Y(n_4326)
);

BUFx3_ASAP7_75t_L g4327 ( 
.A(n_3712),
.Y(n_4327)
);

A2O1A1Ixp33_ASAP7_75t_L g4328 ( 
.A1(n_3895),
.A2(n_2909),
.B(n_2929),
.C(n_2935),
.Y(n_4328)
);

BUFx3_ASAP7_75t_L g4329 ( 
.A(n_3722),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_3518),
.B(n_117),
.Y(n_4330)
);

BUFx3_ASAP7_75t_L g4331 ( 
.A(n_3733),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3939),
.B(n_2935),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_3940),
.B(n_2965),
.Y(n_4333)
);

AND2x6_ASAP7_75t_SL g4334 ( 
.A(n_3803),
.B(n_118),
.Y(n_4334)
);

AOI22xp33_ASAP7_75t_SL g4335 ( 
.A1(n_3421),
.A2(n_3290),
.B1(n_3331),
.B2(n_3273),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_3748),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3750),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3754),
.Y(n_4338)
);

OR2x2_ASAP7_75t_SL g4339 ( 
.A(n_3691),
.B(n_119),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_3761),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_3717),
.Y(n_4341)
);

HB1xp67_ASAP7_75t_L g4342 ( 
.A(n_3725),
.Y(n_4342)
);

INVx2_ASAP7_75t_SL g4343 ( 
.A(n_3839),
.Y(n_4343)
);

O2A1O1Ixp5_ASAP7_75t_L g4344 ( 
.A1(n_3418),
.A2(n_3205),
.B(n_2738),
.C(n_2993),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_3744),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_3746),
.Y(n_4346)
);

AOI22xp5_ASAP7_75t_L g4347 ( 
.A1(n_3743),
.A2(n_2924),
.B1(n_3290),
.B2(n_3273),
.Y(n_4347)
);

AOI21xp5_ASAP7_75t_L g4348 ( 
.A1(n_3442),
.A2(n_3067),
.B(n_3062),
.Y(n_4348)
);

BUFx6f_ASAP7_75t_L g4349 ( 
.A(n_3646),
.Y(n_4349)
);

BUFx3_ASAP7_75t_L g4350 ( 
.A(n_3747),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_3505),
.B(n_2993),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_SL g4352 ( 
.A(n_3664),
.B(n_3062),
.Y(n_4352)
);

AOI22xp5_ASAP7_75t_L g4353 ( 
.A1(n_3751),
.A2(n_2924),
.B1(n_3290),
.B2(n_3273),
.Y(n_4353)
);

INVx2_ASAP7_75t_SL g4354 ( 
.A(n_3466),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_3948),
.Y(n_4355)
);

INVx4_ASAP7_75t_L g4356 ( 
.A(n_3646),
.Y(n_4356)
);

OAI22xp5_ASAP7_75t_SL g4357 ( 
.A1(n_3587),
.A2(n_3015),
.B1(n_3024),
.B2(n_2965),
.Y(n_4357)
);

NOR2xp33_ASAP7_75t_L g4358 ( 
.A(n_3435),
.B(n_3015),
.Y(n_4358)
);

AOI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_3911),
.A2(n_2963),
.B1(n_3024),
.B2(n_3273),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3573),
.Y(n_4360)
);

NAND2xp33_ASAP7_75t_L g4361 ( 
.A(n_3681),
.B(n_3290),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3575),
.Y(n_4362)
);

OAI22xp5_ASAP7_75t_L g4363 ( 
.A1(n_3664),
.A2(n_3062),
.B1(n_3068),
.B2(n_3067),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_3580),
.Y(n_4364)
);

NOR2xp33_ASAP7_75t_R g4365 ( 
.A(n_3681),
.B(n_3331),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_3583),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_3586),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_3736),
.B(n_118),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_SL g4369 ( 
.A(n_3681),
.B(n_3067),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_SL g4370 ( 
.A(n_3830),
.B(n_3068),
.Y(n_4370)
);

NAND2x1_ASAP7_75t_L g4371 ( 
.A(n_3965),
.B(n_3331),
.Y(n_4371)
);

NAND2x1p5_ASAP7_75t_L g4372 ( 
.A(n_3831),
.B(n_2963),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_3830),
.B(n_3068),
.Y(n_4373)
);

INVx1_ASAP7_75t_SL g4374 ( 
.A(n_3407),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_3590),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_3781),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_SL g4377 ( 
.A(n_3453),
.B(n_3077),
.Y(n_4377)
);

BUFx4f_ASAP7_75t_L g4378 ( 
.A(n_3852),
.Y(n_4378)
);

AND2x2_ASAP7_75t_SL g4379 ( 
.A(n_3821),
.B(n_2963),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3597),
.Y(n_4380)
);

AOI22xp33_ASAP7_75t_L g4381 ( 
.A1(n_3912),
.A2(n_2963),
.B1(n_3094),
.B2(n_3077),
.Y(n_4381)
);

BUFx3_ASAP7_75t_L g4382 ( 
.A(n_3790),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_3739),
.B(n_119),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_SL g4384 ( 
.A(n_3821),
.B(n_3077),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_3742),
.B(n_120),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_3791),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_3807),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_3756),
.B(n_121),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_3599),
.Y(n_4389)
);

INVx2_ASAP7_75t_SL g4390 ( 
.A(n_3902),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_3815),
.Y(n_4391)
);

NOR2x1_ASAP7_75t_L g4392 ( 
.A(n_3851),
.B(n_3094),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_3661),
.B(n_121),
.Y(n_4393)
);

AND2x4_ASAP7_75t_L g4394 ( 
.A(n_3720),
.B(n_3094),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_SL g4395 ( 
.A(n_3638),
.B(n_3101),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_3523),
.B(n_122),
.Y(n_4396)
);

INVx3_ASAP7_75t_L g4397 ( 
.A(n_3817),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_3684),
.B(n_122),
.Y(n_4398)
);

OAI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_3914),
.A2(n_3122),
.B(n_3101),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_3604),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_3611),
.Y(n_4401)
);

INVxp67_ASAP7_75t_SL g4402 ( 
.A(n_3968),
.Y(n_4402)
);

INVx3_ASAP7_75t_L g4403 ( 
.A(n_3838),
.Y(n_4403)
);

AND2x2_ASAP7_75t_SL g4404 ( 
.A(n_3638),
.B(n_3101),
.Y(n_4404)
);

INVx4_ASAP7_75t_L g4405 ( 
.A(n_3842),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_3613),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_3686),
.B(n_122),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_L g4408 ( 
.A1(n_3915),
.A2(n_3124),
.B1(n_3133),
.B2(n_3122),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_L g4409 ( 
.A(n_3437),
.B(n_123),
.Y(n_4409)
);

CKINVDCx5p33_ASAP7_75t_R g4410 ( 
.A(n_3398),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_3849),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_SL g4412 ( 
.A(n_3471),
.B(n_3122),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_SL g4413 ( 
.A(n_3870),
.B(n_3124),
.Y(n_4413)
);

HB1xp67_ASAP7_75t_L g4414 ( 
.A(n_3861),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_3871),
.Y(n_4415)
);

AND2x4_ASAP7_75t_L g4416 ( 
.A(n_3877),
.B(n_3124),
.Y(n_4416)
);

NOR2xp67_ASAP7_75t_L g4417 ( 
.A(n_3400),
.B(n_123),
.Y(n_4417)
);

INVxp67_ASAP7_75t_L g4418 ( 
.A(n_3726),
.Y(n_4418)
);

INVx3_ASAP7_75t_L g4419 ( 
.A(n_3894),
.Y(n_4419)
);

AOI21xp5_ASAP7_75t_L g4420 ( 
.A1(n_3486),
.A2(n_3136),
.B(n_3133),
.Y(n_4420)
);

OAI21xp5_ASAP7_75t_L g4421 ( 
.A1(n_3918),
.A2(n_3136),
.B(n_3133),
.Y(n_4421)
);

AND2x4_ASAP7_75t_L g4422 ( 
.A(n_3899),
.B(n_3136),
.Y(n_4422)
);

INVx3_ASAP7_75t_L g4423 ( 
.A(n_3923),
.Y(n_4423)
);

BUFx4f_ASAP7_75t_L g4424 ( 
.A(n_3904),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_3763),
.Y(n_4425)
);

INVx1_ASAP7_75t_SL g4426 ( 
.A(n_3954),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_SL g4427 ( 
.A(n_3683),
.B(n_124),
.Y(n_4427)
);

NOR2x1_ASAP7_75t_L g4428 ( 
.A(n_3859),
.B(n_124),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_3690),
.B(n_124),
.Y(n_4429)
);

INVx1_ASAP7_75t_L g4430 ( 
.A(n_3769),
.Y(n_4430)
);

HB1xp67_ASAP7_75t_L g4431 ( 
.A(n_3920),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_3539),
.Y(n_4432)
);

BUFx12f_ASAP7_75t_L g4433 ( 
.A(n_3749),
.Y(n_4433)
);

OR2x6_ASAP7_75t_L g4434 ( 
.A(n_3784),
.B(n_3801),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_3544),
.Y(n_4435)
);

BUFx12f_ASAP7_75t_L g4436 ( 
.A(n_3757),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_3697),
.B(n_125),
.Y(n_4437)
);

HB1xp67_ASAP7_75t_L g4438 ( 
.A(n_3685),
.Y(n_4438)
);

AND2x6_ASAP7_75t_L g4439 ( 
.A(n_3825),
.B(n_125),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_3933),
.B(n_126),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_SL g4441 ( 
.A(n_3759),
.B(n_126),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_3804),
.B(n_127),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_3775),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_3947),
.Y(n_4444)
);

BUFx4f_ASAP7_75t_L g4445 ( 
.A(n_3860),
.Y(n_4445)
);

INVx5_ASAP7_75t_L g4446 ( 
.A(n_3829),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_SL g4447 ( 
.A(n_3832),
.B(n_127),
.Y(n_4447)
);

AOI22xp5_ASAP7_75t_L g4448 ( 
.A1(n_3702),
.A2(n_3952),
.B1(n_3653),
.B2(n_3431),
.Y(n_4448)
);

NOR2xp33_ASAP7_75t_R g4449 ( 
.A(n_3703),
.B(n_3711),
.Y(n_4449)
);

INVx3_ASAP7_75t_L g4450 ( 
.A(n_3956),
.Y(n_4450)
);

HB1xp67_ASAP7_75t_L g4451 ( 
.A(n_3959),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_3550),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_3967),
.Y(n_4453)
);

AND2x6_ASAP7_75t_SL g4454 ( 
.A(n_3451),
.B(n_127),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_SL g4455 ( 
.A(n_3927),
.B(n_128),
.Y(n_4455)
);

AOI22xp33_ASAP7_75t_L g4456 ( 
.A1(n_3760),
.A2(n_3924),
.B1(n_3957),
.B2(n_3944),
.Y(n_4456)
);

AND2x4_ASAP7_75t_L g4457 ( 
.A(n_3897),
.B(n_128),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3668),
.B(n_128),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_3401),
.B(n_129),
.Y(n_4459)
);

INVx2_ASAP7_75t_SL g4460 ( 
.A(n_3960),
.Y(n_4460)
);

AOI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_3713),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_4461)
);

AND2x4_ASAP7_75t_L g4462 ( 
.A(n_3898),
.B(n_130),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_3670),
.B(n_131),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_3671),
.B(n_133),
.Y(n_4464)
);

INVxp67_ASAP7_75t_SL g4465 ( 
.A(n_3758),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_L g4466 ( 
.A(n_3716),
.B(n_3655),
.Y(n_4466)
);

INVx2_ASAP7_75t_SL g4467 ( 
.A(n_3866),
.Y(n_4467)
);

HB1xp67_ASAP7_75t_L g4468 ( 
.A(n_3469),
.Y(n_4468)
);

INVx3_ASAP7_75t_L g4469 ( 
.A(n_3472),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_SL g4470 ( 
.A(n_3929),
.B(n_133),
.Y(n_4470)
);

BUFx3_ASAP7_75t_L g4471 ( 
.A(n_3473),
.Y(n_4471)
);

AND2x4_ASAP7_75t_SL g4472 ( 
.A(n_3854),
.B(n_133),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_3969),
.Y(n_4473)
);

OAI21xp5_ASAP7_75t_L g4474 ( 
.A1(n_3919),
.A2(n_134),
.B(n_135),
.Y(n_4474)
);

NOR3xp33_ASAP7_75t_SL g4475 ( 
.A(n_3868),
.B(n_134),
.C(n_136),
.Y(n_4475)
);

BUFx12f_ASAP7_75t_L g4476 ( 
.A(n_3872),
.Y(n_4476)
);

A2O1A1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_3629),
.A2(n_137),
.B(n_134),
.C(n_136),
.Y(n_4477)
);

OAI22xp5_ASAP7_75t_L g4478 ( 
.A1(n_3796),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_3462),
.Y(n_4479)
);

BUFx6f_ASAP7_75t_L g4480 ( 
.A(n_3537),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_3553),
.Y(n_4481)
);

CKINVDCx20_ASAP7_75t_R g4482 ( 
.A(n_3468),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_3556),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_3827),
.B(n_137),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_SL g4485 ( 
.A(n_3930),
.B(n_138),
.Y(n_4485)
);

NOR2xp33_ASAP7_75t_L g4486 ( 
.A(n_3812),
.B(n_3907),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_SL g4487 ( 
.A(n_3931),
.B(n_138),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_3558),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_3835),
.B(n_139),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_SL g4490 ( 
.A(n_3811),
.B(n_139),
.Y(n_4490)
);

OR2x2_ASAP7_75t_L g4491 ( 
.A(n_3662),
.B(n_139),
.Y(n_4491)
);

AOI22xp33_ASAP7_75t_L g4492 ( 
.A1(n_3966),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_3645),
.B(n_141),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_3837),
.B(n_141),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_3562),
.Y(n_4495)
);

NOR2xp33_ASAP7_75t_L g4496 ( 
.A(n_3913),
.B(n_142),
.Y(n_4496)
);

INVxp67_ASAP7_75t_L g4497 ( 
.A(n_3651),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_3656),
.B(n_142),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_3564),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_SL g4500 ( 
.A(n_3816),
.B(n_143),
.Y(n_4500)
);

NAND2x1p5_ASAP7_75t_L g4501 ( 
.A(n_3878),
.B(n_143),
.Y(n_4501)
);

INVxp67_ASAP7_75t_L g4502 ( 
.A(n_3652),
.Y(n_4502)
);

BUFx4f_ASAP7_75t_L g4503 ( 
.A(n_3882),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_SL g4504 ( 
.A(n_3700),
.B(n_145),
.Y(n_4504)
);

AO22x1_ASAP7_75t_L g4505 ( 
.A1(n_3958),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_4505)
);

INVx3_ASAP7_75t_L g4506 ( 
.A(n_3570),
.Y(n_4506)
);

CKINVDCx5p33_ASAP7_75t_R g4507 ( 
.A(n_3609),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_3949),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_3585),
.B(n_146),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3950),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_3475),
.Y(n_4511)
);

NOR2x1p5_ASAP7_75t_L g4512 ( 
.A(n_3741),
.B(n_146),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_3840),
.B(n_147),
.Y(n_4513)
);

AO22x1_ASAP7_75t_L g4514 ( 
.A1(n_3737),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4514)
);

INVx2_ASAP7_75t_SL g4515 ( 
.A(n_3887),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_3548),
.A2(n_3864),
.B1(n_3875),
.B2(n_3855),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_3951),
.Y(n_4517)
);

AND2x4_ASAP7_75t_L g4518 ( 
.A(n_3917),
.B(n_148),
.Y(n_4518)
);

BUFx6f_ASAP7_75t_L g4519 ( 
.A(n_3538),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_3478),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_SL g4521 ( 
.A(n_3772),
.B(n_3780),
.Y(n_4521)
);

INVx5_ASAP7_75t_L g4522 ( 
.A(n_3549),
.Y(n_4522)
);

AND2x2_ASAP7_75t_L g4523 ( 
.A(n_3824),
.B(n_149),
.Y(n_4523)
);

OR2x2_ASAP7_75t_L g4524 ( 
.A(n_3953),
.B(n_150),
.Y(n_4524)
);

INVx5_ASAP7_75t_L g4525 ( 
.A(n_3554),
.Y(n_4525)
);

CKINVDCx5p33_ASAP7_75t_R g4526 ( 
.A(n_3964),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_3514),
.A2(n_150),
.B(n_151),
.Y(n_4527)
);

BUFx6f_ASAP7_75t_L g4528 ( 
.A(n_3941),
.Y(n_4528)
);

AOI22xp33_ASAP7_75t_L g4529 ( 
.A1(n_3777),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3521),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_3490),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_3522),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_3432),
.B(n_151),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_3876),
.B(n_3881),
.Y(n_4534)
);

AOI22xp33_ASAP7_75t_L g4535 ( 
.A1(n_3779),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4535)
);

AOI21x1_ASAP7_75t_L g4536 ( 
.A1(n_4030),
.A2(n_3963),
.B(n_3945),
.Y(n_4536)
);

O2A1O1Ixp33_ASAP7_75t_SL g4537 ( 
.A1(n_3984),
.A2(n_3695),
.B(n_3935),
.C(n_3667),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_4114),
.B(n_3426),
.Y(n_4538)
);

A2O1A1Ixp33_ASAP7_75t_L g4539 ( 
.A1(n_4263),
.A2(n_3463),
.B(n_3884),
.C(n_3883),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4116),
.B(n_3496),
.Y(n_4540)
);

BUFx6f_ASAP7_75t_L g4541 ( 
.A(n_4026),
.Y(n_4541)
);

NOR2xp33_ASAP7_75t_L g4542 ( 
.A(n_3983),
.B(n_3937),
.Y(n_4542)
);

INVx2_ASAP7_75t_L g4543 ( 
.A(n_4033),
.Y(n_4543)
);

OAI321xp33_ASAP7_75t_L g4544 ( 
.A1(n_4478),
.A2(n_4474),
.A3(n_4005),
.B1(n_4501),
.B2(n_4124),
.C(n_4133),
.Y(n_4544)
);

AOI22xp5_ASAP7_75t_L g4545 ( 
.A1(n_4433),
.A2(n_3946),
.B1(n_3905),
.B2(n_3906),
.Y(n_4545)
);

AOI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_4313),
.A2(n_3942),
.B(n_3607),
.Y(n_4546)
);

AOI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4280),
.A2(n_3615),
.B(n_3584),
.Y(n_4547)
);

AOI21xp5_ASAP7_75t_L g4548 ( 
.A1(n_4092),
.A2(n_3630),
.B(n_3622),
.Y(n_4548)
);

OAI21xp33_ASAP7_75t_L g4549 ( 
.A1(n_4049),
.A2(n_4137),
.B(n_4486),
.Y(n_4549)
);

NOR2xp33_ASAP7_75t_L g4550 ( 
.A(n_4300),
.B(n_3782),
.Y(n_4550)
);

NAND2x1p5_ASAP7_75t_L g4551 ( 
.A(n_4006),
.B(n_3631),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4033),
.Y(n_4552)
);

AOI22xp5_ASAP7_75t_L g4553 ( 
.A1(n_4436),
.A2(n_3886),
.B1(n_3800),
.B2(n_3808),
.Y(n_4553)
);

AOI21x1_ASAP7_75t_L g4554 ( 
.A1(n_3994),
.A2(n_3639),
.B(n_3637),
.Y(n_4554)
);

AND2x6_ASAP7_75t_L g4555 ( 
.A(n_4259),
.B(n_3502),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4226),
.B(n_152),
.Y(n_4556)
);

BUFx2_ASAP7_75t_L g4557 ( 
.A(n_3987),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4119),
.B(n_3511),
.Y(n_4558)
);

OAI22xp5_ASAP7_75t_L g4559 ( 
.A1(n_4379),
.A2(n_3493),
.B1(n_3809),
.B2(n_3793),
.Y(n_4559)
);

NOR2xp67_ASAP7_75t_L g4560 ( 
.A(n_4006),
.B(n_153),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3988),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_4274),
.B(n_3527),
.Y(n_4562)
);

AOI21xp5_ASAP7_75t_L g4563 ( 
.A1(n_4231),
.A2(n_3677),
.B(n_3647),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_SL g4564 ( 
.A(n_3973),
.B(n_3678),
.Y(n_4564)
);

AOI221xp5_ASAP7_75t_L g4565 ( 
.A1(n_4496),
.A2(n_3532),
.B1(n_3543),
.B2(n_3707),
.C(n_3699),
.Y(n_4565)
);

AOI21x1_ASAP7_75t_L g4566 ( 
.A1(n_4371),
.A2(n_3710),
.B(n_3709),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_4009),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4051),
.Y(n_4568)
);

AOI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_4248),
.A2(n_3731),
.B(n_3727),
.Y(n_4569)
);

NOR2x1_ASAP7_75t_L g4570 ( 
.A(n_3997),
.B(n_154),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4051),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_3970),
.B(n_155),
.Y(n_4572)
);

AND2x4_ASAP7_75t_L g4573 ( 
.A(n_4006),
.B(n_4096),
.Y(n_4573)
);

AOI21xp5_ASAP7_75t_L g4574 ( 
.A1(n_4255),
.A2(n_155),
.B(n_156),
.Y(n_4574)
);

BUFx2_ASAP7_75t_L g4575 ( 
.A(n_4026),
.Y(n_4575)
);

OAI321xp33_ASAP7_75t_L g4576 ( 
.A1(n_3976),
.A2(n_157),
.A3(n_159),
.B1(n_155),
.B2(n_156),
.C(n_158),
.Y(n_4576)
);

BUFx2_ASAP7_75t_L g4577 ( 
.A(n_4026),
.Y(n_4577)
);

OAI21x1_ASAP7_75t_L g4578 ( 
.A1(n_4420),
.A2(n_934),
.B(n_922),
.Y(n_4578)
);

O2A1O1Ixp5_ASAP7_75t_L g4579 ( 
.A1(n_4208),
.A2(n_4521),
.B(n_4504),
.C(n_4427),
.Y(n_4579)
);

O2A1O1Ixp33_ASAP7_75t_SL g4580 ( 
.A1(n_3981),
.A2(n_3992),
.B(n_4028),
.C(n_4044),
.Y(n_4580)
);

AOI21xp5_ASAP7_75t_L g4581 ( 
.A1(n_4074),
.A2(n_156),
.B(n_157),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4093),
.B(n_3993),
.Y(n_4582)
);

NOR2xp33_ASAP7_75t_L g4583 ( 
.A(n_4102),
.B(n_158),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4000),
.B(n_158),
.Y(n_4584)
);

INVx1_ASAP7_75t_SL g4585 ( 
.A(n_4082),
.Y(n_4585)
);

AOI22xp33_ASAP7_75t_L g4586 ( 
.A1(n_4507),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4003),
.B(n_159),
.Y(n_4587)
);

NOR2xp33_ASAP7_75t_L g4588 ( 
.A(n_4032),
.B(n_160),
.Y(n_4588)
);

A2O1A1Ixp33_ASAP7_75t_L g4589 ( 
.A1(n_4167),
.A2(n_4475),
.B(n_4143),
.C(n_4417),
.Y(n_4589)
);

AOI21xp5_ASAP7_75t_L g4590 ( 
.A1(n_4081),
.A2(n_161),
.B(n_162),
.Y(n_4590)
);

INVx1_ASAP7_75t_SL g4591 ( 
.A(n_4015),
.Y(n_4591)
);

AOI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_4101),
.A2(n_162),
.B(n_163),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_SL g4593 ( 
.A(n_4096),
.B(n_163),
.Y(n_4593)
);

INVx2_ASAP7_75t_SL g4594 ( 
.A(n_4197),
.Y(n_4594)
);

AOI21xp33_ASAP7_75t_L g4595 ( 
.A1(n_4516),
.A2(n_163),
.B(n_164),
.Y(n_4595)
);

NOR2xp33_ASAP7_75t_L g4596 ( 
.A(n_4129),
.B(n_4147),
.Y(n_4596)
);

A2O1A1Ixp33_ASAP7_75t_L g4597 ( 
.A1(n_4445),
.A2(n_4503),
.B(n_4424),
.C(n_4472),
.Y(n_4597)
);

NOR2xp33_ASAP7_75t_L g4598 ( 
.A(n_4374),
.B(n_164),
.Y(n_4598)
);

NOR2xp33_ASAP7_75t_L g4599 ( 
.A(n_4191),
.B(n_164),
.Y(n_4599)
);

AOI21xp5_ASAP7_75t_L g4600 ( 
.A1(n_4128),
.A2(n_165),
.B(n_166),
.Y(n_4600)
);

INVx3_ASAP7_75t_L g4601 ( 
.A(n_4096),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4088),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4004),
.Y(n_4603)
);

AOI21xp5_ASAP7_75t_L g4604 ( 
.A1(n_4276),
.A2(n_165),
.B(n_166),
.Y(n_4604)
);

AOI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_4361),
.A2(n_165),
.B(n_167),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_L g4606 ( 
.A(n_4007),
.B(n_167),
.Y(n_4606)
);

INVxp67_ASAP7_75t_L g4607 ( 
.A(n_4299),
.Y(n_4607)
);

AOI22x1_ASAP7_75t_L g4608 ( 
.A1(n_4267),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_4608)
);

AOI21xp5_ASAP7_75t_L g4609 ( 
.A1(n_4113),
.A2(n_168),
.B(n_169),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4016),
.B(n_168),
.Y(n_4610)
);

AOI21xp5_ASAP7_75t_L g4611 ( 
.A1(n_4258),
.A2(n_170),
.B(n_171),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4277),
.B(n_170),
.Y(n_4612)
);

AOI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4439),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_4613)
);

AOI21xp5_ASAP7_75t_L g4614 ( 
.A1(n_4369),
.A2(n_172),
.B(n_173),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4034),
.Y(n_4615)
);

NOR2xp33_ASAP7_75t_L g4616 ( 
.A(n_4142),
.B(n_173),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4046),
.B(n_173),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4054),
.B(n_174),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4056),
.B(n_174),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4019),
.Y(n_4620)
);

AO32x1_ASAP7_75t_L g4621 ( 
.A1(n_4363),
.A2(n_176),
.A3(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_4621)
);

NOR2x1_ASAP7_75t_L g4622 ( 
.A(n_3972),
.B(n_175),
.Y(n_4622)
);

AOI21xp5_ASAP7_75t_L g4623 ( 
.A1(n_4193),
.A2(n_176),
.B(n_177),
.Y(n_4623)
);

OAI22xp5_ASAP7_75t_L g4624 ( 
.A1(n_4404),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_4624)
);

AOI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4199),
.A2(n_178),
.B(n_179),
.Y(n_4625)
);

CKINVDCx10_ASAP7_75t_R g4626 ( 
.A(n_4011),
.Y(n_4626)
);

NOR2xp67_ASAP7_75t_L g4627 ( 
.A(n_4108),
.B(n_178),
.Y(n_4627)
);

NOR2x1_ASAP7_75t_L g4628 ( 
.A(n_4014),
.B(n_179),
.Y(n_4628)
);

NAND3xp33_ASAP7_75t_L g4629 ( 
.A(n_3996),
.B(n_179),
.C(n_180),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_SL g4630 ( 
.A(n_4108),
.B(n_180),
.Y(n_4630)
);

NOR2xp33_ASAP7_75t_L g4631 ( 
.A(n_4148),
.B(n_180),
.Y(n_4631)
);

CKINVDCx20_ASAP7_75t_R g4632 ( 
.A(n_4197),
.Y(n_4632)
);

OAI21x1_ASAP7_75t_L g4633 ( 
.A1(n_3986),
.A2(n_924),
.B(n_915),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_L g4634 ( 
.A(n_4061),
.B(n_181),
.Y(n_4634)
);

HB1xp67_ASAP7_75t_L g4635 ( 
.A(n_4027),
.Y(n_4635)
);

NOR2xp33_ASAP7_75t_L g4636 ( 
.A(n_4151),
.B(n_181),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_SL g4637 ( 
.A(n_4108),
.B(n_182),
.Y(n_4637)
);

OAI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_4339),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_4638)
);

AOI21xp5_ASAP7_75t_L g4639 ( 
.A1(n_4211),
.A2(n_183),
.B(n_184),
.Y(n_4639)
);

AOI22x1_ASAP7_75t_L g4640 ( 
.A1(n_4047),
.A2(n_4372),
.B1(n_4024),
.B2(n_4178),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_SL g4641 ( 
.A(n_4173),
.B(n_183),
.Y(n_4641)
);

HB1xp67_ASAP7_75t_L g4642 ( 
.A(n_4298),
.Y(n_4642)
);

OAI21xp33_ASAP7_75t_L g4643 ( 
.A1(n_4440),
.A2(n_4448),
.B(n_4409),
.Y(n_4643)
);

A2O1A1Ixp33_ASAP7_75t_L g4644 ( 
.A1(n_4230),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4067),
.B(n_186),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4069),
.B(n_186),
.Y(n_4646)
);

NOR2xp33_ASAP7_75t_L g4647 ( 
.A(n_4526),
.B(n_187),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4213),
.A2(n_187),
.B(n_188),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4071),
.B(n_187),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4084),
.B(n_4090),
.Y(n_4650)
);

BUFx3_ASAP7_75t_L g4651 ( 
.A(n_4011),
.Y(n_4651)
);

O2A1O1Ixp33_ASAP7_75t_L g4652 ( 
.A1(n_4497),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_4652)
);

AOI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4214),
.A2(n_188),
.B(n_189),
.Y(n_4653)
);

AOI21xp5_ASAP7_75t_L g4654 ( 
.A1(n_4413),
.A2(n_189),
.B(n_190),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_3974),
.Y(n_4655)
);

AOI22xp5_ASAP7_75t_L g4656 ( 
.A1(n_4439),
.A2(n_194),
.B1(n_191),
.B2(n_192),
.Y(n_4656)
);

AOI22xp5_ASAP7_75t_L g4657 ( 
.A1(n_4439),
.A2(n_194),
.B1(n_191),
.B2(n_192),
.Y(n_4657)
);

INVx3_ASAP7_75t_L g4658 ( 
.A(n_4173),
.Y(n_4658)
);

AOI22x1_ASAP7_75t_L g4659 ( 
.A1(n_4053),
.A2(n_195),
.B1(n_191),
.B2(n_194),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4111),
.B(n_195),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4035),
.B(n_196),
.Y(n_4661)
);

AOI21xp5_ASAP7_75t_L g4662 ( 
.A1(n_4086),
.A2(n_196),
.B(n_197),
.Y(n_4662)
);

BUFx6f_ASAP7_75t_L g4663 ( 
.A(n_4173),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4279),
.B(n_4138),
.Y(n_4664)
);

NOR2xp33_ASAP7_75t_L g4665 ( 
.A(n_4282),
.B(n_197),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4149),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4156),
.B(n_197),
.Y(n_4667)
);

AOI21xp5_ASAP7_75t_L g4668 ( 
.A1(n_4348),
.A2(n_198),
.B(n_199),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_L g4669 ( 
.A(n_4159),
.B(n_198),
.Y(n_4669)
);

O2A1O1Ixp33_ASAP7_75t_L g4670 ( 
.A1(n_4502),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_4670)
);

AOI21xp5_ASAP7_75t_L g4671 ( 
.A1(n_4370),
.A2(n_199),
.B(n_200),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4172),
.B(n_200),
.Y(n_4672)
);

A2O1A1Ixp33_ASAP7_75t_L g4673 ( 
.A1(n_4378),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_4673)
);

A2O1A1Ixp33_ASAP7_75t_L g4674 ( 
.A1(n_4477),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4174),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4180),
.Y(n_4676)
);

OAI21xp5_ASAP7_75t_L g4677 ( 
.A1(n_4527),
.A2(n_201),
.B(n_202),
.Y(n_4677)
);

AOI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_4373),
.A2(n_204),
.B(n_205),
.Y(n_4678)
);

NOR2xp67_ASAP7_75t_L g4679 ( 
.A(n_4198),
.B(n_204),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4321),
.B(n_204),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4352),
.A2(n_206),
.B(n_207),
.Y(n_4681)
);

AOI21xp5_ASAP7_75t_L g4682 ( 
.A1(n_4179),
.A2(n_207),
.B(n_208),
.Y(n_4682)
);

OAI22xp5_ASAP7_75t_L g4683 ( 
.A1(n_4243),
.A2(n_210),
.B1(n_207),
.B2(n_209),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4181),
.Y(n_4684)
);

AOI21xp5_ASAP7_75t_L g4685 ( 
.A1(n_4287),
.A2(n_209),
.B(n_210),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4217),
.B(n_4223),
.Y(n_4686)
);

AOI21xp5_ASAP7_75t_L g4687 ( 
.A1(n_4295),
.A2(n_209),
.B(n_210),
.Y(n_4687)
);

NOR2xp33_ASAP7_75t_L g4688 ( 
.A(n_4055),
.B(n_211),
.Y(n_4688)
);

OAI21xp5_ASAP7_75t_L g4689 ( 
.A1(n_4456),
.A2(n_212),
.B(n_213),
.Y(n_4689)
);

AOI21xp5_ASAP7_75t_L g4690 ( 
.A1(n_4017),
.A2(n_212),
.B(n_213),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_3980),
.Y(n_4691)
);

AOI21xp5_ASAP7_75t_L g4692 ( 
.A1(n_4322),
.A2(n_212),
.B(n_214),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4327),
.B(n_4329),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_4228),
.B(n_214),
.Y(n_4694)
);

AOI21xp5_ASAP7_75t_L g4695 ( 
.A1(n_4141),
.A2(n_215),
.B(n_216),
.Y(n_4695)
);

OA22x2_ASAP7_75t_L g4696 ( 
.A1(n_4094),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_4696)
);

NOR2xp33_ASAP7_75t_L g4697 ( 
.A(n_4196),
.B(n_216),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4232),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4242),
.Y(n_4699)
);

NAND2x1_ASAP7_75t_L g4700 ( 
.A(n_4219),
.B(n_217),
.Y(n_4700)
);

NOR2xp67_ASAP7_75t_L g4701 ( 
.A(n_4198),
.B(n_218),
.Y(n_4701)
);

NOR3xp33_ASAP7_75t_L g4702 ( 
.A(n_4291),
.B(n_227),
.C(n_219),
.Y(n_4702)
);

AOI21xp5_ASAP7_75t_L g4703 ( 
.A1(n_4154),
.A2(n_220),
.B(n_221),
.Y(n_4703)
);

AOI21x1_ASAP7_75t_L g4704 ( 
.A1(n_4162),
.A2(n_220),
.B(n_221),
.Y(n_4704)
);

AOI21xp5_ASAP7_75t_L g4705 ( 
.A1(n_4163),
.A2(n_221),
.B(n_222),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4256),
.B(n_4264),
.Y(n_4706)
);

OAI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4323),
.A2(n_222),
.B(n_223),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4269),
.B(n_222),
.Y(n_4708)
);

A2O1A1Ixp33_ASAP7_75t_L g4709 ( 
.A1(n_4125),
.A2(n_4045),
.B(n_4512),
.C(n_4428),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4281),
.B(n_223),
.Y(n_4710)
);

O2A1O1Ixp5_ASAP7_75t_L g4711 ( 
.A1(n_4395),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_4711)
);

CKINVDCx8_ASAP7_75t_R g4712 ( 
.A(n_4050),
.Y(n_4712)
);

AOI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4164),
.A2(n_224),
.B(n_225),
.Y(n_4713)
);

AOI21xp5_ASAP7_75t_L g4714 ( 
.A1(n_3977),
.A2(n_225),
.B(n_226),
.Y(n_4714)
);

AOI22xp33_ASAP7_75t_L g4715 ( 
.A1(n_4438),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_L g4716 ( 
.A(n_4303),
.B(n_226),
.Y(n_4716)
);

O2A1O1Ixp33_ASAP7_75t_L g4717 ( 
.A1(n_4534),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4306),
.B(n_228),
.Y(n_4718)
);

O2A1O1Ixp33_ASAP7_75t_SL g4719 ( 
.A1(n_4018),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_4719)
);

NOR2xp33_ASAP7_75t_L g4720 ( 
.A(n_4309),
.B(n_230),
.Y(n_4720)
);

AOI21xp5_ASAP7_75t_L g4721 ( 
.A1(n_4402),
.A2(n_231),
.B(n_232),
.Y(n_4721)
);

O2A1O1Ixp33_ASAP7_75t_L g4722 ( 
.A1(n_4118),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_4722)
);

AOI21xp5_ASAP7_75t_L g4723 ( 
.A1(n_3971),
.A2(n_233),
.B(n_234),
.Y(n_4723)
);

OAI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_4233),
.A2(n_236),
.B(n_237),
.Y(n_4724)
);

INVx3_ASAP7_75t_L g4725 ( 
.A(n_4198),
.Y(n_4725)
);

OAI22x1_ASAP7_75t_L g4726 ( 
.A1(n_4237),
.A2(n_3999),
.B1(n_4070),
.B2(n_4123),
.Y(n_4726)
);

AND2x2_ASAP7_75t_L g4727 ( 
.A(n_4331),
.B(n_236),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4307),
.B(n_236),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4318),
.B(n_237),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4200),
.B(n_237),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4330),
.B(n_238),
.Y(n_4731)
);

NOR2xp33_ASAP7_75t_L g4732 ( 
.A(n_4296),
.B(n_4301),
.Y(n_4732)
);

INVx1_ASAP7_75t_SL g4733 ( 
.A(n_4254),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_L g4734 ( 
.A(n_4319),
.B(n_238),
.Y(n_4734)
);

BUFx3_ASAP7_75t_L g4735 ( 
.A(n_4077),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_L g4736 ( 
.A(n_4454),
.B(n_238),
.Y(n_4736)
);

OAI22xp5_ASAP7_75t_L g4737 ( 
.A1(n_4253),
.A2(n_4002),
.B1(n_4171),
.B2(n_4209),
.Y(n_4737)
);

CKINVDCx10_ASAP7_75t_R g4738 ( 
.A(n_4203),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_4468),
.B(n_239),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_SL g4740 ( 
.A(n_4446),
.B(n_239),
.Y(n_4740)
);

AND2x6_ASAP7_75t_L g4741 ( 
.A(n_4347),
.B(n_239),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4324),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4132),
.Y(n_4743)
);

O2A1O1Ixp33_ASAP7_75t_L g4744 ( 
.A1(n_4010),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4360),
.B(n_240),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_SL g4746 ( 
.A(n_4446),
.B(n_240),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_4377),
.A2(n_241),
.B(n_243),
.Y(n_4747)
);

OAI22xp5_ASAP7_75t_L g4748 ( 
.A1(n_4335),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_SL g4749 ( 
.A(n_4446),
.B(n_243),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4136),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4396),
.B(n_244),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4362),
.B(n_244),
.Y(n_4752)
);

OAI22xp5_ASAP7_75t_L g4753 ( 
.A1(n_4185),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_4753)
);

AOI21xp5_ASAP7_75t_L g4754 ( 
.A1(n_4271),
.A2(n_246),
.B(n_247),
.Y(n_4754)
);

OAI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_4471),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_4755)
);

INVxp67_ASAP7_75t_SL g4756 ( 
.A(n_4342),
.Y(n_4756)
);

AO21x1_ASAP7_75t_L g4757 ( 
.A1(n_4384),
.A2(n_248),
.B(n_249),
.Y(n_4757)
);

AOI21x1_ASAP7_75t_L g4758 ( 
.A1(n_3986),
.A2(n_249),
.B(n_250),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4364),
.B(n_250),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4366),
.B(n_251),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4367),
.B(n_251),
.Y(n_4761)
);

AOI21xp5_ASAP7_75t_L g4762 ( 
.A1(n_4412),
.A2(n_252),
.B(n_253),
.Y(n_4762)
);

AOI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4235),
.A2(n_4272),
.B(n_4031),
.Y(n_4763)
);

OAI22xp5_ASAP7_75t_L g4764 ( 
.A1(n_4482),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_4764)
);

AOI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4399),
.A2(n_253),
.B(n_254),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_4060),
.Y(n_4766)
);

AOI21xp5_ASAP7_75t_L g4767 ( 
.A1(n_4421),
.A2(n_254),
.B(n_255),
.Y(n_4767)
);

AOI21x1_ASAP7_75t_L g4768 ( 
.A1(n_4394),
.A2(n_256),
.B(n_257),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4375),
.B(n_256),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4315),
.A2(n_257),
.B(n_258),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4380),
.B(n_257),
.Y(n_4771)
);

INVxp67_ASAP7_75t_L g4772 ( 
.A(n_4192),
.Y(n_4772)
);

AOI21x1_ASAP7_75t_L g4773 ( 
.A1(n_4394),
.A2(n_258),
.B(n_259),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4350),
.B(n_258),
.Y(n_4774)
);

A2O1A1Ixp33_ASAP7_75t_L g4775 ( 
.A1(n_4459),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_4775)
);

OAI21xp5_ASAP7_75t_L g4776 ( 
.A1(n_4022),
.A2(n_260),
.B(n_261),
.Y(n_4776)
);

AOI21xp5_ASAP7_75t_L g4777 ( 
.A1(n_4328),
.A2(n_4344),
.B(n_4357),
.Y(n_4777)
);

AOI21xp5_ASAP7_75t_L g4778 ( 
.A1(n_3982),
.A2(n_261),
.B(n_262),
.Y(n_4778)
);

A2O1A1Ixp33_ASAP7_75t_L g4779 ( 
.A1(n_4065),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_4779)
);

OAI21x1_ASAP7_75t_L g4780 ( 
.A1(n_4079),
.A2(n_931),
.B(n_917),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_3985),
.Y(n_4781)
);

O2A1O1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_4506),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4389),
.B(n_263),
.Y(n_4783)
);

O2A1O1Ixp33_ASAP7_75t_L g4784 ( 
.A1(n_4207),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_4784)
);

AOI21xp5_ASAP7_75t_L g4785 ( 
.A1(n_3982),
.A2(n_266),
.B(n_267),
.Y(n_4785)
);

NOR2xp33_ASAP7_75t_R g4786 ( 
.A(n_4020),
.B(n_267),
.Y(n_4786)
);

NOR2xp33_ASAP7_75t_L g4787 ( 
.A(n_4418),
.B(n_267),
.Y(n_4787)
);

AOI21xp5_ASAP7_75t_L g4788 ( 
.A1(n_3989),
.A2(n_268),
.B(n_269),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_SL g4789 ( 
.A(n_4285),
.B(n_268),
.Y(n_4789)
);

NOR2xp67_ASAP7_75t_L g4790 ( 
.A(n_4221),
.B(n_4239),
.Y(n_4790)
);

INVx1_ASAP7_75t_SL g4791 ( 
.A(n_4150),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4400),
.B(n_268),
.Y(n_4792)
);

NOR2xp33_ASAP7_75t_L g4793 ( 
.A(n_4161),
.B(n_269),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4401),
.B(n_269),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4336),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4406),
.B(n_270),
.Y(n_4796)
);

AOI21xp5_ASAP7_75t_L g4797 ( 
.A1(n_3989),
.A2(n_270),
.B(n_271),
.Y(n_4797)
);

A2O1A1Ixp33_ASAP7_75t_L g4798 ( 
.A1(n_4457),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_4798)
);

INVxp67_ASAP7_75t_L g4799 ( 
.A(n_4059),
.Y(n_4799)
);

BUFx3_ASAP7_75t_L g4800 ( 
.A(n_4073),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_SL g4801 ( 
.A(n_4285),
.B(n_272),
.Y(n_4801)
);

INVx2_ASAP7_75t_SL g4802 ( 
.A(n_4062),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4425),
.B(n_273),
.Y(n_4803)
);

INVx11_ASAP7_75t_L g4804 ( 
.A(n_3975),
.Y(n_4804)
);

OAI21x1_ASAP7_75t_SL g4805 ( 
.A1(n_4343),
.A2(n_273),
.B(n_274),
.Y(n_4805)
);

NOR2xp33_ASAP7_75t_L g4806 ( 
.A(n_4117),
.B(n_274),
.Y(n_4806)
);

OAI22xp5_ASAP7_75t_L g4807 ( 
.A1(n_4457),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4430),
.B(n_4443),
.Y(n_4808)
);

NAND3xp33_ASAP7_75t_L g4809 ( 
.A(n_4206),
.B(n_275),
.C(n_276),
.Y(n_4809)
);

OAI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4465),
.A2(n_275),
.B(n_277),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4444),
.B(n_277),
.Y(n_4811)
);

AOI21xp5_ASAP7_75t_L g4812 ( 
.A1(n_4218),
.A2(n_278),
.B(n_279),
.Y(n_4812)
);

AOI21xp5_ASAP7_75t_L g4813 ( 
.A1(n_4218),
.A2(n_279),
.B(n_280),
.Y(n_4813)
);

NAND3xp33_ASAP7_75t_L g4814 ( 
.A(n_4529),
.B(n_279),
.C(n_280),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4382),
.B(n_281),
.Y(n_4815)
);

AOI22xp33_ASAP7_75t_L g4816 ( 
.A1(n_4442),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_4816)
);

OAI22xp5_ASAP7_75t_L g4817 ( 
.A1(n_4462),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_SL g4818 ( 
.A(n_4285),
.B(n_283),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_4405),
.B(n_284),
.Y(n_4819)
);

BUFx3_ASAP7_75t_L g4820 ( 
.A(n_4039),
.Y(n_4820)
);

NOR2xp33_ASAP7_75t_L g4821 ( 
.A(n_4160),
.B(n_287),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4479),
.B(n_287),
.Y(n_4822)
);

AOI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4466),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_4823)
);

OAI22xp5_ASAP7_75t_L g4824 ( 
.A1(n_4462),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_4824)
);

O2A1O1Ixp33_ASAP7_75t_L g4825 ( 
.A1(n_4490),
.A2(n_292),
.B(n_289),
.C(n_291),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4481),
.B(n_291),
.Y(n_4826)
);

O2A1O1Ixp33_ASAP7_75t_SL g4827 ( 
.A1(n_4455),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_SL g4828 ( 
.A(n_4285),
.B(n_292),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_L g4829 ( 
.A(n_4488),
.B(n_293),
.Y(n_4829)
);

BUFx4f_ASAP7_75t_L g4830 ( 
.A(n_4012),
.Y(n_4830)
);

BUFx2_ASAP7_75t_L g4831 ( 
.A(n_3979),
.Y(n_4831)
);

NOR2xp33_ASAP7_75t_L g4832 ( 
.A(n_4135),
.B(n_293),
.Y(n_4832)
);

AND2x2_ASAP7_75t_L g4833 ( 
.A(n_4414),
.B(n_294),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4227),
.A2(n_294),
.B(n_295),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4097),
.B(n_295),
.Y(n_4835)
);

NAND3xp33_ASAP7_75t_SL g4836 ( 
.A(n_4449),
.B(n_295),
.C(n_296),
.Y(n_4836)
);

BUFx5_ASAP7_75t_L g4837 ( 
.A(n_4089),
.Y(n_4837)
);

OAI22xp5_ASAP7_75t_L g4838 ( 
.A1(n_4518),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_4838)
);

OAI22xp5_ASAP7_75t_L g4839 ( 
.A1(n_4518),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_4839)
);

NAND3xp33_ASAP7_75t_L g4840 ( 
.A(n_4535),
.B(n_297),
.C(n_298),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4337),
.Y(n_4841)
);

OAI22xp5_ASAP7_75t_L g4842 ( 
.A1(n_4043),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_4842)
);

OAI22xp5_ASAP7_75t_L g4843 ( 
.A1(n_4434),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_4523),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_4844)
);

AOI21xp5_ASAP7_75t_L g4845 ( 
.A1(n_4227),
.A2(n_302),
.B(n_303),
.Y(n_4845)
);

O2A1O1Ixp33_ASAP7_75t_L g4846 ( 
.A1(n_4500),
.A2(n_4398),
.B(n_4407),
.C(n_4393),
.Y(n_4846)
);

AOI21xp5_ASAP7_75t_L g4847 ( 
.A1(n_4261),
.A2(n_303),
.B(n_304),
.Y(n_4847)
);

INVx11_ASAP7_75t_L g4848 ( 
.A(n_4476),
.Y(n_4848)
);

INVx4_ASAP7_75t_L g4849 ( 
.A(n_4221),
.Y(n_4849)
);

HB1xp67_ASAP7_75t_L g4850 ( 
.A(n_4216),
.Y(n_4850)
);

AND2x4_ASAP7_75t_L g4851 ( 
.A(n_4221),
.B(n_304),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4495),
.B(n_305),
.Y(n_4852)
);

O2A1O1Ixp33_ASAP7_75t_SL g4853 ( 
.A1(n_4470),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4451),
.B(n_305),
.Y(n_4854)
);

OAI21xp5_ASAP7_75t_L g4855 ( 
.A1(n_4485),
.A2(n_306),
.B(n_307),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4338),
.B(n_307),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4340),
.Y(n_4857)
);

INVx1_ASAP7_75t_SL g4858 ( 
.A(n_4052),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4261),
.A2(n_308),
.B(n_309),
.Y(n_4859)
);

INVx1_ASAP7_75t_SL g4860 ( 
.A(n_4107),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4131),
.B(n_308),
.Y(n_4861)
);

AOI21xp5_ASAP7_75t_L g4862 ( 
.A1(n_4416),
.A2(n_308),
.B(n_309),
.Y(n_4862)
);

OA22x2_ASAP7_75t_L g4863 ( 
.A1(n_4085),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_4863)
);

O2A1O1Ixp5_ASAP7_75t_L g4864 ( 
.A1(n_4514),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_4864)
);

NAND3xp33_ASAP7_75t_L g4865 ( 
.A(n_4484),
.B(n_310),
.C(n_311),
.Y(n_4865)
);

BUFx6f_ASAP7_75t_L g4866 ( 
.A(n_4057),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_SL g4867 ( 
.A(n_4365),
.B(n_313),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_L g4868 ( 
.A(n_4426),
.B(n_313),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4453),
.B(n_314),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4063),
.Y(n_4870)
);

A2O1A1Ixp33_ASAP7_75t_L g4871 ( 
.A1(n_4353),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_4871)
);

AO22x1_ASAP7_75t_L g4872 ( 
.A1(n_4080),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_4872)
);

AOI21xp5_ASAP7_75t_L g4873 ( 
.A1(n_4416),
.A2(n_315),
.B(n_317),
.Y(n_4873)
);

AOI21x1_ASAP7_75t_L g4874 ( 
.A1(n_4041),
.A2(n_317),
.B(n_318),
.Y(n_4874)
);

AOI21xp5_ASAP7_75t_L g4875 ( 
.A1(n_4422),
.A2(n_317),
.B(n_319),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4473),
.B(n_319),
.Y(n_4876)
);

OAI22xp5_ASAP7_75t_L g4877 ( 
.A1(n_4434),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4877)
);

AOI21xp5_ASAP7_75t_L g4878 ( 
.A1(n_4422),
.A2(n_320),
.B(n_321),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_L g4879 ( 
.A(n_4157),
.B(n_322),
.Y(n_4879)
);

NOR2xp67_ASAP7_75t_L g4880 ( 
.A(n_4239),
.B(n_4058),
.Y(n_4880)
);

AOI21xp5_ASAP7_75t_L g4881 ( 
.A1(n_4408),
.A2(n_322),
.B(n_323),
.Y(n_4881)
);

AOI22x1_ASAP7_75t_L g4882 ( 
.A1(n_4316),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4508),
.B(n_4510),
.Y(n_4883)
);

OAI22xp5_ASAP7_75t_L g4884 ( 
.A1(n_4359),
.A2(n_327),
.B1(n_323),
.B2(n_326),
.Y(n_4884)
);

OAI21xp5_ASAP7_75t_L g4885 ( 
.A1(n_4487),
.A2(n_326),
.B(n_327),
.Y(n_4885)
);

INVx3_ASAP7_75t_L g4886 ( 
.A(n_4089),
.Y(n_4886)
);

AND2x2_ASAP7_75t_SL g4887 ( 
.A(n_4210),
.B(n_326),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_SL g4888 ( 
.A(n_4250),
.B(n_327),
.Y(n_4888)
);

OAI22xp5_ASAP7_75t_L g4889 ( 
.A1(n_4127),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_4889)
);

NAND2xp33_ASAP7_75t_L g4890 ( 
.A(n_4166),
.B(n_329),
.Y(n_4890)
);

NOR2xp33_ASAP7_75t_SL g4891 ( 
.A(n_4203),
.B(n_4249),
.Y(n_4891)
);

AOI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4381),
.A2(n_4351),
.B(n_4013),
.Y(n_4892)
);

AOI22xp5_ASAP7_75t_L g4893 ( 
.A1(n_4001),
.A2(n_333),
.B1(n_330),
.B2(n_331),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4037),
.B(n_4040),
.Y(n_4894)
);

HB1xp67_ASAP7_75t_L g4895 ( 
.A(n_3991),
.Y(n_4895)
);

NOR2xp33_ASAP7_75t_L g4896 ( 
.A(n_4410),
.B(n_331),
.Y(n_4896)
);

A2O1A1Ixp33_ASAP7_75t_L g4897 ( 
.A1(n_4467),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_4897)
);

AOI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4498),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4517),
.B(n_4432),
.Y(n_4899)
);

OAI22xp5_ASAP7_75t_L g4900 ( 
.A1(n_4222),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_4900)
);

O2A1O1Ixp5_ASAP7_75t_L g4901 ( 
.A1(n_4505),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_4901)
);

INVx2_ASAP7_75t_L g4902 ( 
.A(n_4023),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4144),
.A2(n_337),
.B(n_338),
.Y(n_4903)
);

NAND3xp33_ASAP7_75t_L g4904 ( 
.A(n_4489),
.B(n_337),
.C(n_339),
.Y(n_4904)
);

INVx5_ASAP7_75t_L g4905 ( 
.A(n_4249),
.Y(n_4905)
);

AND2x4_ASAP7_75t_L g4906 ( 
.A(n_4239),
.B(n_339),
.Y(n_4906)
);

O2A1O1Ixp5_ASAP7_75t_L g4907 ( 
.A1(n_4441),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4152),
.A2(n_340),
.B(n_341),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4435),
.B(n_342),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4341),
.Y(n_4910)
);

AOI22x1_ASAP7_75t_L g4911 ( 
.A1(n_4515),
.A2(n_4356),
.B1(n_4297),
.B2(n_4294),
.Y(n_4911)
);

AOI21x1_ASAP7_75t_L g4912 ( 
.A1(n_4392),
.A2(n_4447),
.B(n_3990),
.Y(n_4912)
);

OAI21x1_ASAP7_75t_L g4913 ( 
.A1(n_4284),
.A2(n_935),
.B(n_921),
.Y(n_4913)
);

AOI22xp5_ASAP7_75t_L g4914 ( 
.A1(n_4078),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4345),
.Y(n_4915)
);

OAI22x1_ASAP7_75t_L g4916 ( 
.A1(n_4265),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4452),
.B(n_343),
.Y(n_4917)
);

AOI21xp5_ASAP7_75t_L g4918 ( 
.A1(n_4305),
.A2(n_344),
.B(n_345),
.Y(n_4918)
);

AOI21xp5_ASAP7_75t_L g4919 ( 
.A1(n_4025),
.A2(n_346),
.B(n_347),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_4029),
.A2(n_346),
.B(n_347),
.Y(n_4920)
);

OR2x2_ASAP7_75t_L g4921 ( 
.A(n_4415),
.B(n_346),
.Y(n_4921)
);

BUFx2_ASAP7_75t_SL g4922 ( 
.A(n_4219),
.Y(n_4922)
);

O2A1O1Ixp33_ASAP7_75t_L g4923 ( 
.A1(n_4429),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_4923)
);

AOI21xp5_ASAP7_75t_L g4924 ( 
.A1(n_4036),
.A2(n_348),
.B(n_349),
.Y(n_4924)
);

NOR2xp33_ASAP7_75t_L g4925 ( 
.A(n_4109),
.B(n_348),
.Y(n_4925)
);

NOR2xp33_ASAP7_75t_L g4926 ( 
.A(n_4121),
.B(n_350),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4064),
.Y(n_4927)
);

A2O1A1Ixp33_ASAP7_75t_L g4928 ( 
.A1(n_4289),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_4928)
);

AOI21xp5_ASAP7_75t_L g4929 ( 
.A1(n_4083),
.A2(n_351),
.B(n_352),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_SL g4930 ( 
.A(n_4250),
.B(n_351),
.Y(n_4930)
);

BUFx12f_ASAP7_75t_L g4931 ( 
.A(n_4008),
.Y(n_4931)
);

OAI22xp5_ASAP7_75t_SL g4932 ( 
.A1(n_4292),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_4932)
);

OR2x2_ASAP7_75t_L g4933 ( 
.A(n_4104),
.B(n_353),
.Y(n_4933)
);

AOI21xp5_ASAP7_75t_L g4934 ( 
.A1(n_4120),
.A2(n_353),
.B(n_354),
.Y(n_4934)
);

AOI221xp5_ASAP7_75t_L g4935 ( 
.A1(n_3998),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.C(n_358),
.Y(n_4935)
);

OAI21xp5_ASAP7_75t_L g4936 ( 
.A1(n_4494),
.A2(n_4513),
.B(n_4383),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4483),
.B(n_355),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_SL g4938 ( 
.A1(n_4189),
.A2(n_355),
.B(n_356),
.Y(n_4938)
);

AOI22xp5_ASAP7_75t_L g4939 ( 
.A1(n_4493),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_4939)
);

AOI21xp5_ASAP7_75t_L g4940 ( 
.A1(n_4511),
.A2(n_357),
.B(n_358),
.Y(n_4940)
);

INVx3_ASAP7_75t_L g4941 ( 
.A(n_4089),
.Y(n_4941)
);

BUFx4f_ASAP7_75t_L g4942 ( 
.A(n_4189),
.Y(n_4942)
);

NAND3xp33_ASAP7_75t_L g4943 ( 
.A(n_4458),
.B(n_359),
.C(n_360),
.Y(n_4943)
);

NOR3xp33_ASAP7_75t_L g4944 ( 
.A(n_4463),
.B(n_368),
.C(n_359),
.Y(n_4944)
);

AOI21xp5_ASAP7_75t_L g4945 ( 
.A1(n_4520),
.A2(n_360),
.B(n_361),
.Y(n_4945)
);

OAI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4368),
.A2(n_360),
.B(n_361),
.Y(n_4946)
);

OAI21xp5_ASAP7_75t_L g4947 ( 
.A1(n_4385),
.A2(n_361),
.B(n_362),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_4499),
.B(n_362),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4158),
.Y(n_4949)
);

NOR2xp67_ASAP7_75t_L g4950 ( 
.A(n_4139),
.B(n_363),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_4170),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_3978),
.B(n_363),
.Y(n_4952)
);

O2A1O1Ixp33_ASAP7_75t_SL g4953 ( 
.A1(n_4205),
.A2(n_367),
.B(n_364),
.C(n_366),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_SL g4954 ( 
.A(n_4250),
.B(n_364),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_SL g4955 ( 
.A(n_3990),
.B(n_367),
.Y(n_4955)
);

CKINVDCx10_ASAP7_75t_R g4956 ( 
.A(n_4038),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4460),
.B(n_367),
.Y(n_4957)
);

AOI21xp5_ASAP7_75t_L g4958 ( 
.A1(n_4531),
.A2(n_368),
.B(n_369),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4450),
.B(n_368),
.Y(n_4959)
);

INVx2_ASAP7_75t_SL g4960 ( 
.A(n_4168),
.Y(n_4960)
);

INVx4_ASAP7_75t_L g4961 ( 
.A(n_4219),
.Y(n_4961)
);

A2O1A1Ixp33_ASAP7_75t_L g4962 ( 
.A1(n_4186),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_L g4963 ( 
.A(n_4530),
.B(n_370),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_SL g4964 ( 
.A(n_4266),
.B(n_370),
.Y(n_4964)
);

NAND2xp5_ASAP7_75t_L g4965 ( 
.A(n_4532),
.B(n_371),
.Y(n_4965)
);

O2A1O1Ixp33_ASAP7_75t_SL g4966 ( 
.A1(n_4238),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_4966)
);

NAND2xp33_ASAP7_75t_L g4967 ( 
.A(n_4098),
.B(n_373),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4115),
.B(n_373),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4183),
.B(n_374),
.Y(n_4969)
);

AOI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4190),
.A2(n_374),
.B(n_375),
.Y(n_4970)
);

CKINVDCx5p33_ASAP7_75t_R g4971 ( 
.A(n_4334),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4187),
.B(n_375),
.Y(n_4972)
);

NOR2xp33_ASAP7_75t_L g4973 ( 
.A(n_4175),
.B(n_375),
.Y(n_4973)
);

AOI21x1_ASAP7_75t_L g4974 ( 
.A1(n_3995),
.A2(n_376),
.B(n_378),
.Y(n_4974)
);

AOI221xp5_ASAP7_75t_L g4975 ( 
.A1(n_4437),
.A2(n_380),
.B1(n_376),
.B2(n_379),
.C(n_381),
.Y(n_4975)
);

BUFx6f_ASAP7_75t_L g4976 ( 
.A(n_4057),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4087),
.B(n_4397),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4215),
.B(n_376),
.Y(n_4978)
);

OAI22xp5_ASAP7_75t_L g4979 ( 
.A1(n_4212),
.A2(n_4461),
.B1(n_4201),
.B2(n_4134),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4244),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4246),
.Y(n_4981)
);

A2O1A1Ixp33_ASAP7_75t_L g4982 ( 
.A1(n_4106),
.A2(n_381),
.B(n_379),
.C(n_380),
.Y(n_4982)
);

OR2x2_ASAP7_75t_SL g4983 ( 
.A(n_4075),
.B(n_379),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_SL g4984 ( 
.A(n_4528),
.B(n_380),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4403),
.B(n_382),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4251),
.A2(n_382),
.B(n_383),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_4252),
.A2(n_383),
.B(n_384),
.Y(n_4987)
);

O2A1O1Ixp5_ASAP7_75t_L g4988 ( 
.A1(n_4388),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_4988)
);

O2A1O1Ixp33_ASAP7_75t_SL g4989 ( 
.A1(n_4241),
.A2(n_4245),
.B(n_4354),
.C(n_4095),
.Y(n_4989)
);

AOI21xp5_ASAP7_75t_L g4990 ( 
.A1(n_4257),
.A2(n_384),
.B(n_385),
.Y(n_4990)
);

OAI22xp5_ASAP7_75t_L g4991 ( 
.A1(n_4325),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4278),
.A2(n_387),
.B(n_388),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4290),
.B(n_387),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4308),
.A2(n_388),
.B(n_389),
.Y(n_4994)
);

AOI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4310),
.A2(n_389),
.B(n_390),
.Y(n_4995)
);

OAI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4492),
.A2(n_4464),
.B(n_4184),
.Y(n_4996)
);

INVx4_ASAP7_75t_L g4997 ( 
.A(n_4146),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4312),
.B(n_390),
.Y(n_4998)
);

BUFx8_ASAP7_75t_L g4999 ( 
.A(n_4262),
.Y(n_4999)
);

BUFx6f_ASAP7_75t_SL g5000 ( 
.A(n_4234),
.Y(n_5000)
);

OAI22xp5_ASAP7_75t_L g5001 ( 
.A1(n_4325),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_5001)
);

O2A1O1Ixp5_ASAP7_75t_L g5002 ( 
.A1(n_4202),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_5002)
);

OAI22xp5_ASAP7_75t_L g5003 ( 
.A1(n_4469),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4317),
.A2(n_393),
.B(n_394),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4320),
.B(n_394),
.Y(n_5005)
);

INVx3_ASAP7_75t_L g5006 ( 
.A(n_4146),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4326),
.B(n_395),
.Y(n_5007)
);

A2O1A1Ixp33_ASAP7_75t_L g5008 ( 
.A1(n_4188),
.A2(n_398),
.B(n_396),
.C(n_397),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4346),
.B(n_396),
.Y(n_5009)
);

AOI21xp33_ASAP7_75t_L g5010 ( 
.A1(n_4549),
.A2(n_4491),
.B(n_4524),
.Y(n_5010)
);

NAND2x1p5_ASAP7_75t_L g5011 ( 
.A(n_4942),
.B(n_4195),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4742),
.B(n_4431),
.Y(n_5012)
);

OAI21x1_ASAP7_75t_L g5013 ( 
.A1(n_4758),
.A2(n_4286),
.B(n_4204),
.Y(n_5013)
);

INVx4_ASAP7_75t_L g5014 ( 
.A(n_4942),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4561),
.Y(n_5015)
);

OAI21x1_ASAP7_75t_L g5016 ( 
.A1(n_4633),
.A2(n_4332),
.B(n_4314),
.Y(n_5016)
);

AOI21x1_ASAP7_75t_SL g5017 ( 
.A1(n_4851),
.A2(n_4105),
.B(n_4100),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4756),
.B(n_4229),
.Y(n_5018)
);

OA21x2_ASAP7_75t_L g5019 ( 
.A1(n_4777),
.A2(n_4155),
.B(n_4333),
.Y(n_5019)
);

AND2x2_ASAP7_75t_L g5020 ( 
.A(n_4894),
.B(n_4288),
.Y(n_5020)
);

OAI21x1_ASAP7_75t_L g5021 ( 
.A1(n_4780),
.A2(n_4247),
.B(n_4240),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_SL g5022 ( 
.A(n_4726),
.B(n_4528),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4603),
.Y(n_5023)
);

OAI21xp5_ASAP7_75t_L g5024 ( 
.A1(n_4836),
.A2(n_4066),
.B(n_4533),
.Y(n_5024)
);

AOI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4580),
.A2(n_4525),
.B(n_4522),
.Y(n_5025)
);

AOI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_4763),
.A2(n_4525),
.B(n_4522),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4977),
.B(n_4419),
.Y(n_5027)
);

INVx2_ASAP7_75t_SL g5028 ( 
.A(n_4626),
.Y(n_5028)
);

BUFx6f_ASAP7_75t_L g5029 ( 
.A(n_4541),
.Y(n_5029)
);

AOI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_4546),
.A2(n_4525),
.B(n_4522),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4642),
.B(n_4355),
.Y(n_5031)
);

A2O1A1Ixp33_ASAP7_75t_L g5032 ( 
.A1(n_4890),
.A2(n_4509),
.B(n_4176),
.C(n_4220),
.Y(n_5032)
);

HB1xp67_ASAP7_75t_L g5033 ( 
.A(n_4895),
.Y(n_5033)
);

BUFx3_ASAP7_75t_L g5034 ( 
.A(n_4632),
.Y(n_5034)
);

AOI21xp5_ASAP7_75t_L g5035 ( 
.A1(n_4544),
.A2(n_4122),
.B(n_4110),
.Y(n_5035)
);

INVx4_ASAP7_75t_L g5036 ( 
.A(n_4905),
.Y(n_5036)
);

OAI22x1_ASAP7_75t_L g5037 ( 
.A1(n_4831),
.A2(n_4130),
.B1(n_4225),
.B2(n_4236),
.Y(n_5037)
);

OAI21xp5_ASAP7_75t_L g5038 ( 
.A1(n_4864),
.A2(n_4112),
.B(n_4302),
.Y(n_5038)
);

OAI21x1_ASAP7_75t_SL g5039 ( 
.A1(n_4640),
.A2(n_4390),
.B(n_4311),
.Y(n_5039)
);

INVx3_ASAP7_75t_L g5040 ( 
.A(n_4999),
.Y(n_5040)
);

OAI21x1_ASAP7_75t_L g5041 ( 
.A1(n_4911),
.A2(n_4554),
.B(n_4912),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4615),
.Y(n_5042)
);

NAND2x1_ASAP7_75t_L g5043 ( 
.A(n_4961),
.B(n_4146),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4870),
.B(n_4376),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4666),
.Y(n_5045)
);

AND2x2_ASAP7_75t_L g5046 ( 
.A(n_4693),
.B(n_4423),
.Y(n_5046)
);

AOI221x1_ASAP7_75t_L g5047 ( 
.A1(n_4938),
.A2(n_4224),
.B1(n_4528),
.B2(n_4358),
.C(n_4110),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_4772),
.B(n_4386),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4675),
.Y(n_5049)
);

OR2x2_ASAP7_75t_L g5050 ( 
.A(n_4567),
.B(n_4387),
.Y(n_5050)
);

AND2x4_ASAP7_75t_L g5051 ( 
.A(n_4557),
.B(n_4283),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4661),
.B(n_4391),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4582),
.B(n_4411),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4655),
.Y(n_5054)
);

A2O1A1Ixp33_ASAP7_75t_L g5055 ( 
.A1(n_4967),
.A2(n_4126),
.B(n_4145),
.C(n_4122),
.Y(n_5055)
);

OAI21x1_ASAP7_75t_L g5056 ( 
.A1(n_4566),
.A2(n_4268),
.B(n_4260),
.Y(n_5056)
);

INVxp67_ASAP7_75t_L g5057 ( 
.A(n_4635),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_L g5058 ( 
.A(n_4910),
.B(n_4293),
.Y(n_5058)
);

NAND2xp5_ASAP7_75t_SL g5059 ( 
.A(n_4830),
.B(n_3995),
.Y(n_5059)
);

AOI211x1_ASAP7_75t_L g5060 ( 
.A1(n_4872),
.A2(n_4182),
.B(n_4275),
.C(n_4270),
.Y(n_5060)
);

AND2x2_ASAP7_75t_L g5061 ( 
.A(n_4556),
.B(n_4293),
.Y(n_5061)
);

OAI21xp5_ASAP7_75t_L g5062 ( 
.A1(n_4901),
.A2(n_4048),
.B(n_4042),
.Y(n_5062)
);

INVx5_ASAP7_75t_L g5063 ( 
.A(n_4849),
.Y(n_5063)
);

OAI21x1_ASAP7_75t_L g5064 ( 
.A1(n_4536),
.A2(n_4068),
.B(n_4057),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4915),
.B(n_4042),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_4743),
.B(n_4048),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_4750),
.B(n_4099),
.Y(n_5067)
);

AND2x4_ASAP7_75t_L g5068 ( 
.A(n_4575),
.B(n_4126),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4691),
.Y(n_5069)
);

AOI21x1_ASAP7_75t_L g5070 ( 
.A1(n_4547),
.A2(n_4021),
.B(n_4145),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_4795),
.B(n_4099),
.Y(n_5071)
);

AOI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4989),
.A2(n_4519),
.B(n_4480),
.Y(n_5072)
);

INVx2_ASAP7_75t_L g5073 ( 
.A(n_4781),
.Y(n_5073)
);

OAI21x1_ASAP7_75t_L g5074 ( 
.A1(n_4601),
.A2(n_4072),
.B(n_4068),
.Y(n_5074)
);

AND2x4_ASAP7_75t_L g5075 ( 
.A(n_4577),
.B(n_4021),
.Y(n_5075)
);

NAND2xp33_ASAP7_75t_SL g5076 ( 
.A(n_4961),
.B(n_4068),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4841),
.B(n_4103),
.Y(n_5077)
);

NAND2x1p5_ASAP7_75t_L g5078 ( 
.A(n_4905),
.B(n_4072),
.Y(n_5078)
);

INVx2_ASAP7_75t_L g5079 ( 
.A(n_4620),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4857),
.B(n_4103),
.Y(n_5080)
);

NOR2xp67_ASAP7_75t_L g5081 ( 
.A(n_4905),
.B(n_396),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4676),
.B(n_4153),
.Y(n_5082)
);

INVx2_ASAP7_75t_L g5083 ( 
.A(n_4902),
.Y(n_5083)
);

INVx5_ASAP7_75t_L g5084 ( 
.A(n_4849),
.Y(n_5084)
);

AND2x4_ASAP7_75t_L g5085 ( 
.A(n_4594),
.B(n_4153),
.Y(n_5085)
);

OAI21x1_ASAP7_75t_L g5086 ( 
.A1(n_4601),
.A2(n_4076),
.B(n_4072),
.Y(n_5086)
);

NAND2x1p5_ASAP7_75t_L g5087 ( 
.A(n_4790),
.B(n_4076),
.Y(n_5087)
);

OAI21x1_ASAP7_75t_L g5088 ( 
.A1(n_4658),
.A2(n_4091),
.B(n_4076),
.Y(n_5088)
);

BUFx3_ASAP7_75t_L g5089 ( 
.A(n_4999),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4684),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_4730),
.B(n_4165),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4789),
.A2(n_4519),
.B(n_4480),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4698),
.Y(n_5093)
);

OA22x2_ASAP7_75t_L g5094 ( 
.A1(n_4613),
.A2(n_4177),
.B1(n_4194),
.B2(n_4165),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_4699),
.B(n_4177),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4801),
.A2(n_4519),
.B(n_4480),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_L g5097 ( 
.A(n_4850),
.B(n_4194),
.Y(n_5097)
);

OAI21x1_ASAP7_75t_L g5098 ( 
.A1(n_4658),
.A2(n_4140),
.B(n_4091),
.Y(n_5098)
);

INVx3_ASAP7_75t_L g5099 ( 
.A(n_4800),
.Y(n_5099)
);

AOI21xp5_ASAP7_75t_SL g5100 ( 
.A1(n_4709),
.A2(n_4140),
.B(n_4091),
.Y(n_5100)
);

OAI21x1_ASAP7_75t_L g5101 ( 
.A1(n_4725),
.A2(n_4169),
.B(n_4140),
.Y(n_5101)
);

NAND2xp5_ASAP7_75t_SL g5102 ( 
.A(n_4830),
.B(n_4169),
.Y(n_5102)
);

NAND2xp5_ASAP7_75t_SL g5103 ( 
.A(n_4891),
.B(n_4169),
.Y(n_5103)
);

OAI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4629),
.A2(n_4644),
.B(n_4589),
.Y(n_5104)
);

BUFx4f_ASAP7_75t_L g5105 ( 
.A(n_4887),
.Y(n_5105)
);

INVx2_ASAP7_75t_SL g5106 ( 
.A(n_4738),
.Y(n_5106)
);

OAI21x1_ASAP7_75t_L g5107 ( 
.A1(n_4725),
.A2(n_4548),
.B(n_4578),
.Y(n_5107)
);

AND2x4_ASAP7_75t_L g5108 ( 
.A(n_4651),
.B(n_4273),
.Y(n_5108)
);

OAI21x1_ASAP7_75t_L g5109 ( 
.A1(n_4892),
.A2(n_4304),
.B(n_4273),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_4899),
.B(n_397),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_SL g5111 ( 
.A(n_4837),
.B(n_4273),
.Y(n_5111)
);

INVx5_ASAP7_75t_L g5112 ( 
.A(n_4573),
.Y(n_5112)
);

BUFx4f_ASAP7_75t_L g5113 ( 
.A(n_4931),
.Y(n_5113)
);

AOI22xp5_ASAP7_75t_L g5114 ( 
.A1(n_4643),
.A2(n_4349),
.B1(n_4304),
.B2(n_400),
.Y(n_5114)
);

AOI21xp5_ASAP7_75t_SL g5115 ( 
.A1(n_4573),
.A2(n_4349),
.B(n_4304),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4818),
.A2(n_4349),
.B(n_398),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_4949),
.Y(n_5117)
);

AOI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_4828),
.A2(n_398),
.B(n_399),
.Y(n_5118)
);

OAI21x1_ASAP7_75t_L g5119 ( 
.A1(n_4563),
.A2(n_917),
.B(n_916),
.Y(n_5119)
);

INVx1_ASAP7_75t_SL g5120 ( 
.A(n_4591),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_4650),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_4951),
.Y(n_5122)
);

INVx3_ASAP7_75t_L g5123 ( 
.A(n_4541),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_4808),
.B(n_399),
.Y(n_5124)
);

OAI21x1_ASAP7_75t_L g5125 ( 
.A1(n_4569),
.A2(n_919),
.B(n_918),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_4883),
.B(n_399),
.Y(n_5126)
);

NOR2xp33_ASAP7_75t_L g5127 ( 
.A(n_4971),
.B(n_400),
.Y(n_5127)
);

AND2x2_ASAP7_75t_L g5128 ( 
.A(n_4543),
.B(n_400),
.Y(n_5128)
);

AND2x4_ASAP7_75t_L g5129 ( 
.A(n_4791),
.B(n_401),
.Y(n_5129)
);

OAI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4704),
.A2(n_919),
.B(n_918),
.Y(n_5130)
);

AND2x4_ASAP7_75t_L g5131 ( 
.A(n_4735),
.B(n_402),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4927),
.B(n_402),
.Y(n_5132)
);

AOI21xp5_ASAP7_75t_L g5133 ( 
.A1(n_4539),
.A2(n_402),
.B(n_403),
.Y(n_5133)
);

OAI21xp5_ASAP7_75t_L g5134 ( 
.A1(n_4809),
.A2(n_403),
.B(n_404),
.Y(n_5134)
);

OAI21x1_ASAP7_75t_L g5135 ( 
.A1(n_4913),
.A2(n_923),
.B(n_920),
.Y(n_5135)
);

AOI21xp5_ASAP7_75t_L g5136 ( 
.A1(n_4537),
.A2(n_404),
.B(n_405),
.Y(n_5136)
);

AND2x4_ASAP7_75t_L g5137 ( 
.A(n_4860),
.B(n_405),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4686),
.Y(n_5138)
);

OAI21x1_ASAP7_75t_SL g5139 ( 
.A1(n_4757),
.A2(n_413),
.B(n_405),
.Y(n_5139)
);

NOR2xp33_ASAP7_75t_SL g5140 ( 
.A(n_4597),
.B(n_406),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4706),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4980),
.B(n_406),
.Y(n_5142)
);

AOI221xp5_ASAP7_75t_L g5143 ( 
.A1(n_4764),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.C(n_409),
.Y(n_5143)
);

OR2x2_ASAP7_75t_L g5144 ( 
.A(n_4664),
.B(n_408),
.Y(n_5144)
);

AOI21x1_ASAP7_75t_SL g5145 ( 
.A1(n_4851),
.A2(n_409),
.B(n_410),
.Y(n_5145)
);

AND2x4_ASAP7_75t_L g5146 ( 
.A(n_4880),
.B(n_410),
.Y(n_5146)
);

OAI21x1_ASAP7_75t_L g5147 ( 
.A1(n_4551),
.A2(n_927),
.B(n_923),
.Y(n_5147)
);

AOI221xp5_ASAP7_75t_L g5148 ( 
.A1(n_4683),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.C(n_414),
.Y(n_5148)
);

INVx3_ASAP7_75t_L g5149 ( 
.A(n_4541),
.Y(n_5149)
);

OAI21x1_ASAP7_75t_L g5150 ( 
.A1(n_4886),
.A2(n_931),
.B(n_930),
.Y(n_5150)
);

OAI21x1_ASAP7_75t_L g5151 ( 
.A1(n_4886),
.A2(n_5006),
.B(n_4941),
.Y(n_5151)
);

BUFx2_ASAP7_75t_L g5152 ( 
.A(n_4866),
.Y(n_5152)
);

INVx4_ASAP7_75t_L g5153 ( 
.A(n_5000),
.Y(n_5153)
);

HB1xp67_ASAP7_75t_L g5154 ( 
.A(n_4602),
.Y(n_5154)
);

BUFx6f_ASAP7_75t_L g5155 ( 
.A(n_4820),
.Y(n_5155)
);

INVx3_ASAP7_75t_L g5156 ( 
.A(n_5000),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4981),
.B(n_411),
.Y(n_5157)
);

OAI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_5002),
.A2(n_411),
.B(n_412),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4552),
.Y(n_5159)
);

A2O1A1Ixp33_ASAP7_75t_L g5160 ( 
.A1(n_4700),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_5160)
);

NOR2x1_ASAP7_75t_SL g5161 ( 
.A(n_4922),
.B(n_415),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_4833),
.B(n_415),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4568),
.Y(n_5163)
);

AND2x2_ASAP7_75t_L g5164 ( 
.A(n_4571),
.B(n_415),
.Y(n_5164)
);

OAI21x1_ASAP7_75t_SL g5165 ( 
.A1(n_4997),
.A2(n_424),
.B(n_416),
.Y(n_5165)
);

AOI21x1_ASAP7_75t_L g5166 ( 
.A1(n_4874),
.A2(n_416),
.B(n_417),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_SL g5167 ( 
.A(n_4837),
.B(n_416),
.Y(n_5167)
);

AOI21x1_ASAP7_75t_L g5168 ( 
.A1(n_4627),
.A2(n_417),
.B(n_418),
.Y(n_5168)
);

A2O1A1Ixp33_ASAP7_75t_L g5169 ( 
.A1(n_4744),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_5169)
);

OAI21x1_ASAP7_75t_L g5170 ( 
.A1(n_4941),
.A2(n_933),
.B(n_932),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_4559),
.A2(n_419),
.B(n_420),
.Y(n_5171)
);

AOI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_4737),
.A2(n_420),
.B(n_421),
.Y(n_5172)
);

AND2x2_ASAP7_75t_L g5173 ( 
.A(n_4612),
.B(n_421),
.Y(n_5173)
);

AO21x2_ASAP7_75t_L g5174 ( 
.A1(n_4740),
.A2(n_421),
.B(n_422),
.Y(n_5174)
);

OAI21x1_ASAP7_75t_L g5175 ( 
.A1(n_5006),
.A2(n_934),
.B(n_933),
.Y(n_5175)
);

OAI21x1_ASAP7_75t_L g5176 ( 
.A1(n_4579),
.A2(n_936),
.B(n_935),
.Y(n_5176)
);

OAI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_4798),
.A2(n_422),
.B(n_423),
.Y(n_5177)
);

INVx1_ASAP7_75t_L g5178 ( 
.A(n_4921),
.Y(n_5178)
);

OAI21x1_ASAP7_75t_L g5179 ( 
.A1(n_4690),
.A2(n_937),
.B(n_936),
.Y(n_5179)
);

HB1xp67_ASAP7_75t_L g5180 ( 
.A(n_4680),
.Y(n_5180)
);

AO21x2_ASAP7_75t_L g5181 ( 
.A1(n_4746),
.A2(n_422),
.B(n_423),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_4727),
.B(n_423),
.Y(n_5182)
);

OAI21x1_ASAP7_75t_L g5183 ( 
.A1(n_4682),
.A2(n_939),
.B(n_938),
.Y(n_5183)
);

XNOR2xp5_ASAP7_75t_L g5184 ( 
.A(n_4983),
.B(n_424),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_4835),
.B(n_425),
.Y(n_5185)
);

AOI21xp5_ASAP7_75t_L g5186 ( 
.A1(n_4564),
.A2(n_425),
.B(n_426),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_4724),
.A2(n_425),
.B(n_426),
.Y(n_5187)
);

NOR2xp33_ASAP7_75t_L g5188 ( 
.A(n_4596),
.B(n_426),
.Y(n_5188)
);

INVx4_ASAP7_75t_L g5189 ( 
.A(n_4848),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_4731),
.B(n_427),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_4866),
.Y(n_5191)
);

OAI21x1_ASAP7_75t_L g5192 ( 
.A1(n_4768),
.A2(n_939),
.B(n_938),
.Y(n_5192)
);

OAI21x1_ASAP7_75t_L g5193 ( 
.A1(n_4773),
.A2(n_941),
.B(n_940),
.Y(n_5193)
);

AO31x2_ASAP7_75t_L g5194 ( 
.A1(n_4624),
.A2(n_4979),
.A3(n_4779),
.B(n_4871),
.Y(n_5194)
);

OAI22x1_ASAP7_75t_L g5195 ( 
.A1(n_4585),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_4751),
.B(n_427),
.Y(n_5196)
);

A2O1A1Ixp33_ASAP7_75t_L g5197 ( 
.A1(n_4560),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_5197)
);

AOI21x1_ASAP7_75t_L g5198 ( 
.A1(n_4679),
.A2(n_428),
.B(n_429),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_4572),
.B(n_430),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_4774),
.B(n_430),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4933),
.Y(n_5201)
);

OAI21x1_ASAP7_75t_L g5202 ( 
.A1(n_4711),
.A2(n_944),
.B(n_943),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_4815),
.B(n_431),
.Y(n_5203)
);

AOI211x1_ASAP7_75t_L g5204 ( 
.A1(n_4810),
.A2(n_433),
.B(n_431),
.C(n_432),
.Y(n_5204)
);

NAND2xp33_ASAP7_75t_SL g5205 ( 
.A(n_4786),
.B(n_431),
.Y(n_5205)
);

AO31x2_ASAP7_75t_L g5206 ( 
.A1(n_4754),
.A2(n_434),
.A3(n_432),
.B(n_433),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_L g5207 ( 
.A(n_4540),
.B(n_433),
.Y(n_5207)
);

AOI21xp5_ASAP7_75t_L g5208 ( 
.A1(n_4595),
.A2(n_434),
.B(n_435),
.Y(n_5208)
);

NAND2x1p5_ASAP7_75t_L g5209 ( 
.A(n_4906),
.B(n_435),
.Y(n_5209)
);

NOR2xp33_ASAP7_75t_SL g5210 ( 
.A(n_4712),
.B(n_435),
.Y(n_5210)
);

HB1xp67_ASAP7_75t_L g5211 ( 
.A(n_4985),
.Y(n_5211)
);

OAI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4944),
.A2(n_4702),
.B(n_4673),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_4558),
.B(n_436),
.Y(n_5213)
);

AND2x2_ASAP7_75t_L g5214 ( 
.A(n_4732),
.B(n_4819),
.Y(n_5214)
);

CKINVDCx20_ASAP7_75t_R g5215 ( 
.A(n_4766),
.Y(n_5215)
);

OAI21x1_ASAP7_75t_L g5216 ( 
.A1(n_4600),
.A2(n_4604),
.B(n_4671),
.Y(n_5216)
);

O2A1O1Ixp5_ASAP7_75t_L g5217 ( 
.A1(n_4867),
.A2(n_438),
.B(n_436),
.C(n_437),
.Y(n_5217)
);

INVx3_ASAP7_75t_L g5218 ( 
.A(n_4802),
.Y(n_5218)
);

OAI21x1_ASAP7_75t_L g5219 ( 
.A1(n_4678),
.A2(n_944),
.B(n_943),
.Y(n_5219)
);

OAI21x1_ASAP7_75t_L g5220 ( 
.A1(n_4654),
.A2(n_948),
.B(n_946),
.Y(n_5220)
);

BUFx2_ASAP7_75t_L g5221 ( 
.A(n_4866),
.Y(n_5221)
);

OAI21x1_ASAP7_75t_L g5222 ( 
.A1(n_4765),
.A2(n_948),
.B(n_946),
.Y(n_5222)
);

AND2x4_ASAP7_75t_L g5223 ( 
.A(n_4960),
.B(n_436),
.Y(n_5223)
);

AOI21xp33_ASAP7_75t_L g5224 ( 
.A1(n_4846),
.A2(n_437),
.B(n_438),
.Y(n_5224)
);

AOI21xp5_ASAP7_75t_L g5225 ( 
.A1(n_4593),
.A2(n_438),
.B(n_439),
.Y(n_5225)
);

AOI21xp5_ASAP7_75t_L g5226 ( 
.A1(n_4630),
.A2(n_439),
.B(n_440),
.Y(n_5226)
);

BUFx2_ASAP7_75t_L g5227 ( 
.A(n_4976),
.Y(n_5227)
);

AOI21xp5_ASAP7_75t_L g5228 ( 
.A1(n_4637),
.A2(n_439),
.B(n_440),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_4854),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4584),
.Y(n_5230)
);

INVx4_ASAP7_75t_L g5231 ( 
.A(n_4804),
.Y(n_5231)
);

NOR2x1p5_ASAP7_75t_L g5232 ( 
.A(n_4997),
.B(n_440),
.Y(n_5232)
);

BUFx6f_ASAP7_75t_L g5233 ( 
.A(n_4663),
.Y(n_5233)
);

AOI21xp5_ASAP7_75t_L g5234 ( 
.A1(n_4641),
.A2(n_441),
.B(n_442),
.Y(n_5234)
);

NAND2x1_ASAP7_75t_L g5235 ( 
.A(n_4741),
.B(n_442),
.Y(n_5235)
);

NAND2xp5_ASAP7_75t_L g5236 ( 
.A(n_4545),
.B(n_443),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_4587),
.Y(n_5237)
);

AOI21xp5_ASAP7_75t_L g5238 ( 
.A1(n_4770),
.A2(n_443),
.B(n_444),
.Y(n_5238)
);

AO31x2_ASAP7_75t_L g5239 ( 
.A1(n_4753),
.A2(n_445),
.A3(n_443),
.B(n_444),
.Y(n_5239)
);

INVx3_ASAP7_75t_L g5240 ( 
.A(n_4858),
.Y(n_5240)
);

BUFx4_ASAP7_75t_SL g5241 ( 
.A(n_4956),
.Y(n_5241)
);

OAI21x1_ASAP7_75t_L g5242 ( 
.A1(n_4767),
.A2(n_950),
.B(n_949),
.Y(n_5242)
);

A2O1A1Ixp33_ASAP7_75t_L g5243 ( 
.A1(n_4717),
.A2(n_446),
.B(n_444),
.C(n_445),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_4599),
.B(n_445),
.Y(n_5244)
);

AND2x2_ASAP7_75t_SL g5245 ( 
.A(n_4906),
.B(n_4663),
.Y(n_5245)
);

BUFx2_ASAP7_75t_L g5246 ( 
.A(n_4976),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_4606),
.Y(n_5247)
);

OAI21x1_ASAP7_75t_L g5248 ( 
.A1(n_4605),
.A2(n_950),
.B(n_949),
.Y(n_5248)
);

OAI21x1_ASAP7_75t_L g5249 ( 
.A1(n_4681),
.A2(n_952),
.B(n_951),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4553),
.B(n_4562),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_4610),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_4617),
.B(n_446),
.Y(n_5252)
);

AOI21x1_ASAP7_75t_SL g5253 ( 
.A1(n_4868),
.A2(n_446),
.B(n_447),
.Y(n_5253)
);

NOR2x1_ASAP7_75t_L g5254 ( 
.A(n_4701),
.B(n_447),
.Y(n_5254)
);

OAI21xp5_ASAP7_75t_L g5255 ( 
.A1(n_4865),
.A2(n_448),
.B(n_449),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_4618),
.B(n_448),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_4619),
.B(n_448),
.Y(n_5257)
);

OAI21x1_ASAP7_75t_L g5258 ( 
.A1(n_4685),
.A2(n_4692),
.B(n_4687),
.Y(n_5258)
);

OAI21x1_ASAP7_75t_L g5259 ( 
.A1(n_4623),
.A2(n_952),
.B(n_951),
.Y(n_5259)
);

BUFx3_ASAP7_75t_L g5260 ( 
.A(n_4733),
.Y(n_5260)
);

OAI21x1_ASAP7_75t_L g5261 ( 
.A1(n_4625),
.A2(n_955),
.B(n_953),
.Y(n_5261)
);

AND2x2_ASAP7_75t_L g5262 ( 
.A(n_4550),
.B(n_449),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4634),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_4645),
.B(n_449),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_4646),
.B(n_450),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_4649),
.Y(n_5266)
);

OAI21x1_ASAP7_75t_L g5267 ( 
.A1(n_4639),
.A2(n_956),
.B(n_953),
.Y(n_5267)
);

AO31x2_ASAP7_75t_L g5268 ( 
.A1(n_4638),
.A2(n_4748),
.A3(n_4884),
.B(n_4842),
.Y(n_5268)
);

OAI21x1_ASAP7_75t_L g5269 ( 
.A1(n_4648),
.A2(n_957),
.B(n_956),
.Y(n_5269)
);

OAI21x1_ASAP7_75t_L g5270 ( 
.A1(n_4653),
.A2(n_958),
.B(n_957),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_4976),
.Y(n_5271)
);

AND3x4_ASAP7_75t_L g5272 ( 
.A(n_4950),
.B(n_450),
.C(n_451),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_L g5273 ( 
.A(n_4660),
.B(n_451),
.Y(n_5273)
);

NAND2xp33_ASAP7_75t_L g5274 ( 
.A(n_4837),
.B(n_452),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_4667),
.B(n_452),
.Y(n_5275)
);

AOI21x1_ASAP7_75t_L g5276 ( 
.A1(n_4749),
.A2(n_453),
.B(n_454),
.Y(n_5276)
);

AOI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_4719),
.A2(n_453),
.B(n_454),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4669),
.Y(n_5278)
);

OAI21x1_ASAP7_75t_L g5279 ( 
.A1(n_4974),
.A2(n_960),
.B(n_959),
.Y(n_5279)
);

AND2x2_ASAP7_75t_L g5280 ( 
.A(n_4688),
.B(n_453),
.Y(n_5280)
);

OAI21x1_ASAP7_75t_L g5281 ( 
.A1(n_4723),
.A2(n_960),
.B(n_959),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4672),
.Y(n_5282)
);

AOI21x1_ASAP7_75t_L g5283 ( 
.A1(n_4622),
.A2(n_454),
.B(n_455),
.Y(n_5283)
);

NAND2xp5_ASAP7_75t_SL g5284 ( 
.A(n_4837),
.B(n_455),
.Y(n_5284)
);

OA22x2_ASAP7_75t_L g5285 ( 
.A1(n_4656),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_5285)
);

AND2x4_ASAP7_75t_L g5286 ( 
.A(n_4799),
.B(n_456),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_4694),
.B(n_456),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4538),
.A2(n_457),
.B(n_458),
.Y(n_5288)
);

NAND3xp33_ASAP7_75t_L g5289 ( 
.A(n_4697),
.B(n_457),
.C(n_458),
.Y(n_5289)
);

INVx2_ASAP7_75t_SL g5290 ( 
.A(n_4837),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_4588),
.B(n_459),
.Y(n_5291)
);

NOR2x1_ASAP7_75t_L g5292 ( 
.A(n_4628),
.B(n_459),
.Y(n_5292)
);

INVx2_ASAP7_75t_L g5293 ( 
.A(n_4969),
.Y(n_5293)
);

OAI21x1_ASAP7_75t_L g5294 ( 
.A1(n_4714),
.A2(n_963),
.B(n_961),
.Y(n_5294)
);

AOI21xp5_ASAP7_75t_L g5295 ( 
.A1(n_4984),
.A2(n_459),
.B(n_460),
.Y(n_5295)
);

AND2x2_ASAP7_75t_L g5296 ( 
.A(n_4926),
.B(n_460),
.Y(n_5296)
);

AND2x4_ASAP7_75t_L g5297 ( 
.A(n_4607),
.B(n_4663),
.Y(n_5297)
);

OAI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_4904),
.A2(n_460),
.B(n_461),
.Y(n_5298)
);

OAI21x1_ASAP7_75t_L g5299 ( 
.A1(n_4882),
.A2(n_964),
.B(n_963),
.Y(n_5299)
);

OAI21x1_ASAP7_75t_L g5300 ( 
.A1(n_4668),
.A2(n_965),
.B(n_964),
.Y(n_5300)
);

BUFx3_ASAP7_75t_L g5301 ( 
.A(n_4973),
.Y(n_5301)
);

OAI21xp5_ASAP7_75t_L g5302 ( 
.A1(n_4943),
.A2(n_461),
.B(n_462),
.Y(n_5302)
);

AO31x2_ASAP7_75t_L g5303 ( 
.A1(n_4962),
.A2(n_463),
.A3(n_461),
.B(n_462),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_4708),
.B(n_463),
.Y(n_5304)
);

BUFx3_ASAP7_75t_L g5305 ( 
.A(n_4647),
.Y(n_5305)
);

AOI21x1_ASAP7_75t_L g5306 ( 
.A1(n_4955),
.A2(n_464),
.B(n_465),
.Y(n_5306)
);

AOI21xp5_ASAP7_75t_SL g5307 ( 
.A1(n_5008),
.A2(n_464),
.B(n_465),
.Y(n_5307)
);

OAI22xp5_ASAP7_75t_L g5308 ( 
.A1(n_4657),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_5308)
);

BUFx2_ASAP7_75t_L g5309 ( 
.A(n_4741),
.Y(n_5309)
);

INVx4_ASAP7_75t_L g5310 ( 
.A(n_4741),
.Y(n_5310)
);

INVx3_ASAP7_75t_L g5311 ( 
.A(n_4741),
.Y(n_5311)
);

A2O1A1Ixp33_ASAP7_75t_L g5312 ( 
.A1(n_4722),
.A2(n_469),
.B(n_467),
.C(n_468),
.Y(n_5312)
);

OAI21x1_ASAP7_75t_L g5313 ( 
.A1(n_4881),
.A2(n_966),
.B(n_965),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_4710),
.Y(n_5314)
);

AO21x1_ASAP7_75t_L g5315 ( 
.A1(n_4583),
.A2(n_467),
.B(n_468),
.Y(n_5315)
);

AOI221x1_ASAP7_75t_L g5316 ( 
.A1(n_4916),
.A2(n_968),
.B1(n_969),
.B2(n_967),
.C(n_966),
.Y(n_5316)
);

OAI21xp5_ASAP7_75t_L g5317 ( 
.A1(n_4988),
.A2(n_469),
.B(n_470),
.Y(n_5317)
);

NAND2x1_ASAP7_75t_L g5318 ( 
.A(n_4555),
.B(n_470),
.Y(n_5318)
);

NAND2xp5_ASAP7_75t_SL g5319 ( 
.A(n_4570),
.B(n_471),
.Y(n_5319)
);

OAI21x1_ASAP7_75t_L g5320 ( 
.A1(n_4608),
.A2(n_969),
.B(n_967),
.Y(n_5320)
);

OAI21xp5_ASAP7_75t_L g5321 ( 
.A1(n_4928),
.A2(n_471),
.B(n_472),
.Y(n_5321)
);

NAND2xp5_ASAP7_75t_SL g5322 ( 
.A(n_4696),
.B(n_4863),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_4716),
.B(n_471),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_4821),
.B(n_472),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_5033),
.B(n_4787),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5121),
.B(n_4720),
.Y(n_5326)
);

BUFx3_ASAP7_75t_L g5327 ( 
.A(n_5034),
.Y(n_5327)
);

INVx2_ASAP7_75t_SL g5328 ( 
.A(n_5089),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_5015),
.Y(n_5329)
);

HB1xp67_ASAP7_75t_L g5330 ( 
.A(n_5154),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5023),
.Y(n_5331)
);

INVx2_ASAP7_75t_L g5332 ( 
.A(n_5050),
.Y(n_5332)
);

CKINVDCx5p33_ASAP7_75t_R g5333 ( 
.A(n_5241),
.Y(n_5333)
);

INVx3_ASAP7_75t_SL g5334 ( 
.A(n_5189),
.Y(n_5334)
);

BUFx2_ASAP7_75t_L g5335 ( 
.A(n_5051),
.Y(n_5335)
);

INVxp67_ASAP7_75t_SL g5336 ( 
.A(n_5211),
.Y(n_5336)
);

OR2x6_ASAP7_75t_L g5337 ( 
.A(n_5028),
.B(n_4736),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_L g5338 ( 
.A(n_5138),
.B(n_4739),
.Y(n_5338)
);

INVx5_ASAP7_75t_L g5339 ( 
.A(n_5231),
.Y(n_5339)
);

OR2x2_ASAP7_75t_L g5340 ( 
.A(n_5180),
.B(n_5031),
.Y(n_5340)
);

BUFx6f_ASAP7_75t_SL g5341 ( 
.A(n_5106),
.Y(n_5341)
);

INVx2_ASAP7_75t_L g5342 ( 
.A(n_5054),
.Y(n_5342)
);

BUFx3_ASAP7_75t_L g5343 ( 
.A(n_5099),
.Y(n_5343)
);

BUFx3_ASAP7_75t_L g5344 ( 
.A(n_5040),
.Y(n_5344)
);

INVx5_ASAP7_75t_L g5345 ( 
.A(n_5063),
.Y(n_5345)
);

AOI22xp33_ASAP7_75t_SL g5346 ( 
.A1(n_5309),
.A2(n_4555),
.B1(n_4932),
.B2(n_4659),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5042),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_5141),
.B(n_4822),
.Y(n_5348)
);

INVx3_ASAP7_75t_SL g5349 ( 
.A(n_5215),
.Y(n_5349)
);

BUFx12f_ASAP7_75t_L g5350 ( 
.A(n_5153),
.Y(n_5350)
);

BUFx12f_ASAP7_75t_L g5351 ( 
.A(n_5155),
.Y(n_5351)
);

BUFx3_ASAP7_75t_L g5352 ( 
.A(n_5113),
.Y(n_5352)
);

INVx8_ASAP7_75t_L g5353 ( 
.A(n_5155),
.Y(n_5353)
);

AND2x2_ASAP7_75t_L g5354 ( 
.A(n_5020),
.B(n_4665),
.Y(n_5354)
);

INVx3_ASAP7_75t_L g5355 ( 
.A(n_5105),
.Y(n_5355)
);

INVx1_ASAP7_75t_SL g5356 ( 
.A(n_5120),
.Y(n_5356)
);

INVx2_ASAP7_75t_L g5357 ( 
.A(n_5069),
.Y(n_5357)
);

INVx5_ASAP7_75t_L g5358 ( 
.A(n_5063),
.Y(n_5358)
);

INVx2_ASAP7_75t_L g5359 ( 
.A(n_5073),
.Y(n_5359)
);

INVx2_ASAP7_75t_L g5360 ( 
.A(n_5079),
.Y(n_5360)
);

INVx1_ASAP7_75t_SL g5361 ( 
.A(n_5260),
.Y(n_5361)
);

AND2x4_ASAP7_75t_L g5362 ( 
.A(n_5112),
.B(n_4555),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5045),
.Y(n_5363)
);

INVx5_ASAP7_75t_L g5364 ( 
.A(n_5063),
.Y(n_5364)
);

BUFx6f_ASAP7_75t_L g5365 ( 
.A(n_5233),
.Y(n_5365)
);

AND2x4_ASAP7_75t_L g5366 ( 
.A(n_5112),
.B(n_4555),
.Y(n_5366)
);

BUFx2_ASAP7_75t_L g5367 ( 
.A(n_5112),
.Y(n_5367)
);

CKINVDCx5p33_ASAP7_75t_R g5368 ( 
.A(n_5156),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_5178),
.B(n_4598),
.Y(n_5369)
);

INVx5_ASAP7_75t_SL g5370 ( 
.A(n_5131),
.Y(n_5370)
);

INVx3_ASAP7_75t_L g5371 ( 
.A(n_5014),
.Y(n_5371)
);

INVxp67_ASAP7_75t_SL g5372 ( 
.A(n_5057),
.Y(n_5372)
);

INVx5_ASAP7_75t_SL g5373 ( 
.A(n_5146),
.Y(n_5373)
);

INVx5_ASAP7_75t_L g5374 ( 
.A(n_5084),
.Y(n_5374)
);

AOI22xp33_ASAP7_75t_L g5375 ( 
.A1(n_5309),
.A2(n_4707),
.B1(n_4972),
.B2(n_4689),
.Y(n_5375)
);

BUFx8_ASAP7_75t_L g5376 ( 
.A(n_5297),
.Y(n_5376)
);

BUFx6f_ASAP7_75t_L g5377 ( 
.A(n_5233),
.Y(n_5377)
);

INVx2_ASAP7_75t_L g5378 ( 
.A(n_5083),
.Y(n_5378)
);

NAND2x1p5_ASAP7_75t_L g5379 ( 
.A(n_5084),
.B(n_4888),
.Y(n_5379)
);

BUFx12f_ASAP7_75t_L g5380 ( 
.A(n_5223),
.Y(n_5380)
);

BUFx12f_ASAP7_75t_L g5381 ( 
.A(n_5137),
.Y(n_5381)
);

INVx5_ASAP7_75t_L g5382 ( 
.A(n_5084),
.Y(n_5382)
);

BUFx12f_ASAP7_75t_L g5383 ( 
.A(n_5209),
.Y(n_5383)
);

BUFx6f_ASAP7_75t_L g5384 ( 
.A(n_5029),
.Y(n_5384)
);

BUFx4f_ASAP7_75t_SL g5385 ( 
.A(n_5240),
.Y(n_5385)
);

BUFx6f_ASAP7_75t_L g5386 ( 
.A(n_5029),
.Y(n_5386)
);

BUFx3_ASAP7_75t_L g5387 ( 
.A(n_5046),
.Y(n_5387)
);

INVx2_ASAP7_75t_L g5388 ( 
.A(n_5117),
.Y(n_5388)
);

INVxp67_ASAP7_75t_SL g5389 ( 
.A(n_5122),
.Y(n_5389)
);

HB1xp67_ASAP7_75t_L g5390 ( 
.A(n_5048),
.Y(n_5390)
);

BUFx12f_ASAP7_75t_L g5391 ( 
.A(n_5232),
.Y(n_5391)
);

INVx1_ASAP7_75t_SL g5392 ( 
.A(n_5085),
.Y(n_5392)
);

BUFx3_ASAP7_75t_L g5393 ( 
.A(n_5218),
.Y(n_5393)
);

INVx5_ASAP7_75t_L g5394 ( 
.A(n_5036),
.Y(n_5394)
);

BUFx3_ASAP7_75t_L g5395 ( 
.A(n_5075),
.Y(n_5395)
);

INVx3_ASAP7_75t_L g5396 ( 
.A(n_5043),
.Y(n_5396)
);

INVxp67_ASAP7_75t_SL g5397 ( 
.A(n_5018),
.Y(n_5397)
);

BUFx3_ASAP7_75t_L g5398 ( 
.A(n_5068),
.Y(n_5398)
);

BUFx2_ASAP7_75t_SL g5399 ( 
.A(n_5081),
.Y(n_5399)
);

BUFx6f_ASAP7_75t_L g5400 ( 
.A(n_5108),
.Y(n_5400)
);

INVx2_ASAP7_75t_L g5401 ( 
.A(n_5049),
.Y(n_5401)
);

NOR2xp33_ASAP7_75t_L g5402 ( 
.A(n_5305),
.B(n_4542),
.Y(n_5402)
);

INVx2_ASAP7_75t_L g5403 ( 
.A(n_5090),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5093),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_5012),
.Y(n_5405)
);

INVx5_ASAP7_75t_L g5406 ( 
.A(n_5123),
.Y(n_5406)
);

BUFx6f_ASAP7_75t_L g5407 ( 
.A(n_5149),
.Y(n_5407)
);

INVx3_ASAP7_75t_SL g5408 ( 
.A(n_5245),
.Y(n_5408)
);

CKINVDCx11_ASAP7_75t_R g5409 ( 
.A(n_5301),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_5159),
.Y(n_5410)
);

INVx4_ASAP7_75t_L g5411 ( 
.A(n_5272),
.Y(n_5411)
);

INVx2_ASAP7_75t_L g5412 ( 
.A(n_5163),
.Y(n_5412)
);

BUFx12f_ASAP7_75t_L g5413 ( 
.A(n_5129),
.Y(n_5413)
);

INVx2_ASAP7_75t_L g5414 ( 
.A(n_5066),
.Y(n_5414)
);

INVxp67_ASAP7_75t_SL g5415 ( 
.A(n_5053),
.Y(n_5415)
);

BUFx12f_ASAP7_75t_L g5416 ( 
.A(n_5286),
.Y(n_5416)
);

INVx1_ASAP7_75t_SL g5417 ( 
.A(n_5091),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5044),
.Y(n_5418)
);

INVxp67_ASAP7_75t_SL g5419 ( 
.A(n_5097),
.Y(n_5419)
);

NOR2xp33_ASAP7_75t_L g5420 ( 
.A(n_5127),
.B(n_5188),
.Y(n_5420)
);

BUFx2_ASAP7_75t_L g5421 ( 
.A(n_5076),
.Y(n_5421)
);

BUFx6f_ASAP7_75t_L g5422 ( 
.A(n_5087),
.Y(n_5422)
);

BUFx6f_ASAP7_75t_L g5423 ( 
.A(n_5152),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5201),
.Y(n_5424)
);

BUFx3_ASAP7_75t_L g5425 ( 
.A(n_5027),
.Y(n_5425)
);

BUFx2_ASAP7_75t_L g5426 ( 
.A(n_5152),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5067),
.Y(n_5427)
);

CKINVDCx20_ASAP7_75t_R g5428 ( 
.A(n_5205),
.Y(n_5428)
);

NAND2xp5_ASAP7_75t_L g5429 ( 
.A(n_5230),
.B(n_4936),
.Y(n_5429)
);

INVx1_ASAP7_75t_SL g5430 ( 
.A(n_5052),
.Y(n_5430)
);

BUFx2_ASAP7_75t_L g5431 ( 
.A(n_5221),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_5237),
.B(n_4832),
.Y(n_5432)
);

BUFx8_ASAP7_75t_L g5433 ( 
.A(n_5173),
.Y(n_5433)
);

BUFx6f_ASAP7_75t_L g5434 ( 
.A(n_5221),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5071),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_5077),
.Y(n_5436)
);

BUFx12f_ASAP7_75t_L g5437 ( 
.A(n_5011),
.Y(n_5437)
);

INVx3_ASAP7_75t_L g5438 ( 
.A(n_5310),
.Y(n_5438)
);

INVx4_ASAP7_75t_L g5439 ( 
.A(n_5078),
.Y(n_5439)
);

BUFx2_ASAP7_75t_SL g5440 ( 
.A(n_5103),
.Y(n_5440)
);

AOI22xp33_ASAP7_75t_L g5441 ( 
.A1(n_5094),
.A2(n_4877),
.B1(n_4843),
.B2(n_4807),
.Y(n_5441)
);

INVx2_ASAP7_75t_SL g5442 ( 
.A(n_5061),
.Y(n_5442)
);

BUFx3_ASAP7_75t_L g5443 ( 
.A(n_5227),
.Y(n_5443)
);

BUFx8_ASAP7_75t_L g5444 ( 
.A(n_5262),
.Y(n_5444)
);

BUFx3_ASAP7_75t_L g5445 ( 
.A(n_5227),
.Y(n_5445)
);

INVx1_ASAP7_75t_L g5446 ( 
.A(n_5080),
.Y(n_5446)
);

BUFx12f_ASAP7_75t_L g5447 ( 
.A(n_5185),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_L g5448 ( 
.A(n_5247),
.B(n_4745),
.Y(n_5448)
);

AND2x6_ASAP7_75t_L g5449 ( 
.A(n_5311),
.B(n_4896),
.Y(n_5449)
);

BUFx6f_ASAP7_75t_L g5450 ( 
.A(n_5246),
.Y(n_5450)
);

INVx4_ASAP7_75t_L g5451 ( 
.A(n_5246),
.Y(n_5451)
);

BUFx4f_ASAP7_75t_SL g5452 ( 
.A(n_5059),
.Y(n_5452)
);

NOR2xp33_ASAP7_75t_L g5453 ( 
.A(n_5210),
.B(n_4806),
.Y(n_5453)
);

INVx5_ASAP7_75t_L g5454 ( 
.A(n_5290),
.Y(n_5454)
);

BUFx2_ASAP7_75t_L g5455 ( 
.A(n_5151),
.Y(n_5455)
);

BUFx3_ASAP7_75t_L g5456 ( 
.A(n_5214),
.Y(n_5456)
);

BUFx3_ASAP7_75t_L g5457 ( 
.A(n_5199),
.Y(n_5457)
);

BUFx6f_ASAP7_75t_L g5458 ( 
.A(n_5191),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5058),
.Y(n_5459)
);

BUFx6f_ASAP7_75t_L g5460 ( 
.A(n_5271),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5065),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_5082),
.Y(n_5462)
);

BUFx6f_ASAP7_75t_L g5463 ( 
.A(n_5074),
.Y(n_5463)
);

INVx1_ASAP7_75t_SL g5464 ( 
.A(n_5037),
.Y(n_5464)
);

AND2x4_ASAP7_75t_L g5465 ( 
.A(n_5161),
.B(n_5095),
.Y(n_5465)
);

INVx2_ASAP7_75t_L g5466 ( 
.A(n_5293),
.Y(n_5466)
);

BUFx4f_ASAP7_75t_SL g5467 ( 
.A(n_5022),
.Y(n_5467)
);

INVx4_ASAP7_75t_L g5468 ( 
.A(n_5285),
.Y(n_5468)
);

INVx1_ASAP7_75t_SL g5469 ( 
.A(n_5144),
.Y(n_5469)
);

INVx2_ASAP7_75t_SL g5470 ( 
.A(n_5128),
.Y(n_5470)
);

INVx3_ASAP7_75t_L g5471 ( 
.A(n_5235),
.Y(n_5471)
);

AND2x2_ASAP7_75t_L g5472 ( 
.A(n_5229),
.B(n_4925),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_5251),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5263),
.Y(n_5474)
);

AOI22xp33_ASAP7_75t_L g5475 ( 
.A1(n_5322),
.A2(n_4817),
.B1(n_4838),
.B2(n_4824),
.Y(n_5475)
);

BUFx12f_ASAP7_75t_L g5476 ( 
.A(n_5280),
.Y(n_5476)
);

NAND2xp5_ASAP7_75t_L g5477 ( 
.A(n_5266),
.B(n_4752),
.Y(n_5477)
);

INVx3_ASAP7_75t_L g5478 ( 
.A(n_5318),
.Y(n_5478)
);

INVx2_ASAP7_75t_SL g5479 ( 
.A(n_5164),
.Y(n_5479)
);

BUFx3_ASAP7_75t_L g5480 ( 
.A(n_5086),
.Y(n_5480)
);

BUFx2_ASAP7_75t_L g5481 ( 
.A(n_5088),
.Y(n_5481)
);

BUFx2_ASAP7_75t_L g5482 ( 
.A(n_5098),
.Y(n_5482)
);

INVx4_ASAP7_75t_L g5483 ( 
.A(n_5174),
.Y(n_5483)
);

INVx3_ASAP7_75t_L g5484 ( 
.A(n_5101),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5278),
.Y(n_5485)
);

INVx5_ASAP7_75t_L g5486 ( 
.A(n_5244),
.Y(n_5486)
);

BUFx8_ASAP7_75t_SL g5487 ( 
.A(n_5190),
.Y(n_5487)
);

BUFx2_ASAP7_75t_SL g5488 ( 
.A(n_5102),
.Y(n_5488)
);

OAI22xp33_ASAP7_75t_L g5489 ( 
.A1(n_5140),
.A2(n_4776),
.B1(n_4939),
.B2(n_4839),
.Y(n_5489)
);

INVx3_ASAP7_75t_L g5490 ( 
.A(n_5283),
.Y(n_5490)
);

INVx6_ASAP7_75t_L g5491 ( 
.A(n_5291),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_SL g5492 ( 
.A(n_5039),
.B(n_4576),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5109),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_5070),
.Y(n_5494)
);

NAND2x1p5_ASAP7_75t_L g5495 ( 
.A(n_5254),
.B(n_4930),
.Y(n_5495)
);

BUFx6f_ASAP7_75t_L g5496 ( 
.A(n_5150),
.Y(n_5496)
);

INVx3_ASAP7_75t_L g5497 ( 
.A(n_5070),
.Y(n_5497)
);

INVx2_ASAP7_75t_L g5498 ( 
.A(n_5019),
.Y(n_5498)
);

NAND2x1p5_ASAP7_75t_L g5499 ( 
.A(n_5292),
.B(n_4954),
.Y(n_5499)
);

BUFx5_ASAP7_75t_L g5500 ( 
.A(n_5282),
.Y(n_5500)
);

BUFx6f_ASAP7_75t_L g5501 ( 
.A(n_5170),
.Y(n_5501)
);

NAND2x1p5_ASAP7_75t_L g5502 ( 
.A(n_5319),
.B(n_4964),
.Y(n_5502)
);

INVx2_ASAP7_75t_L g5503 ( 
.A(n_5019),
.Y(n_5503)
);

NOR2xp33_ASAP7_75t_SL g5504 ( 
.A(n_5032),
.B(n_4879),
.Y(n_5504)
);

NAND2x1p5_ASAP7_75t_L g5505 ( 
.A(n_5175),
.B(n_4893),
.Y(n_5505)
);

INVx1_ASAP7_75t_L g5506 ( 
.A(n_5314),
.Y(n_5506)
);

BUFx6f_ASAP7_75t_L g5507 ( 
.A(n_5111),
.Y(n_5507)
);

OAI22xp33_ASAP7_75t_SL g5508 ( 
.A1(n_5167),
.A2(n_5001),
.B1(n_4991),
.B2(n_4957),
.Y(n_5508)
);

AND2x2_ASAP7_75t_L g5509 ( 
.A(n_5250),
.B(n_5296),
.Y(n_5509)
);

CKINVDCx20_ASAP7_75t_R g5510 ( 
.A(n_5184),
.Y(n_5510)
);

INVx5_ASAP7_75t_L g5511 ( 
.A(n_5324),
.Y(n_5511)
);

OR2x6_ASAP7_75t_L g5512 ( 
.A(n_5391),
.B(n_5100),
.Y(n_5512)
);

BUFx4f_ASAP7_75t_L g5513 ( 
.A(n_5334),
.Y(n_5513)
);

INVx3_ASAP7_75t_L g5514 ( 
.A(n_5344),
.Y(n_5514)
);

AO31x2_ASAP7_75t_L g5515 ( 
.A1(n_5455),
.A2(n_5047),
.A3(n_5072),
.B(n_5195),
.Y(n_5515)
);

BUFx2_ASAP7_75t_L g5516 ( 
.A(n_5451),
.Y(n_5516)
);

OA21x2_ASAP7_75t_L g5517 ( 
.A1(n_5481),
.A2(n_5041),
.B(n_5064),
.Y(n_5517)
);

HB1xp67_ASAP7_75t_L g5518 ( 
.A(n_5330),
.Y(n_5518)
);

AND2x4_ASAP7_75t_L g5519 ( 
.A(n_5387),
.B(n_5055),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_L g5520 ( 
.A1(n_5468),
.A2(n_5104),
.B1(n_5315),
.B2(n_5212),
.Y(n_5520)
);

INVx3_ASAP7_75t_L g5521 ( 
.A(n_5376),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5329),
.Y(n_5522)
);

OAI21x1_ASAP7_75t_L g5523 ( 
.A1(n_5484),
.A2(n_5039),
.B(n_5025),
.Y(n_5523)
);

OAI22xp5_ASAP7_75t_L g5524 ( 
.A1(n_5346),
.A2(n_5184),
.B1(n_5060),
.B2(n_5035),
.Y(n_5524)
);

INVx1_ASAP7_75t_SL g5525 ( 
.A(n_5409),
.Y(n_5525)
);

OAI22xp5_ASAP7_75t_L g5526 ( 
.A1(n_5428),
.A2(n_5289),
.B1(n_5172),
.B2(n_5204),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_5500),
.Y(n_5527)
);

INVx2_ASAP7_75t_L g5528 ( 
.A(n_5500),
.Y(n_5528)
);

BUFx3_ASAP7_75t_L g5529 ( 
.A(n_5351),
.Y(n_5529)
);

AOI21xp5_ASAP7_75t_SL g5530 ( 
.A1(n_5421),
.A2(n_5197),
.B(n_5160),
.Y(n_5530)
);

AO21x2_ASAP7_75t_L g5531 ( 
.A1(n_5494),
.A2(n_5165),
.B(n_5026),
.Y(n_5531)
);

OAI21x1_ASAP7_75t_L g5532 ( 
.A1(n_5497),
.A2(n_5017),
.B(n_5030),
.Y(n_5532)
);

CKINVDCx20_ASAP7_75t_R g5533 ( 
.A(n_5333),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5500),
.Y(n_5534)
);

OAI21x1_ASAP7_75t_L g5535 ( 
.A1(n_5498),
.A2(n_5107),
.B(n_5115),
.Y(n_5535)
);

INVx2_ASAP7_75t_SL g5536 ( 
.A(n_5353),
.Y(n_5536)
);

OAI21x1_ASAP7_75t_L g5537 ( 
.A1(n_5503),
.A2(n_5165),
.B(n_5145),
.Y(n_5537)
);

O2A1O1Ixp33_ASAP7_75t_L g5538 ( 
.A1(n_5492),
.A2(n_5236),
.B(n_5010),
.C(n_5224),
.Y(n_5538)
);

OAI21xp5_ASAP7_75t_L g5539 ( 
.A1(n_5411),
.A2(n_5274),
.B(n_5217),
.Y(n_5539)
);

AND2x6_ASAP7_75t_L g5540 ( 
.A(n_5362),
.B(n_5114),
.Y(n_5540)
);

NAND2xp5_ASAP7_75t_L g5541 ( 
.A(n_5415),
.B(n_5124),
.Y(n_5541)
);

OAI21xp5_ASAP7_75t_L g5542 ( 
.A1(n_5504),
.A2(n_5136),
.B(n_5316),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_5419),
.B(n_5056),
.Y(n_5543)
);

OAI21x1_ASAP7_75t_L g5544 ( 
.A1(n_5396),
.A2(n_5016),
.B(n_5092),
.Y(n_5544)
);

AOI21xp5_ASAP7_75t_L g5545 ( 
.A1(n_5489),
.A2(n_5284),
.B(n_5096),
.Y(n_5545)
);

INVx2_ASAP7_75t_SL g5546 ( 
.A(n_5339),
.Y(n_5546)
);

AND2x2_ASAP7_75t_L g5547 ( 
.A(n_5456),
.B(n_5013),
.Y(n_5547)
);

OAI22xp5_ASAP7_75t_L g5548 ( 
.A1(n_5375),
.A2(n_5171),
.B1(n_5182),
.B2(n_5200),
.Y(n_5548)
);

NOR2xp33_ASAP7_75t_SL g5549 ( 
.A(n_5339),
.B(n_5196),
.Y(n_5549)
);

OAI21x1_ASAP7_75t_L g5550 ( 
.A1(n_5493),
.A2(n_5253),
.B(n_5166),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_5425),
.B(n_5062),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5331),
.Y(n_5552)
);

O2A1O1Ixp33_ASAP7_75t_L g5553 ( 
.A1(n_5355),
.A2(n_5169),
.B(n_5312),
.C(n_5243),
.Y(n_5553)
);

AO21x2_ASAP7_75t_L g5554 ( 
.A1(n_5429),
.A2(n_5139),
.B(n_5134),
.Y(n_5554)
);

OAI21x1_ASAP7_75t_L g5555 ( 
.A1(n_5471),
.A2(n_5198),
.B(n_5168),
.Y(n_5555)
);

CKINVDCx20_ASAP7_75t_R g5556 ( 
.A(n_5349),
.Y(n_5556)
);

AOI21x1_ASAP7_75t_L g5557 ( 
.A1(n_5367),
.A2(n_5306),
.B(n_5276),
.Y(n_5557)
);

BUFx12f_ASAP7_75t_L g5558 ( 
.A(n_5352),
.Y(n_5558)
);

OAI21x1_ASAP7_75t_L g5559 ( 
.A1(n_5438),
.A2(n_5021),
.B(n_5176),
.Y(n_5559)
);

NOR2xp67_ASAP7_75t_L g5560 ( 
.A(n_5345),
.B(n_5277),
.Y(n_5560)
);

AOI21xp5_ASAP7_75t_L g5561 ( 
.A1(n_5345),
.A2(n_4621),
.B(n_5139),
.Y(n_5561)
);

OAI21x1_ASAP7_75t_L g5562 ( 
.A1(n_5478),
.A2(n_5320),
.B(n_5299),
.Y(n_5562)
);

INVx4_ASAP7_75t_L g5563 ( 
.A(n_5383),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5347),
.Y(n_5564)
);

BUFx3_ASAP7_75t_L g5565 ( 
.A(n_5343),
.Y(n_5565)
);

AND2x2_ASAP7_75t_L g5566 ( 
.A(n_5397),
.B(n_5430),
.Y(n_5566)
);

OAI22xp5_ASAP7_75t_L g5567 ( 
.A1(n_5408),
.A2(n_5203),
.B1(n_5024),
.B2(n_5162),
.Y(n_5567)
);

INVx1_ASAP7_75t_SL g5568 ( 
.A(n_5385),
.Y(n_5568)
);

OAI21xp5_ASAP7_75t_L g5569 ( 
.A1(n_5510),
.A2(n_5133),
.B(n_5307),
.Y(n_5569)
);

AOI21x1_ASAP7_75t_L g5570 ( 
.A1(n_5482),
.A2(n_5337),
.B(n_5465),
.Y(n_5570)
);

BUFx4f_ASAP7_75t_L g5571 ( 
.A(n_5437),
.Y(n_5571)
);

HB1xp67_ASAP7_75t_L g5572 ( 
.A(n_5389),
.Y(n_5572)
);

OAI21x1_ASAP7_75t_L g5573 ( 
.A1(n_5490),
.A2(n_5279),
.B(n_5193),
.Y(n_5573)
);

BUFx2_ASAP7_75t_L g5574 ( 
.A(n_5395),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5363),
.Y(n_5575)
);

OAI21x1_ASAP7_75t_L g5576 ( 
.A1(n_5379),
.A2(n_5192),
.B(n_5147),
.Y(n_5576)
);

AOI22xp5_ASAP7_75t_L g5577 ( 
.A1(n_5449),
.A2(n_4793),
.B1(n_4631),
.B2(n_4636),
.Y(n_5577)
);

OAI21x1_ASAP7_75t_L g5578 ( 
.A1(n_5499),
.A2(n_5125),
.B(n_5119),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_L g5579 ( 
.A(n_5405),
.B(n_5126),
.Y(n_5579)
);

AOI21xp5_ASAP7_75t_L g5580 ( 
.A1(n_5358),
.A2(n_4621),
.B(n_5116),
.Y(n_5580)
);

OAI21x1_ASAP7_75t_L g5581 ( 
.A1(n_5495),
.A2(n_5130),
.B(n_5135),
.Y(n_5581)
);

NAND3xp33_ASAP7_75t_L g5582 ( 
.A(n_5483),
.B(n_5256),
.C(n_5252),
.Y(n_5582)
);

OAI21x1_ASAP7_75t_SL g5583 ( 
.A1(n_5328),
.A2(n_5298),
.B(n_5255),
.Y(n_5583)
);

OAI21x1_ASAP7_75t_L g5584 ( 
.A1(n_5371),
.A2(n_5038),
.B(n_5132),
.Y(n_5584)
);

OAI21x1_ASAP7_75t_L g5585 ( 
.A1(n_5502),
.A2(n_5142),
.B(n_4805),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5332),
.B(n_5181),
.Y(n_5586)
);

A2O1A1Ixp33_ASAP7_75t_L g5587 ( 
.A1(n_5453),
.A2(n_5302),
.B(n_5177),
.C(n_5187),
.Y(n_5587)
);

OAI21x1_ASAP7_75t_L g5588 ( 
.A1(n_5505),
.A2(n_5202),
.B(n_5216),
.Y(n_5588)
);

NAND2x1p5_ASAP7_75t_L g5589 ( 
.A(n_5358),
.B(n_5248),
.Y(n_5589)
);

OAI21x1_ASAP7_75t_L g5590 ( 
.A1(n_5336),
.A2(n_5157),
.B(n_5258),
.Y(n_5590)
);

INVx3_ASAP7_75t_L g5591 ( 
.A(n_5350),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5404),
.Y(n_5592)
);

NOR2xp33_ASAP7_75t_L g5593 ( 
.A(n_5341),
.B(n_5257),
.Y(n_5593)
);

OAI21xp5_ASAP7_75t_L g5594 ( 
.A1(n_5464),
.A2(n_5186),
.B(n_5321),
.Y(n_5594)
);

OR2x6_ASAP7_75t_L g5595 ( 
.A(n_5399),
.B(n_5118),
.Y(n_5595)
);

OAI21x1_ASAP7_75t_L g5596 ( 
.A1(n_5473),
.A2(n_5242),
.B(n_5222),
.Y(n_5596)
);

OAI22xp5_ASAP7_75t_L g5597 ( 
.A1(n_5486),
.A2(n_5110),
.B1(n_4816),
.B2(n_4823),
.Y(n_5597)
);

AOI22xp5_ASAP7_75t_L g5598 ( 
.A1(n_5449),
.A2(n_4616),
.B1(n_5308),
.B2(n_4914),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5342),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5401),
.Y(n_5600)
);

AND2x2_ASAP7_75t_L g5601 ( 
.A(n_5390),
.B(n_5268),
.Y(n_5601)
);

OAI21x1_ASAP7_75t_L g5602 ( 
.A1(n_5474),
.A2(n_5158),
.B(n_5317),
.Y(n_5602)
);

O2A1O1Ixp33_ASAP7_75t_SL g5603 ( 
.A1(n_5361),
.A2(n_4982),
.B(n_4897),
.C(n_4775),
.Y(n_5603)
);

OA21x2_ASAP7_75t_L g5604 ( 
.A1(n_5426),
.A2(n_5213),
.B(n_5207),
.Y(n_5604)
);

OA21x2_ASAP7_75t_L g5605 ( 
.A1(n_5431),
.A2(n_5265),
.B(n_5264),
.Y(n_5605)
);

OAI21x1_ASAP7_75t_L g5606 ( 
.A1(n_5485),
.A2(n_5506),
.B(n_5466),
.Y(n_5606)
);

NOR2xp33_ASAP7_75t_L g5607 ( 
.A(n_5327),
.B(n_5273),
.Y(n_5607)
);

OAI21x1_ASAP7_75t_L g5608 ( 
.A1(n_5325),
.A2(n_5300),
.B(n_5183),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_5403),
.Y(n_5609)
);

AO21x2_ASAP7_75t_L g5610 ( 
.A1(n_5372),
.A2(n_4728),
.B(n_4718),
.Y(n_5610)
);

OAI21x1_ASAP7_75t_L g5611 ( 
.A1(n_5357),
.A2(n_5226),
.B(n_5225),
.Y(n_5611)
);

INVx6_ASAP7_75t_L g5612 ( 
.A(n_5364),
.Y(n_5612)
);

INVx2_ASAP7_75t_L g5613 ( 
.A(n_5359),
.Y(n_5613)
);

AOI21xp5_ASAP7_75t_L g5614 ( 
.A1(n_5364),
.A2(n_4621),
.B(n_4953),
.Y(n_5614)
);

INVx3_ASAP7_75t_L g5615 ( 
.A(n_5374),
.Y(n_5615)
);

INVx2_ASAP7_75t_L g5616 ( 
.A(n_5360),
.Y(n_5616)
);

AND2x2_ASAP7_75t_L g5617 ( 
.A(n_5417),
.B(n_5268),
.Y(n_5617)
);

OA21x2_ASAP7_75t_L g5618 ( 
.A1(n_5338),
.A2(n_5287),
.B(n_5275),
.Y(n_5618)
);

OAI21x1_ASAP7_75t_L g5619 ( 
.A1(n_5378),
.A2(n_5234),
.B(n_5228),
.Y(n_5619)
);

OAI21xp5_ASAP7_75t_L g5620 ( 
.A1(n_5420),
.A2(n_5288),
.B(n_4784),
.Y(n_5620)
);

AO21x2_ASAP7_75t_L g5621 ( 
.A1(n_5348),
.A2(n_4734),
.B(n_4729),
.Y(n_5621)
);

OAI21x1_ASAP7_75t_L g5622 ( 
.A1(n_5388),
.A2(n_5294),
.B(n_5281),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_5418),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5424),
.Y(n_5624)
);

OAI21xp5_ASAP7_75t_L g5625 ( 
.A1(n_5508),
.A2(n_4923),
.B(n_5208),
.Y(n_5625)
);

NOR2xp33_ASAP7_75t_L g5626 ( 
.A(n_5511),
.B(n_5304),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5410),
.Y(n_5627)
);

CKINVDCx5p33_ASAP7_75t_R g5628 ( 
.A(n_5433),
.Y(n_5628)
);

NOR2x1_ASAP7_75t_R g5629 ( 
.A(n_5416),
.B(n_5323),
.Y(n_5629)
);

OAI21xp5_ASAP7_75t_L g5630 ( 
.A1(n_5432),
.A2(n_4907),
.B(n_5295),
.Y(n_5630)
);

OAI21x1_ASAP7_75t_L g5631 ( 
.A1(n_5412),
.A2(n_5313),
.B(n_5219),
.Y(n_5631)
);

INVx3_ASAP7_75t_L g5632 ( 
.A(n_5374),
.Y(n_5632)
);

OAI21x1_ASAP7_75t_L g5633 ( 
.A1(n_5448),
.A2(n_5249),
.B(n_5179),
.Y(n_5633)
);

HB1xp67_ASAP7_75t_L g5634 ( 
.A(n_5340),
.Y(n_5634)
);

NOR2xp33_ASAP7_75t_L g5635 ( 
.A(n_5511),
.B(n_4759),
.Y(n_5635)
);

OA21x2_ASAP7_75t_L g5636 ( 
.A1(n_5477),
.A2(n_4856),
.B(n_4761),
.Y(n_5636)
);

AND2x4_ASAP7_75t_L g5637 ( 
.A(n_5335),
.B(n_5194),
.Y(n_5637)
);

OAI21xp5_ASAP7_75t_L g5638 ( 
.A1(n_5475),
.A2(n_4785),
.B(n_4778),
.Y(n_5638)
);

INVx2_ASAP7_75t_L g5639 ( 
.A(n_5443),
.Y(n_5639)
);

CKINVDCx5p33_ASAP7_75t_R g5640 ( 
.A(n_5368),
.Y(n_5640)
);

INVx6_ASAP7_75t_L g5641 ( 
.A(n_5382),
.Y(n_5641)
);

OAI21x1_ASAP7_75t_L g5642 ( 
.A1(n_5369),
.A2(n_5261),
.B(n_5259),
.Y(n_5642)
);

OAI21x1_ASAP7_75t_L g5643 ( 
.A1(n_5326),
.A2(n_5462),
.B(n_5427),
.Y(n_5643)
);

NAND2xp5_ASAP7_75t_L g5644 ( 
.A(n_5459),
.B(n_5435),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5572),
.Y(n_5645)
);

INVx1_ASAP7_75t_SL g5646 ( 
.A(n_5525),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5606),
.Y(n_5647)
);

AOI22xp33_ASAP7_75t_L g5648 ( 
.A1(n_5524),
.A2(n_5486),
.B1(n_5441),
.B2(n_5491),
.Y(n_5648)
);

BUFx2_ASAP7_75t_L g5649 ( 
.A(n_5516),
.Y(n_5649)
);

BUFx2_ASAP7_75t_SL g5650 ( 
.A(n_5521),
.Y(n_5650)
);

OAI21x1_ASAP7_75t_L g5651 ( 
.A1(n_5570),
.A2(n_5414),
.B(n_5436),
.Y(n_5651)
);

INVx1_ASAP7_75t_SL g5652 ( 
.A(n_5565),
.Y(n_5652)
);

HB1xp67_ASAP7_75t_L g5653 ( 
.A(n_5516),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5627),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5566),
.Y(n_5655)
);

INVx2_ASAP7_75t_L g5656 ( 
.A(n_5518),
.Y(n_5656)
);

INVx2_ASAP7_75t_SL g5657 ( 
.A(n_5513),
.Y(n_5657)
);

BUFx3_ASAP7_75t_L g5658 ( 
.A(n_5571),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5600),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_5574),
.Y(n_5660)
);

INVx1_ASAP7_75t_SL g5661 ( 
.A(n_5556),
.Y(n_5661)
);

AND2x2_ASAP7_75t_L g5662 ( 
.A(n_5574),
.B(n_5442),
.Y(n_5662)
);

OAI22xp5_ASAP7_75t_L g5663 ( 
.A1(n_5519),
.A2(n_5467),
.B1(n_5392),
.B2(n_5452),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5609),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5623),
.Y(n_5665)
);

AND2x2_ASAP7_75t_L g5666 ( 
.A(n_5634),
.B(n_5356),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_5522),
.Y(n_5667)
);

INVx2_ASAP7_75t_L g5668 ( 
.A(n_5643),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_5599),
.Y(n_5669)
);

INVx2_ASAP7_75t_L g5670 ( 
.A(n_5613),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5552),
.Y(n_5671)
);

OAI21x1_ASAP7_75t_L g5672 ( 
.A1(n_5523),
.A2(n_5461),
.B(n_5446),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_5616),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5564),
.Y(n_5674)
);

INVx1_ASAP7_75t_SL g5675 ( 
.A(n_5514),
.Y(n_5675)
);

OAI22xp33_ASAP7_75t_L g5676 ( 
.A1(n_5549),
.A2(n_5382),
.B1(n_5454),
.B2(n_5394),
.Y(n_5676)
);

AOI22xp33_ASAP7_75t_L g5677 ( 
.A1(n_5637),
.A2(n_5509),
.B1(n_5413),
.B2(n_5457),
.Y(n_5677)
);

INVx1_ASAP7_75t_SL g5678 ( 
.A(n_5529),
.Y(n_5678)
);

INVx2_ASAP7_75t_L g5679 ( 
.A(n_5586),
.Y(n_5679)
);

HB1xp67_ASAP7_75t_L g5680 ( 
.A(n_5617),
.Y(n_5680)
);

BUFx3_ASAP7_75t_L g5681 ( 
.A(n_5558),
.Y(n_5681)
);

HB1xp67_ASAP7_75t_L g5682 ( 
.A(n_5618),
.Y(n_5682)
);

BUFx2_ASAP7_75t_L g5683 ( 
.A(n_5546),
.Y(n_5683)
);

NOR2xp33_ASAP7_75t_L g5684 ( 
.A(n_5563),
.B(n_5487),
.Y(n_5684)
);

INVx3_ASAP7_75t_L g5685 ( 
.A(n_5612),
.Y(n_5685)
);

INVx4_ASAP7_75t_L g5686 ( 
.A(n_5628),
.Y(n_5686)
);

OA21x2_ASAP7_75t_L g5687 ( 
.A1(n_5532),
.A2(n_5472),
.B(n_5469),
.Y(n_5687)
);

BUFx5_ASAP7_75t_L g5688 ( 
.A(n_5540),
.Y(n_5688)
);

OAI21x1_ASAP7_75t_L g5689 ( 
.A1(n_5535),
.A2(n_5402),
.B(n_5354),
.Y(n_5689)
);

BUFx5_ASAP7_75t_L g5690 ( 
.A(n_5540),
.Y(n_5690)
);

INVx4_ASAP7_75t_L g5691 ( 
.A(n_5591),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5575),
.Y(n_5692)
);

AND2x4_ASAP7_75t_L g5693 ( 
.A(n_5551),
.B(n_5398),
.Y(n_5693)
);

INVx6_ASAP7_75t_L g5694 ( 
.A(n_5612),
.Y(n_5694)
);

INVx2_ASAP7_75t_L g5695 ( 
.A(n_5592),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_5624),
.Y(n_5696)
);

INVx2_ASAP7_75t_L g5697 ( 
.A(n_5543),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5644),
.Y(n_5698)
);

NAND2xp5_ASAP7_75t_L g5699 ( 
.A(n_5601),
.B(n_5470),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5541),
.Y(n_5700)
);

OAI21x1_ASAP7_75t_L g5701 ( 
.A1(n_5544),
.A2(n_5269),
.B(n_5267),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5547),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5579),
.Y(n_5703)
);

INVx4_ASAP7_75t_L g5704 ( 
.A(n_5640),
.Y(n_5704)
);

INVx1_ASAP7_75t_SL g5705 ( 
.A(n_5568),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5618),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5605),
.Y(n_5707)
);

OAI22xp5_ASAP7_75t_SL g5708 ( 
.A1(n_5533),
.A2(n_5381),
.B1(n_5380),
.B2(n_5447),
.Y(n_5708)
);

HB1xp67_ASAP7_75t_L g5709 ( 
.A(n_5605),
.Y(n_5709)
);

BUFx3_ASAP7_75t_L g5710 ( 
.A(n_5536),
.Y(n_5710)
);

AOI22xp33_ASAP7_75t_L g5711 ( 
.A1(n_5540),
.A2(n_5476),
.B1(n_5479),
.B2(n_5496),
.Y(n_5711)
);

BUFx6f_ASAP7_75t_SL g5712 ( 
.A(n_5512),
.Y(n_5712)
);

BUFx2_ASAP7_75t_L g5713 ( 
.A(n_5641),
.Y(n_5713)
);

HB1xp67_ASAP7_75t_L g5714 ( 
.A(n_5604),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_5639),
.B(n_5445),
.Y(n_5715)
);

AOI22xp5_ASAP7_75t_L g5716 ( 
.A1(n_5520),
.A2(n_5440),
.B1(n_5366),
.B2(n_5373),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_5604),
.Y(n_5717)
);

AOI22xp33_ASAP7_75t_L g5718 ( 
.A1(n_5569),
.A2(n_5501),
.B1(n_5496),
.B2(n_5393),
.Y(n_5718)
);

INVx3_ASAP7_75t_L g5719 ( 
.A(n_5641),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5636),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5636),
.Y(n_5721)
);

OAI21xp5_ASAP7_75t_L g5722 ( 
.A1(n_5530),
.A2(n_5545),
.B(n_5539),
.Y(n_5722)
);

INVx3_ASAP7_75t_L g5723 ( 
.A(n_5615),
.Y(n_5723)
);

INVx6_ASAP7_75t_L g5724 ( 
.A(n_5512),
.Y(n_5724)
);

OA21x2_ASAP7_75t_L g5725 ( 
.A1(n_5590),
.A2(n_4917),
.B(n_4909),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5621),
.Y(n_5726)
);

BUFx3_ASAP7_75t_L g5727 ( 
.A(n_5632),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_5527),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5596),
.Y(n_5729)
);

AOI22xp33_ASAP7_75t_L g5730 ( 
.A1(n_5595),
.A2(n_5501),
.B1(n_5444),
.B2(n_5488),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_5528),
.Y(n_5731)
);

INVx2_ASAP7_75t_L g5732 ( 
.A(n_5534),
.Y(n_5732)
);

BUFx2_ASAP7_75t_L g5733 ( 
.A(n_5595),
.Y(n_5733)
);

AOI22xp33_ASAP7_75t_SL g5734 ( 
.A1(n_5583),
.A2(n_5370),
.B1(n_5454),
.B2(n_5394),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_L g5735 ( 
.A1(n_5625),
.A2(n_5148),
.B1(n_5143),
.B2(n_4996),
.Y(n_5735)
);

OAI22xp33_ASAP7_75t_L g5736 ( 
.A1(n_5560),
.A2(n_5439),
.B1(n_5400),
.B2(n_5406),
.Y(n_5736)
);

BUFx3_ASAP7_75t_L g5737 ( 
.A(n_5593),
.Y(n_5737)
);

INVx2_ASAP7_75t_L g5738 ( 
.A(n_5517),
.Y(n_5738)
);

BUFx4f_ASAP7_75t_SL g5739 ( 
.A(n_5629),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5517),
.Y(n_5740)
);

INVx5_ASAP7_75t_L g5741 ( 
.A(n_5557),
.Y(n_5741)
);

BUFx12f_ASAP7_75t_L g5742 ( 
.A(n_5589),
.Y(n_5742)
);

AOI21x1_ASAP7_75t_L g5743 ( 
.A1(n_5555),
.A2(n_4769),
.B(n_4760),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5610),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5550),
.Y(n_5745)
);

OAI22xp33_ASAP7_75t_L g5746 ( 
.A1(n_5567),
.A2(n_5400),
.B1(n_5406),
.B2(n_5507),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5537),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5633),
.Y(n_5748)
);

INVx4_ASAP7_75t_L g5749 ( 
.A(n_5531),
.Y(n_5749)
);

HB1xp67_ASAP7_75t_L g5750 ( 
.A(n_5642),
.Y(n_5750)
);

CKINVDCx11_ASAP7_75t_R g5751 ( 
.A(n_5548),
.Y(n_5751)
);

HB1xp67_ASAP7_75t_L g5752 ( 
.A(n_5608),
.Y(n_5752)
);

NAND2xp5_ASAP7_75t_L g5753 ( 
.A(n_5582),
.B(n_5423),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5584),
.Y(n_5754)
);

AND2x4_ASAP7_75t_L g5755 ( 
.A(n_5626),
.B(n_5423),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5588),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5515),
.Y(n_5757)
);

HB1xp67_ASAP7_75t_L g5758 ( 
.A(n_5622),
.Y(n_5758)
);

INVx2_ASAP7_75t_L g5759 ( 
.A(n_5515),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5573),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_5631),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_5559),
.Y(n_5762)
);

OAI22xp33_ASAP7_75t_R g5763 ( 
.A1(n_5607),
.A2(n_5194),
.B1(n_4586),
.B2(n_4670),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_5562),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5554),
.Y(n_5765)
);

BUFx2_ASAP7_75t_L g5766 ( 
.A(n_5581),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5635),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_5576),
.Y(n_5768)
);

AOI22xp33_ASAP7_75t_SL g5769 ( 
.A1(n_5526),
.A2(n_5480),
.B1(n_5434),
.B2(n_5450),
.Y(n_5769)
);

INVx2_ASAP7_75t_SL g5770 ( 
.A(n_5585),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5578),
.Y(n_5771)
);

BUFx6f_ASAP7_75t_L g5772 ( 
.A(n_5611),
.Y(n_5772)
);

INVx5_ASAP7_75t_SL g5773 ( 
.A(n_5650),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5649),
.Y(n_5774)
);

AND2x2_ASAP7_75t_L g5775 ( 
.A(n_5683),
.B(n_5713),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5649),
.Y(n_5776)
);

BUFx2_ASAP7_75t_L g5777 ( 
.A(n_5653),
.Y(n_5777)
);

AND2x2_ASAP7_75t_L g5778 ( 
.A(n_5683),
.B(n_5434),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5669),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5706),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5645),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5670),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_5713),
.B(n_5450),
.Y(n_5783)
);

NAND2x1p5_ASAP7_75t_L g5784 ( 
.A(n_5691),
.B(n_5422),
.Y(n_5784)
);

OR2x6_ASAP7_75t_L g5785 ( 
.A(n_5742),
.B(n_5594),
.Y(n_5785)
);

HB1xp67_ASAP7_75t_L g5786 ( 
.A(n_5660),
.Y(n_5786)
);

OAI21x1_ASAP7_75t_L g5787 ( 
.A1(n_5651),
.A2(n_5689),
.B(n_5672),
.Y(n_5787)
);

AOI22xp5_ASAP7_75t_L g5788 ( 
.A1(n_5763),
.A2(n_5598),
.B1(n_5577),
.B2(n_5597),
.Y(n_5788)
);

OAI22xp5_ASAP7_75t_L g5789 ( 
.A1(n_5733),
.A2(n_5587),
.B1(n_5542),
.B2(n_5638),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5673),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5720),
.Y(n_5791)
);

INVx4_ASAP7_75t_L g5792 ( 
.A(n_5658),
.Y(n_5792)
);

INVx2_ASAP7_75t_L g5793 ( 
.A(n_5656),
.Y(n_5793)
);

OR2x2_ASAP7_75t_L g5794 ( 
.A(n_5700),
.B(n_5458),
.Y(n_5794)
);

INVx2_ASAP7_75t_L g5795 ( 
.A(n_5728),
.Y(n_5795)
);

HB1xp67_ASAP7_75t_L g5796 ( 
.A(n_5721),
.Y(n_5796)
);

INVx1_ASAP7_75t_L g5797 ( 
.A(n_5682),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5695),
.Y(n_5798)
);

NAND2xp5_ASAP7_75t_L g5799 ( 
.A(n_5707),
.B(n_5538),
.Y(n_5799)
);

BUFx3_ASAP7_75t_L g5800 ( 
.A(n_5681),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5731),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5654),
.Y(n_5802)
);

INVx2_ASAP7_75t_L g5803 ( 
.A(n_5732),
.Y(n_5803)
);

AOI22xp33_ASAP7_75t_L g5804 ( 
.A1(n_5751),
.A2(n_5620),
.B1(n_5630),
.B2(n_5619),
.Y(n_5804)
);

BUFx2_ASAP7_75t_R g5805 ( 
.A(n_5710),
.Y(n_5805)
);

INVx2_ASAP7_75t_L g5806 ( 
.A(n_5679),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5761),
.Y(n_5807)
);

BUFx3_ASAP7_75t_L g5808 ( 
.A(n_5657),
.Y(n_5808)
);

INVx2_ASAP7_75t_SL g5809 ( 
.A(n_5652),
.Y(n_5809)
);

OR2x2_ASAP7_75t_L g5810 ( 
.A(n_5703),
.B(n_5458),
.Y(n_5810)
);

INVx2_ASAP7_75t_SL g5811 ( 
.A(n_5694),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5659),
.Y(n_5812)
);

AND2x2_ASAP7_75t_L g5813 ( 
.A(n_5733),
.B(n_5463),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5664),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5667),
.Y(n_5815)
);

HB1xp67_ASAP7_75t_L g5816 ( 
.A(n_5666),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_5671),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5748),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5655),
.Y(n_5819)
);

AND2x4_ASAP7_75t_L g5820 ( 
.A(n_5770),
.B(n_5463),
.Y(n_5820)
);

BUFx3_ASAP7_75t_L g5821 ( 
.A(n_5678),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5674),
.Y(n_5822)
);

INVx2_ASAP7_75t_SL g5823 ( 
.A(n_5694),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5692),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5696),
.Y(n_5825)
);

AOI22xp33_ASAP7_75t_SL g5826 ( 
.A1(n_5722),
.A2(n_5602),
.B1(n_5507),
.B2(n_5407),
.Y(n_5826)
);

INVx3_ASAP7_75t_L g5827 ( 
.A(n_5712),
.Y(n_5827)
);

NAND2x1p5_ASAP7_75t_L g5828 ( 
.A(n_5727),
.B(n_5422),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5665),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5717),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_5726),
.Y(n_5831)
);

AOI22xp33_ASAP7_75t_L g5832 ( 
.A1(n_5648),
.A2(n_5580),
.B1(n_5561),
.B2(n_5614),
.Y(n_5832)
);

INVx1_ASAP7_75t_SL g5833 ( 
.A(n_5661),
.Y(n_5833)
);

AO21x2_ASAP7_75t_L g5834 ( 
.A1(n_5757),
.A2(n_4947),
.B(n_4946),
.Y(n_5834)
);

BUFx2_ASAP7_75t_L g5835 ( 
.A(n_5687),
.Y(n_5835)
);

INVx3_ASAP7_75t_L g5836 ( 
.A(n_5724),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5698),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5709),
.Y(n_5838)
);

INVx2_ASAP7_75t_L g5839 ( 
.A(n_5729),
.Y(n_5839)
);

INVx2_ASAP7_75t_L g5840 ( 
.A(n_5647),
.Y(n_5840)
);

INVx2_ASAP7_75t_L g5841 ( 
.A(n_5756),
.Y(n_5841)
);

BUFx2_ASAP7_75t_L g5842 ( 
.A(n_5687),
.Y(n_5842)
);

BUFx3_ASAP7_75t_L g5843 ( 
.A(n_5686),
.Y(n_5843)
);

AOI21x1_ASAP7_75t_L g5844 ( 
.A1(n_5759),
.A2(n_4959),
.B(n_4813),
.Y(n_5844)
);

INVx2_ASAP7_75t_L g5845 ( 
.A(n_5760),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5714),
.Y(n_5846)
);

INVx3_ASAP7_75t_L g5847 ( 
.A(n_5724),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5771),
.Y(n_5848)
);

AND2x4_ASAP7_75t_L g5849 ( 
.A(n_5693),
.B(n_5460),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5662),
.Y(n_5850)
);

AND2x2_ASAP7_75t_L g5851 ( 
.A(n_5677),
.B(n_5460),
.Y(n_5851)
);

OR2x2_ASAP7_75t_L g5852 ( 
.A(n_5697),
.B(n_5407),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5744),
.Y(n_5853)
);

AO21x2_ASAP7_75t_L g5854 ( 
.A1(n_5765),
.A2(n_4885),
.B(n_4855),
.Y(n_5854)
);

INVx1_ASAP7_75t_L g5855 ( 
.A(n_5768),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5745),
.Y(n_5856)
);

AOI222xp33_ASAP7_75t_L g5857 ( 
.A1(n_5739),
.A2(n_4889),
.B1(n_4900),
.B2(n_4755),
.C1(n_4783),
.C2(n_4794),
.Y(n_5857)
);

CKINVDCx5p33_ASAP7_75t_R g5858 ( 
.A(n_5646),
.Y(n_5858)
);

BUFx3_ASAP7_75t_L g5859 ( 
.A(n_5684),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5758),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_5738),
.Y(n_5861)
);

AOI21xp5_ASAP7_75t_L g5862 ( 
.A1(n_5676),
.A2(n_5603),
.B(n_5553),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5740),
.Y(n_5863)
);

NOR2xp33_ASAP7_75t_L g5864 ( 
.A(n_5704),
.B(n_5365),
.Y(n_5864)
);

AND2x4_ASAP7_75t_L g5865 ( 
.A(n_5723),
.B(n_5719),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5764),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5747),
.Y(n_5867)
);

AND2x2_ASAP7_75t_L g5868 ( 
.A(n_5685),
.B(n_5675),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5702),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5668),
.Y(n_5870)
);

INVxp67_ASAP7_75t_SL g5871 ( 
.A(n_5752),
.Y(n_5871)
);

OR2x2_ASAP7_75t_L g5872 ( 
.A(n_5680),
.B(n_5384),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5753),
.Y(n_5873)
);

AND2x4_ASAP7_75t_L g5874 ( 
.A(n_5755),
.B(n_5365),
.Y(n_5874)
);

OAI21x1_ASAP7_75t_L g5875 ( 
.A1(n_5754),
.A2(n_5762),
.B(n_5663),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5772),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5750),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5699),
.Y(n_5878)
);

AOI22xp33_ASAP7_75t_SL g5879 ( 
.A1(n_5789),
.A2(n_5688),
.B1(n_5690),
.B2(n_5741),
.Y(n_5879)
);

AND2x2_ASAP7_75t_L g5880 ( 
.A(n_5775),
.B(n_5688),
.Y(n_5880)
);

OAI21x1_ASAP7_75t_L g5881 ( 
.A1(n_5875),
.A2(n_5730),
.B(n_5718),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5797),
.Y(n_5882)
);

INVx2_ASAP7_75t_SL g5883 ( 
.A(n_5821),
.Y(n_5883)
);

BUFx3_ASAP7_75t_L g5884 ( 
.A(n_5800),
.Y(n_5884)
);

INVx2_ASAP7_75t_L g5885 ( 
.A(n_5777),
.Y(n_5885)
);

AO21x2_ASAP7_75t_L g5886 ( 
.A1(n_5799),
.A2(n_5746),
.B(n_5743),
.Y(n_5886)
);

AO21x2_ASAP7_75t_L g5887 ( 
.A1(n_5860),
.A2(n_5743),
.B(n_5716),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5777),
.Y(n_5888)
);

INVx3_ASAP7_75t_L g5889 ( 
.A(n_5773),
.Y(n_5889)
);

OR2x6_ASAP7_75t_L g5890 ( 
.A(n_5827),
.B(n_5708),
.Y(n_5890)
);

INVx3_ASAP7_75t_L g5891 ( 
.A(n_5773),
.Y(n_5891)
);

BUFx2_ASAP7_75t_L g5892 ( 
.A(n_5785),
.Y(n_5892)
);

AOI21x1_ASAP7_75t_L g5893 ( 
.A1(n_5785),
.A2(n_5766),
.B(n_5725),
.Y(n_5893)
);

HB1xp67_ASAP7_75t_L g5894 ( 
.A(n_5796),
.Y(n_5894)
);

AO21x2_ASAP7_75t_L g5895 ( 
.A1(n_5860),
.A2(n_5877),
.B(n_5871),
.Y(n_5895)
);

AND2x2_ASAP7_75t_L g5896 ( 
.A(n_5836),
.B(n_5688),
.Y(n_5896)
);

AO21x2_ASAP7_75t_L g5897 ( 
.A1(n_5838),
.A2(n_5736),
.B(n_5701),
.Y(n_5897)
);

AND2x4_ASAP7_75t_L g5898 ( 
.A(n_5836),
.B(n_5737),
.Y(n_5898)
);

OA21x2_ASAP7_75t_L g5899 ( 
.A1(n_5862),
.A2(n_5766),
.B(n_5711),
.Y(n_5899)
);

INVx3_ASAP7_75t_L g5900 ( 
.A(n_5784),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5863),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5837),
.Y(n_5902)
);

INVx2_ASAP7_75t_L g5903 ( 
.A(n_5774),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_L g5904 ( 
.A(n_5832),
.B(n_5788),
.Y(n_5904)
);

OR2x2_ASAP7_75t_L g5905 ( 
.A(n_5780),
.B(n_5725),
.Y(n_5905)
);

BUFx2_ASAP7_75t_L g5906 ( 
.A(n_5827),
.Y(n_5906)
);

BUFx3_ASAP7_75t_L g5907 ( 
.A(n_5843),
.Y(n_5907)
);

INVx3_ASAP7_75t_L g5908 ( 
.A(n_5792),
.Y(n_5908)
);

INVx2_ASAP7_75t_L g5909 ( 
.A(n_5776),
.Y(n_5909)
);

AND2x2_ASAP7_75t_L g5910 ( 
.A(n_5847),
.B(n_5688),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5795),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5846),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5816),
.Y(n_5913)
);

AND2x2_ASAP7_75t_L g5914 ( 
.A(n_5847),
.B(n_5690),
.Y(n_5914)
);

NAND2xp5_ASAP7_75t_L g5915 ( 
.A(n_5781),
.B(n_5769),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_5811),
.B(n_5823),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5802),
.Y(n_5917)
);

AND2x2_ASAP7_75t_L g5918 ( 
.A(n_5868),
.B(n_5690),
.Y(n_5918)
);

AND2x2_ASAP7_75t_L g5919 ( 
.A(n_5865),
.B(n_5690),
.Y(n_5919)
);

AND2x2_ASAP7_75t_L g5920 ( 
.A(n_5865),
.B(n_5715),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5783),
.B(n_5767),
.Y(n_5921)
);

OR2x6_ASAP7_75t_L g5922 ( 
.A(n_5792),
.B(n_5734),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5812),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5814),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_5873),
.B(n_5834),
.Y(n_5925)
);

AND2x2_ASAP7_75t_L g5926 ( 
.A(n_5778),
.B(n_5705),
.Y(n_5926)
);

AOI22xp33_ASAP7_75t_L g5927 ( 
.A1(n_5804),
.A2(n_5772),
.B1(n_5735),
.B2(n_5741),
.Y(n_5927)
);

HB1xp67_ASAP7_75t_L g5928 ( 
.A(n_5830),
.Y(n_5928)
);

INVx1_ASAP7_75t_SL g5929 ( 
.A(n_5805),
.Y(n_5929)
);

NAND2xp5_ASAP7_75t_L g5930 ( 
.A(n_5878),
.B(n_5741),
.Y(n_5930)
);

INVx3_ASAP7_75t_L g5931 ( 
.A(n_5808),
.Y(n_5931)
);

INVx2_ASAP7_75t_L g5932 ( 
.A(n_5801),
.Y(n_5932)
);

OA21x2_ASAP7_75t_L g5933 ( 
.A1(n_5835),
.A2(n_5842),
.B(n_5787),
.Y(n_5933)
);

HB1xp67_ASAP7_75t_L g5934 ( 
.A(n_5791),
.Y(n_5934)
);

OAI21x1_ASAP7_75t_L g5935 ( 
.A1(n_5861),
.A2(n_5749),
.B(n_4797),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5803),
.Y(n_5936)
);

AO21x2_ASAP7_75t_L g5937 ( 
.A1(n_5853),
.A2(n_4792),
.B(n_4771),
.Y(n_5937)
);

AND2x2_ASAP7_75t_L g5938 ( 
.A(n_5851),
.B(n_5377),
.Y(n_5938)
);

AND2x2_ASAP7_75t_L g5939 ( 
.A(n_5813),
.B(n_5377),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5825),
.Y(n_5940)
);

AOI21x1_ASAP7_75t_L g5941 ( 
.A1(n_5835),
.A2(n_4834),
.B(n_4812),
.Y(n_5941)
);

INVx2_ASAP7_75t_L g5942 ( 
.A(n_5779),
.Y(n_5942)
);

INVx2_ASAP7_75t_L g5943 ( 
.A(n_5782),
.Y(n_5943)
);

INVxp33_ASAP7_75t_L g5944 ( 
.A(n_5828),
.Y(n_5944)
);

INVx2_ASAP7_75t_L g5945 ( 
.A(n_5790),
.Y(n_5945)
);

INVx2_ASAP7_75t_SL g5946 ( 
.A(n_5849),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5825),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5849),
.B(n_5384),
.Y(n_5948)
);

INVx2_ASAP7_75t_L g5949 ( 
.A(n_5793),
.Y(n_5949)
);

AND2x2_ASAP7_75t_L g5950 ( 
.A(n_5809),
.B(n_5386),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5815),
.Y(n_5951)
);

AND2x2_ASAP7_75t_L g5952 ( 
.A(n_5850),
.B(n_5386),
.Y(n_5952)
);

INVx1_ASAP7_75t_SL g5953 ( 
.A(n_5858),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5817),
.Y(n_5954)
);

BUFx2_ASAP7_75t_L g5955 ( 
.A(n_5859),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5824),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5829),
.Y(n_5957)
);

HB1xp67_ASAP7_75t_L g5958 ( 
.A(n_5845),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5869),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5822),
.Y(n_5960)
);

OR2x2_ASAP7_75t_L g5961 ( 
.A(n_5819),
.B(n_5206),
.Y(n_5961)
);

NAND2xp5_ASAP7_75t_L g5962 ( 
.A(n_5867),
.B(n_5206),
.Y(n_5962)
);

INVx2_ASAP7_75t_L g5963 ( 
.A(n_5861),
.Y(n_5963)
);

HB1xp67_ASAP7_75t_L g5964 ( 
.A(n_5839),
.Y(n_5964)
);

INVx2_ASAP7_75t_SL g5965 ( 
.A(n_5833),
.Y(n_5965)
);

OR2x2_ASAP7_75t_L g5966 ( 
.A(n_5786),
.B(n_5239),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5856),
.Y(n_5967)
);

INVx3_ASAP7_75t_L g5968 ( 
.A(n_5842),
.Y(n_5968)
);

INVx2_ASAP7_75t_L g5969 ( 
.A(n_5806),
.Y(n_5969)
);

OA21x2_ASAP7_75t_L g5970 ( 
.A1(n_5876),
.A2(n_5866),
.B(n_5841),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5848),
.Y(n_5971)
);

INVx3_ASAP7_75t_L g5972 ( 
.A(n_5874),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5798),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5818),
.Y(n_5974)
);

BUFx2_ASAP7_75t_L g5975 ( 
.A(n_5874),
.Y(n_5975)
);

OAI21xp5_ASAP7_75t_L g5976 ( 
.A1(n_5826),
.A2(n_4788),
.B(n_4845),
.Y(n_5976)
);

HB1xp67_ASAP7_75t_L g5977 ( 
.A(n_5855),
.Y(n_5977)
);

OR2x2_ASAP7_75t_L g5978 ( 
.A(n_5840),
.B(n_5239),
.Y(n_5978)
);

HB1xp67_ASAP7_75t_L g5979 ( 
.A(n_5831),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5810),
.Y(n_5980)
);

OAI21x1_ASAP7_75t_L g5981 ( 
.A1(n_5870),
.A2(n_4859),
.B(n_4847),
.Y(n_5981)
);

AND2x2_ASAP7_75t_L g5982 ( 
.A(n_5872),
.B(n_5303),
.Y(n_5982)
);

AO21x2_ASAP7_75t_L g5983 ( 
.A1(n_5807),
.A2(n_4803),
.B(n_4796),
.Y(n_5983)
);

AOI22xp33_ASAP7_75t_L g5984 ( 
.A1(n_5854),
.A2(n_4968),
.B1(n_4662),
.B2(n_4611),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5794),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5844),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5844),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5852),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5820),
.Y(n_5989)
);

INVx2_ASAP7_75t_L g5990 ( 
.A(n_5820),
.Y(n_5990)
);

INVx2_ASAP7_75t_L g5991 ( 
.A(n_5864),
.Y(n_5991)
);

HB1xp67_ASAP7_75t_L g5992 ( 
.A(n_5857),
.Y(n_5992)
);

AO21x1_ASAP7_75t_SL g5993 ( 
.A1(n_5773),
.A2(n_4948),
.B(n_4937),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5797),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5797),
.Y(n_5995)
);

HB1xp67_ASAP7_75t_L g5996 ( 
.A(n_5777),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5777),
.Y(n_5997)
);

INVx2_ASAP7_75t_L g5998 ( 
.A(n_5777),
.Y(n_5998)
);

AND2x2_ASAP7_75t_L g5999 ( 
.A(n_5775),
.B(n_5303),
.Y(n_5999)
);

AND2x2_ASAP7_75t_L g6000 ( 
.A(n_5775),
.B(n_4811),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5797),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5775),
.B(n_4826),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5830),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5799),
.B(n_4829),
.Y(n_6004)
);

BUFx6f_ASAP7_75t_L g6005 ( 
.A(n_5800),
.Y(n_6005)
);

BUFx6f_ASAP7_75t_L g6006 ( 
.A(n_5800),
.Y(n_6006)
);

OR2x2_ASAP7_75t_L g6007 ( 
.A(n_5799),
.B(n_4852),
.Y(n_6007)
);

INVx2_ASAP7_75t_L g6008 ( 
.A(n_5777),
.Y(n_6008)
);

NOR2xp67_ASAP7_75t_L g6009 ( 
.A(n_5862),
.B(n_473),
.Y(n_6009)
);

AO21x2_ASAP7_75t_L g6010 ( 
.A1(n_5799),
.A2(n_4876),
.B(n_4869),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5797),
.Y(n_6011)
);

BUFx2_ASAP7_75t_L g6012 ( 
.A(n_5785),
.Y(n_6012)
);

INVxp67_ASAP7_75t_SL g6013 ( 
.A(n_5821),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_6013),
.Y(n_6014)
);

INVx2_ASAP7_75t_SL g6015 ( 
.A(n_5884),
.Y(n_6015)
);

OR2x2_ASAP7_75t_L g6016 ( 
.A(n_5913),
.B(n_4963),
.Y(n_6016)
);

HB1xp67_ASAP7_75t_L g6017 ( 
.A(n_5996),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5955),
.Y(n_6018)
);

HB1xp67_ASAP7_75t_L g6019 ( 
.A(n_5894),
.Y(n_6019)
);

BUFx3_ASAP7_75t_L g6020 ( 
.A(n_6005),
.Y(n_6020)
);

NAND2xp5_ASAP7_75t_L g6021 ( 
.A(n_5904),
.B(n_4965),
.Y(n_6021)
);

INVx5_ASAP7_75t_L g6022 ( 
.A(n_6005),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5955),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_6010),
.B(n_4861),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5888),
.Y(n_6025)
);

OR2x2_ASAP7_75t_L g6026 ( 
.A(n_5966),
.B(n_4952),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_5965),
.Y(n_6027)
);

BUFx2_ASAP7_75t_L g6028 ( 
.A(n_5922),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5906),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5906),
.Y(n_6030)
);

NOR2x1p5_ASAP7_75t_L g6031 ( 
.A(n_5889),
.B(n_4814),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5908),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5908),
.Y(n_6033)
);

OR2x2_ASAP7_75t_L g6034 ( 
.A(n_5885),
.B(n_4978),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5883),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5928),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5931),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_5934),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5931),
.B(n_5270),
.Y(n_6039)
);

NOR2x1_ASAP7_75t_SL g6040 ( 
.A(n_5922),
.B(n_5003),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5892),
.B(n_5220),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5892),
.B(n_4993),
.Y(n_6042)
);

INVx2_ASAP7_75t_L g6043 ( 
.A(n_5997),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5998),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_6008),
.Y(n_6045)
);

INVx2_ASAP7_75t_L g6046 ( 
.A(n_5968),
.Y(n_6046)
);

INVx2_ASAP7_75t_SL g6047 ( 
.A(n_5907),
.Y(n_6047)
);

INVx2_ASAP7_75t_SL g6048 ( 
.A(n_6005),
.Y(n_6048)
);

INVx1_ASAP7_75t_L g6049 ( 
.A(n_5882),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5912),
.Y(n_6050)
);

INVx4_ASAP7_75t_L g6051 ( 
.A(n_6006),
.Y(n_6051)
);

AOI22xp33_ASAP7_75t_L g6052 ( 
.A1(n_5992),
.A2(n_4935),
.B1(n_4918),
.B2(n_4975),
.Y(n_6052)
);

INVx1_ASAP7_75t_SL g6053 ( 
.A(n_5953),
.Y(n_6053)
);

NAND2x1_ASAP7_75t_L g6054 ( 
.A(n_5975),
.B(n_4721),
.Y(n_6054)
);

INVx3_ASAP7_75t_L g6055 ( 
.A(n_6006),
.Y(n_6055)
);

INVx4_ASAP7_75t_SL g6056 ( 
.A(n_6006),
.Y(n_6056)
);

INVx2_ASAP7_75t_SL g6057 ( 
.A(n_5889),
.Y(n_6057)
);

INVx2_ASAP7_75t_SL g6058 ( 
.A(n_5891),
.Y(n_6058)
);

AND2x2_ASAP7_75t_L g6059 ( 
.A(n_6012),
.B(n_5916),
.Y(n_6059)
);

NAND2x1_ASAP7_75t_L g6060 ( 
.A(n_5975),
.B(n_4862),
.Y(n_6060)
);

AND2x4_ASAP7_75t_L g6061 ( 
.A(n_5891),
.B(n_4677),
.Y(n_6061)
);

INVxp67_ASAP7_75t_L g6062 ( 
.A(n_6012),
.Y(n_6062)
);

AOI22xp33_ASAP7_75t_L g6063 ( 
.A1(n_5890),
.A2(n_4840),
.B1(n_5238),
.B2(n_4715),
.Y(n_6063)
);

OR2x2_ASAP7_75t_L g6064 ( 
.A(n_5961),
.B(n_4998),
.Y(n_6064)
);

NOR2x1_ASAP7_75t_SL g6065 ( 
.A(n_5890),
.B(n_5005),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_5994),
.Y(n_6066)
);

AND2x2_ASAP7_75t_L g6067 ( 
.A(n_5900),
.B(n_5007),
.Y(n_6067)
);

BUFx2_ASAP7_75t_L g6068 ( 
.A(n_5929),
.Y(n_6068)
);

INVx5_ASAP7_75t_L g6069 ( 
.A(n_5900),
.Y(n_6069)
);

OR2x6_ASAP7_75t_L g6070 ( 
.A(n_6009),
.B(n_4652),
.Y(n_6070)
);

INVx2_ASAP7_75t_L g6071 ( 
.A(n_5968),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5995),
.Y(n_6072)
);

INVx2_ASAP7_75t_SL g6073 ( 
.A(n_5898),
.Y(n_6073)
);

INVx2_ASAP7_75t_L g6074 ( 
.A(n_5901),
.Y(n_6074)
);

OR2x2_ASAP7_75t_L g6075 ( 
.A(n_5962),
.B(n_5009),
.Y(n_6075)
);

AND2x4_ASAP7_75t_L g6076 ( 
.A(n_5898),
.B(n_4614),
.Y(n_6076)
);

OR2x2_ASAP7_75t_L g6077 ( 
.A(n_6007),
.B(n_5978),
.Y(n_6077)
);

INVx2_ASAP7_75t_L g6078 ( 
.A(n_5963),
.Y(n_6078)
);

OR2x2_ASAP7_75t_L g6079 ( 
.A(n_6001),
.B(n_473),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_6011),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5977),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_5979),
.Y(n_6082)
);

INVx2_ASAP7_75t_SL g6083 ( 
.A(n_5926),
.Y(n_6083)
);

AND2x2_ASAP7_75t_L g6084 ( 
.A(n_5918),
.B(n_4898),
.Y(n_6084)
);

INVx2_ASAP7_75t_L g6085 ( 
.A(n_5911),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5919),
.B(n_5896),
.Y(n_6086)
);

AND2x4_ASAP7_75t_SL g6087 ( 
.A(n_5991),
.B(n_4844),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5932),
.Y(n_6088)
);

OR2x6_ASAP7_75t_L g6089 ( 
.A(n_5946),
.B(n_4782),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5902),
.Y(n_6090)
);

AND2x2_ASAP7_75t_L g6091 ( 
.A(n_5910),
.B(n_4873),
.Y(n_6091)
);

BUFx2_ASAP7_75t_L g6092 ( 
.A(n_5933),
.Y(n_6092)
);

INVx2_ASAP7_75t_L g6093 ( 
.A(n_5936),
.Y(n_6093)
);

AND2x2_ASAP7_75t_L g6094 ( 
.A(n_5914),
.B(n_4875),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5917),
.Y(n_6095)
);

AND2x2_ASAP7_75t_L g6096 ( 
.A(n_5880),
.B(n_4878),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5923),
.Y(n_6097)
);

AND2x2_ASAP7_75t_L g6098 ( 
.A(n_5972),
.B(n_4581),
.Y(n_6098)
);

INVxp67_ASAP7_75t_SL g6099 ( 
.A(n_5933),
.Y(n_6099)
);

INVx1_ASAP7_75t_SL g6100 ( 
.A(n_5950),
.Y(n_6100)
);

AND2x2_ASAP7_75t_L g6101 ( 
.A(n_5972),
.B(n_4590),
.Y(n_6101)
);

INVx1_ASAP7_75t_SL g6102 ( 
.A(n_5948),
.Y(n_6102)
);

AND2x4_ASAP7_75t_L g6103 ( 
.A(n_5920),
.B(n_4592),
.Y(n_6103)
);

INVx1_ASAP7_75t_L g6104 ( 
.A(n_5924),
.Y(n_6104)
);

BUFx2_ASAP7_75t_L g6105 ( 
.A(n_5899),
.Y(n_6105)
);

OR2x2_ASAP7_75t_L g6106 ( 
.A(n_6004),
.B(n_473),
.Y(n_6106)
);

INVx2_ASAP7_75t_L g6107 ( 
.A(n_5942),
.Y(n_6107)
);

HB1xp67_ASAP7_75t_L g6108 ( 
.A(n_5903),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_5944),
.B(n_4574),
.Y(n_6109)
);

AND2x2_ASAP7_75t_L g6110 ( 
.A(n_5999),
.B(n_4609),
.Y(n_6110)
);

AO21x2_ASAP7_75t_L g6111 ( 
.A1(n_5893),
.A2(n_4966),
.B(n_4703),
.Y(n_6111)
);

BUFx2_ASAP7_75t_L g6112 ( 
.A(n_5899),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5943),
.Y(n_6113)
);

OAI21x1_ASAP7_75t_L g6114 ( 
.A1(n_5893),
.A2(n_4825),
.B(n_4705),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_5938),
.B(n_4695),
.Y(n_6115)
);

INVx2_ASAP7_75t_L g6116 ( 
.A(n_5945),
.Y(n_6116)
);

NAND2xp5_ASAP7_75t_L g6117 ( 
.A(n_5937),
.B(n_4713),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_5982),
.B(n_4762),
.Y(n_6118)
);

INVx3_ASAP7_75t_L g6119 ( 
.A(n_5897),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_5951),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5949),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5954),
.Y(n_6122)
);

NAND2xp5_ASAP7_75t_L g6123 ( 
.A(n_5983),
.B(n_4747),
.Y(n_6123)
);

HB1xp67_ASAP7_75t_L g6124 ( 
.A(n_5909),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_5956),
.Y(n_6125)
);

AND2x2_ASAP7_75t_L g6126 ( 
.A(n_5881),
.B(n_474),
.Y(n_6126)
);

AND2x2_ASAP7_75t_L g6127 ( 
.A(n_5927),
.B(n_474),
.Y(n_6127)
);

INVx2_ASAP7_75t_SL g6128 ( 
.A(n_5939),
.Y(n_6128)
);

OR2x2_ASAP7_75t_L g6129 ( 
.A(n_5915),
.B(n_475),
.Y(n_6129)
);

CKINVDCx12_ASAP7_75t_R g6130 ( 
.A(n_5921),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5957),
.Y(n_6131)
);

AND2x4_ASAP7_75t_L g6132 ( 
.A(n_5980),
.B(n_475),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_6003),
.Y(n_6133)
);

AND2x2_ASAP7_75t_L g6134 ( 
.A(n_5989),
.B(n_475),
.Y(n_6134)
);

NAND2xp5_ASAP7_75t_L g6135 ( 
.A(n_6000),
.B(n_4940),
.Y(n_6135)
);

AND2x2_ASAP7_75t_L g6136 ( 
.A(n_5990),
.B(n_476),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_6003),
.Y(n_6137)
);

AND2x2_ASAP7_75t_L g6138 ( 
.A(n_5988),
.B(n_476),
.Y(n_6138)
);

INVx2_ASAP7_75t_L g6139 ( 
.A(n_5959),
.Y(n_6139)
);

INVx4_ASAP7_75t_L g6140 ( 
.A(n_5952),
.Y(n_6140)
);

AND2x4_ASAP7_75t_L g6141 ( 
.A(n_5985),
.B(n_476),
.Y(n_6141)
);

AO21x2_ASAP7_75t_L g6142 ( 
.A1(n_5925),
.A2(n_4853),
.B(n_4827),
.Y(n_6142)
);

AND2x2_ASAP7_75t_L g6143 ( 
.A(n_5879),
.B(n_477),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_5940),
.Y(n_6144)
);

INVx2_ASAP7_75t_SL g6145 ( 
.A(n_5930),
.Y(n_6145)
);

INVx2_ASAP7_75t_L g6146 ( 
.A(n_5969),
.Y(n_6146)
);

AND2x2_ASAP7_75t_L g6147 ( 
.A(n_6002),
.B(n_477),
.Y(n_6147)
);

BUFx2_ASAP7_75t_L g6148 ( 
.A(n_5886),
.Y(n_6148)
);

AND2x2_ASAP7_75t_L g6149 ( 
.A(n_5993),
.B(n_477),
.Y(n_6149)
);

INVx2_ASAP7_75t_L g6150 ( 
.A(n_5974),
.Y(n_6150)
);

AND2x2_ASAP7_75t_L g6151 ( 
.A(n_5993),
.B(n_478),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_5970),
.Y(n_6152)
);

NAND2xp5_ASAP7_75t_SL g6153 ( 
.A(n_5905),
.B(n_4674),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_5887),
.B(n_478),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_5970),
.Y(n_6155)
);

AO31x2_ASAP7_75t_L g6156 ( 
.A1(n_5986),
.A2(n_4958),
.A3(n_4945),
.B(n_4908),
.Y(n_6156)
);

NAND2xp5_ASAP7_75t_L g6157 ( 
.A(n_5984),
.B(n_4903),
.Y(n_6157)
);

HB1xp67_ASAP7_75t_L g6158 ( 
.A(n_5973),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_5947),
.Y(n_6159)
);

AND2x2_ASAP7_75t_L g6160 ( 
.A(n_5960),
.B(n_478),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_5973),
.Y(n_6161)
);

INVx2_ASAP7_75t_L g6162 ( 
.A(n_5987),
.Y(n_6162)
);

INVx4_ASAP7_75t_L g6163 ( 
.A(n_5895),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_5967),
.Y(n_6164)
);

NAND2xp5_ASAP7_75t_L g6165 ( 
.A(n_5971),
.B(n_5958),
.Y(n_6165)
);

NOR2xp67_ASAP7_75t_L g6166 ( 
.A(n_5964),
.B(n_5941),
.Y(n_6166)
);

AND2x2_ASAP7_75t_L g6167 ( 
.A(n_5935),
.B(n_479),
.Y(n_6167)
);

HB1xp67_ASAP7_75t_L g6168 ( 
.A(n_5981),
.Y(n_6168)
);

HB1xp67_ASAP7_75t_L g6169 ( 
.A(n_5941),
.Y(n_6169)
);

AND2x4_ASAP7_75t_L g6170 ( 
.A(n_5976),
.B(n_479),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_6013),
.Y(n_6171)
);

INVx2_ASAP7_75t_L g6172 ( 
.A(n_5955),
.Y(n_6172)
);

NAND2xp5_ASAP7_75t_L g6173 ( 
.A(n_5904),
.B(n_4919),
.Y(n_6173)
);

INVx3_ASAP7_75t_L g6174 ( 
.A(n_5884),
.Y(n_6174)
);

INVx2_ASAP7_75t_L g6175 ( 
.A(n_5955),
.Y(n_6175)
);

NAND2xp5_ASAP7_75t_L g6176 ( 
.A(n_5904),
.B(n_4920),
.Y(n_6176)
);

INVxp67_ASAP7_75t_SL g6177 ( 
.A(n_6013),
.Y(n_6177)
);

HB1xp67_ASAP7_75t_L g6178 ( 
.A(n_6014),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_6177),
.Y(n_6179)
);

INVx2_ASAP7_75t_L g6180 ( 
.A(n_6171),
.Y(n_6180)
);

AND2x4_ASAP7_75t_L g6181 ( 
.A(n_6020),
.B(n_6022),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_6018),
.Y(n_6182)
);

INVx2_ASAP7_75t_L g6183 ( 
.A(n_6023),
.Y(n_6183)
);

INVx3_ASAP7_75t_L g6184 ( 
.A(n_6174),
.Y(n_6184)
);

AND2x2_ASAP7_75t_L g6185 ( 
.A(n_6068),
.B(n_479),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_6172),
.Y(n_6186)
);

INVx4_ASAP7_75t_L g6187 ( 
.A(n_6051),
.Y(n_6187)
);

INVx1_ASAP7_75t_L g6188 ( 
.A(n_6017),
.Y(n_6188)
);

INVxp67_ASAP7_75t_SL g6189 ( 
.A(n_6068),
.Y(n_6189)
);

AND2x2_ASAP7_75t_L g6190 ( 
.A(n_6047),
.B(n_480),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_6019),
.Y(n_6191)
);

BUFx2_ASAP7_75t_L g6192 ( 
.A(n_6055),
.Y(n_6192)
);

BUFx3_ASAP7_75t_L g6193 ( 
.A(n_6015),
.Y(n_6193)
);

AND2x2_ASAP7_75t_L g6194 ( 
.A(n_6059),
.B(n_480),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_6175),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_6092),
.Y(n_6196)
);

OR2x2_ASAP7_75t_L g6197 ( 
.A(n_6062),
.B(n_480),
.Y(n_6197)
);

AND2x2_ASAP7_75t_L g6198 ( 
.A(n_6057),
.B(n_481),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_6035),
.Y(n_6199)
);

AND2x4_ASAP7_75t_L g6200 ( 
.A(n_6022),
.B(n_481),
.Y(n_6200)
);

INVx2_ASAP7_75t_L g6201 ( 
.A(n_6027),
.Y(n_6201)
);

INVx2_ASAP7_75t_L g6202 ( 
.A(n_6152),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_6058),
.B(n_481),
.Y(n_6203)
);

INVx2_ASAP7_75t_SL g6204 ( 
.A(n_6022),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_6092),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_6099),
.Y(n_6206)
);

INVx2_ASAP7_75t_L g6207 ( 
.A(n_6155),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_6029),
.Y(n_6208)
);

INVx3_ASAP7_75t_L g6209 ( 
.A(n_6140),
.Y(n_6209)
);

INVx2_ASAP7_75t_L g6210 ( 
.A(n_6032),
.Y(n_6210)
);

HB1xp67_ASAP7_75t_L g6211 ( 
.A(n_6030),
.Y(n_6211)
);

NAND2x1_ASAP7_75t_L g6212 ( 
.A(n_6028),
.B(n_4924),
.Y(n_6212)
);

AO21x2_ASAP7_75t_L g6213 ( 
.A1(n_6040),
.A2(n_4934),
.B(n_4929),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_6033),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_6162),
.Y(n_6215)
);

AND2x4_ASAP7_75t_L g6216 ( 
.A(n_6056),
.B(n_482),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_6073),
.B(n_482),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_6158),
.Y(n_6218)
);

AND2x2_ASAP7_75t_L g6219 ( 
.A(n_6037),
.B(n_483),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_6044),
.Y(n_6220)
);

AND2x2_ASAP7_75t_L g6221 ( 
.A(n_6048),
.B(n_483),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_6046),
.Y(n_6222)
);

AND2x2_ASAP7_75t_L g6223 ( 
.A(n_6053),
.B(n_483),
.Y(n_6223)
);

AND2x2_ASAP7_75t_L g6224 ( 
.A(n_6086),
.B(n_484),
.Y(n_6224)
);

INVx1_ASAP7_75t_L g6225 ( 
.A(n_6045),
.Y(n_6225)
);

INVx2_ASAP7_75t_L g6226 ( 
.A(n_6071),
.Y(n_6226)
);

AND2x2_ASAP7_75t_L g6227 ( 
.A(n_6028),
.B(n_485),
.Y(n_6227)
);

AND2x2_ASAP7_75t_L g6228 ( 
.A(n_6083),
.B(n_485),
.Y(n_6228)
);

AND2x2_ASAP7_75t_L g6229 ( 
.A(n_6143),
.B(n_486),
.Y(n_6229)
);

AND2x2_ASAP7_75t_L g6230 ( 
.A(n_6100),
.B(n_487),
.Y(n_6230)
);

AOI22xp33_ASAP7_75t_SL g6231 ( 
.A1(n_6065),
.A2(n_4970),
.B1(n_4987),
.B2(n_4986),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_6043),
.Y(n_6232)
);

AND2x2_ASAP7_75t_L g6233 ( 
.A(n_6102),
.B(n_487),
.Y(n_6233)
);

INVx2_ASAP7_75t_L g6234 ( 
.A(n_6074),
.Y(n_6234)
);

HB1xp67_ASAP7_75t_L g6235 ( 
.A(n_6036),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_6038),
.Y(n_6236)
);

NAND2xp5_ASAP7_75t_L g6237 ( 
.A(n_6154),
.B(n_4990),
.Y(n_6237)
);

INVx2_ASAP7_75t_L g6238 ( 
.A(n_6085),
.Y(n_6238)
);

OR2x2_ASAP7_75t_L g6239 ( 
.A(n_6173),
.B(n_488),
.Y(n_6239)
);

INVx1_ASAP7_75t_L g6240 ( 
.A(n_6081),
.Y(n_6240)
);

BUFx6f_ASAP7_75t_L g6241 ( 
.A(n_6069),
.Y(n_6241)
);

INVx3_ASAP7_75t_L g6242 ( 
.A(n_6069),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_6082),
.Y(n_6243)
);

HB1xp67_ASAP7_75t_L g6244 ( 
.A(n_6025),
.Y(n_6244)
);

INVxp67_ASAP7_75t_L g6245 ( 
.A(n_6149),
.Y(n_6245)
);

OR2x2_ASAP7_75t_L g6246 ( 
.A(n_6176),
.B(n_488),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_6034),
.Y(n_6247)
);

AND2x2_ASAP7_75t_L g6248 ( 
.A(n_6128),
.B(n_488),
.Y(n_6248)
);

AO31x2_ASAP7_75t_L g6249 ( 
.A1(n_6163),
.A2(n_6148),
.A3(n_6105),
.B(n_6112),
.Y(n_6249)
);

OR2x2_ASAP7_75t_L g6250 ( 
.A(n_6026),
.B(n_489),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_6165),
.Y(n_6251)
);

AND2x4_ASAP7_75t_SL g6252 ( 
.A(n_6061),
.B(n_489),
.Y(n_6252)
);

NAND2xp33_ASAP7_75t_SL g6253 ( 
.A(n_6060),
.B(n_490),
.Y(n_6253)
);

INVx1_ASAP7_75t_L g6254 ( 
.A(n_6087),
.Y(n_6254)
);

AND2x4_ASAP7_75t_L g6255 ( 
.A(n_6056),
.B(n_490),
.Y(n_6255)
);

NAND2xp5_ASAP7_75t_L g6256 ( 
.A(n_6126),
.B(n_4992),
.Y(n_6256)
);

BUFx3_ASAP7_75t_L g6257 ( 
.A(n_6069),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6127),
.B(n_491),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_6077),
.Y(n_6259)
);

HB1xp67_ASAP7_75t_L g6260 ( 
.A(n_6088),
.Y(n_6260)
);

HB1xp67_ASAP7_75t_L g6261 ( 
.A(n_6093),
.Y(n_6261)
);

INVx3_ASAP7_75t_L g6262 ( 
.A(n_6132),
.Y(n_6262)
);

AND2x4_ASAP7_75t_L g6263 ( 
.A(n_6031),
.B(n_491),
.Y(n_6263)
);

HB1xp67_ASAP7_75t_L g6264 ( 
.A(n_6107),
.Y(n_6264)
);

INVx2_ASAP7_75t_L g6265 ( 
.A(n_6113),
.Y(n_6265)
);

OR2x2_ASAP7_75t_L g6266 ( 
.A(n_6024),
.B(n_492),
.Y(n_6266)
);

AOI22xp5_ASAP7_75t_L g6267 ( 
.A1(n_6170),
.A2(n_4565),
.B1(n_4995),
.B2(n_4994),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_6160),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_6138),
.Y(n_6269)
);

AND2x4_ASAP7_75t_SL g6270 ( 
.A(n_6134),
.B(n_492),
.Y(n_6270)
);

AND2x2_ASAP7_75t_L g6271 ( 
.A(n_6042),
.B(n_6110),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_6064),
.Y(n_6272)
);

AND2x2_ASAP7_75t_L g6273 ( 
.A(n_6118),
.B(n_492),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_6108),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_6124),
.Y(n_6275)
);

AND2x2_ASAP7_75t_L g6276 ( 
.A(n_6109),
.B(n_493),
.Y(n_6276)
);

AND2x2_ASAP7_75t_L g6277 ( 
.A(n_6145),
.B(n_494),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_6116),
.Y(n_6278)
);

NOR2xp33_ASAP7_75t_L g6279 ( 
.A(n_6130),
.B(n_494),
.Y(n_6279)
);

AND2x2_ASAP7_75t_L g6280 ( 
.A(n_6039),
.B(n_494),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6167),
.Y(n_6281)
);

NAND2xp5_ASAP7_75t_L g6282 ( 
.A(n_6041),
.B(n_6021),
.Y(n_6282)
);

INVx4_ASAP7_75t_L g6283 ( 
.A(n_6141),
.Y(n_6283)
);

BUFx2_ASAP7_75t_L g6284 ( 
.A(n_6105),
.Y(n_6284)
);

AND2x2_ASAP7_75t_L g6285 ( 
.A(n_6098),
.B(n_6101),
.Y(n_6285)
);

AO21x2_ASAP7_75t_L g6286 ( 
.A1(n_6166),
.A2(n_5004),
.B(n_495),
.Y(n_6286)
);

INVx2_ASAP7_75t_L g6287 ( 
.A(n_6121),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_6135),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6016),
.Y(n_6289)
);

INVxp67_ASAP7_75t_SL g6290 ( 
.A(n_6151),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_6079),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_6157),
.Y(n_6292)
);

INVx2_ASAP7_75t_L g6293 ( 
.A(n_6139),
.Y(n_6293)
);

HB1xp67_ASAP7_75t_L g6294 ( 
.A(n_6146),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_6106),
.Y(n_6295)
);

NAND2xp5_ASAP7_75t_L g6296 ( 
.A(n_6089),
.B(n_495),
.Y(n_6296)
);

AND2x2_ASAP7_75t_L g6297 ( 
.A(n_6091),
.B(n_496),
.Y(n_6297)
);

INVx5_ASAP7_75t_L g6298 ( 
.A(n_6089),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6123),
.Y(n_6299)
);

BUFx3_ASAP7_75t_L g6300 ( 
.A(n_6136),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_6133),
.Y(n_6301)
);

AND2x4_ASAP7_75t_L g6302 ( 
.A(n_6076),
.B(n_496),
.Y(n_6302)
);

NAND2xp5_ASAP7_75t_L g6303 ( 
.A(n_6084),
.B(n_497),
.Y(n_6303)
);

INVx2_ASAP7_75t_L g6304 ( 
.A(n_6150),
.Y(n_6304)
);

AND2x2_ASAP7_75t_L g6305 ( 
.A(n_6094),
.B(n_497),
.Y(n_6305)
);

NAND2xp5_ASAP7_75t_SL g6306 ( 
.A(n_6112),
.B(n_498),
.Y(n_6306)
);

BUFx2_ASAP7_75t_L g6307 ( 
.A(n_6169),
.Y(n_6307)
);

INVx2_ASAP7_75t_L g6308 ( 
.A(n_6067),
.Y(n_6308)
);

AND2x2_ASAP7_75t_L g6309 ( 
.A(n_6096),
.B(n_498),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_6137),
.Y(n_6310)
);

OR2x2_ASAP7_75t_L g6311 ( 
.A(n_6075),
.B(n_498),
.Y(n_6311)
);

OR2x2_ASAP7_75t_SL g6312 ( 
.A(n_6129),
.B(n_499),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_6049),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_6050),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_6078),
.Y(n_6315)
);

AND2x4_ASAP7_75t_SL g6316 ( 
.A(n_6147),
.B(n_6103),
.Y(n_6316)
);

INVx3_ASAP7_75t_L g6317 ( 
.A(n_6161),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6066),
.Y(n_6318)
);

OR2x2_ASAP7_75t_L g6319 ( 
.A(n_6153),
.B(n_500),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_6115),
.B(n_500),
.Y(n_6320)
);

OR2x2_ASAP7_75t_L g6321 ( 
.A(n_6179),
.B(n_6117),
.Y(n_6321)
);

INVx1_ASAP7_75t_SL g6322 ( 
.A(n_6193),
.Y(n_6322)
);

OAI21xp33_ASAP7_75t_L g6323 ( 
.A1(n_6189),
.A2(n_6054),
.B(n_6119),
.Y(n_6323)
);

INVx1_ASAP7_75t_L g6324 ( 
.A(n_6307),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6307),
.Y(n_6325)
);

NAND2xp5_ASAP7_75t_L g6326 ( 
.A(n_6227),
.B(n_6072),
.Y(n_6326)
);

NAND2xp5_ASAP7_75t_L g6327 ( 
.A(n_6298),
.B(n_6080),
.Y(n_6327)
);

INVxp67_ASAP7_75t_L g6328 ( 
.A(n_6185),
.Y(n_6328)
);

OAI21xp5_ASAP7_75t_SL g6329 ( 
.A1(n_6181),
.A2(n_6063),
.B(n_6052),
.Y(n_6329)
);

INVxp67_ASAP7_75t_SL g6330 ( 
.A(n_6279),
.Y(n_6330)
);

NAND2xp5_ASAP7_75t_L g6331 ( 
.A(n_6298),
.B(n_6090),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_6223),
.Y(n_6332)
);

INVx2_ASAP7_75t_L g6333 ( 
.A(n_6200),
.Y(n_6333)
);

HB1xp67_ASAP7_75t_L g6334 ( 
.A(n_6178),
.Y(n_6334)
);

INVx2_ASAP7_75t_L g6335 ( 
.A(n_6200),
.Y(n_6335)
);

NOR2xp33_ASAP7_75t_L g6336 ( 
.A(n_6187),
.B(n_6148),
.Y(n_6336)
);

HB1xp67_ASAP7_75t_L g6337 ( 
.A(n_6206),
.Y(n_6337)
);

AOI211x1_ASAP7_75t_SL g6338 ( 
.A1(n_6199),
.A2(n_6168),
.B(n_6070),
.C(n_6054),
.Y(n_6338)
);

INVx2_ASAP7_75t_SL g6339 ( 
.A(n_6181),
.Y(n_6339)
);

INVx2_ASAP7_75t_L g6340 ( 
.A(n_6192),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6230),
.Y(n_6341)
);

OR2x2_ASAP7_75t_L g6342 ( 
.A(n_6195),
.B(n_6164),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_6233),
.Y(n_6343)
);

HB1xp67_ASAP7_75t_L g6344 ( 
.A(n_6202),
.Y(n_6344)
);

BUFx2_ASAP7_75t_L g6345 ( 
.A(n_6184),
.Y(n_6345)
);

INVx2_ASAP7_75t_SL g6346 ( 
.A(n_6209),
.Y(n_6346)
);

INVx1_ASAP7_75t_L g6347 ( 
.A(n_6217),
.Y(n_6347)
);

NAND2xp5_ASAP7_75t_L g6348 ( 
.A(n_6298),
.B(n_6290),
.Y(n_6348)
);

INVx1_ASAP7_75t_L g6349 ( 
.A(n_6198),
.Y(n_6349)
);

AO21x2_ASAP7_75t_L g6350 ( 
.A1(n_6196),
.A2(n_6097),
.B(n_6095),
.Y(n_6350)
);

BUFx3_ASAP7_75t_L g6351 ( 
.A(n_6216),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_6203),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_6192),
.Y(n_6353)
);

AOI21x1_ASAP7_75t_L g6354 ( 
.A1(n_6284),
.A2(n_6060),
.B(n_6070),
.Y(n_6354)
);

NAND2xp5_ASAP7_75t_L g6355 ( 
.A(n_6276),
.B(n_6104),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_6228),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_6216),
.Y(n_6357)
);

BUFx6f_ASAP7_75t_L g6358 ( 
.A(n_6241),
.Y(n_6358)
);

INVx2_ASAP7_75t_L g6359 ( 
.A(n_6255),
.Y(n_6359)
);

INVx1_ASAP7_75t_L g6360 ( 
.A(n_6207),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_6255),
.Y(n_6361)
);

A2O1A1Ixp33_ASAP7_75t_L g6362 ( 
.A1(n_6263),
.A2(n_6114),
.B(n_6122),
.C(n_6120),
.Y(n_6362)
);

OR2x2_ASAP7_75t_L g6363 ( 
.A(n_6183),
.B(n_6125),
.Y(n_6363)
);

HB1xp67_ASAP7_75t_L g6364 ( 
.A(n_6188),
.Y(n_6364)
);

INVx2_ASAP7_75t_L g6365 ( 
.A(n_6186),
.Y(n_6365)
);

INVx2_ASAP7_75t_L g6366 ( 
.A(n_6190),
.Y(n_6366)
);

INVx1_ASAP7_75t_SL g6367 ( 
.A(n_6221),
.Y(n_6367)
);

NAND2xp5_ASAP7_75t_L g6368 ( 
.A(n_6320),
.B(n_6131),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_6210),
.Y(n_6369)
);

INVxp67_ASAP7_75t_L g6370 ( 
.A(n_6229),
.Y(n_6370)
);

INVx2_ASAP7_75t_L g6371 ( 
.A(n_6214),
.Y(n_6371)
);

A2O1A1Ixp33_ASAP7_75t_L g6372 ( 
.A1(n_6263),
.A2(n_6144),
.B(n_6159),
.C(n_6111),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_6254),
.B(n_6142),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_6277),
.Y(n_6374)
);

NAND2xp5_ASAP7_75t_L g6375 ( 
.A(n_6271),
.B(n_6156),
.Y(n_6375)
);

OA21x2_ASAP7_75t_L g6376 ( 
.A1(n_6284),
.A2(n_6156),
.B(n_500),
.Y(n_6376)
);

CKINVDCx20_ASAP7_75t_R g6377 ( 
.A(n_6312),
.Y(n_6377)
);

AND2x2_ASAP7_75t_L g6378 ( 
.A(n_6285),
.B(n_501),
.Y(n_6378)
);

A2O1A1Ixp33_ASAP7_75t_L g6379 ( 
.A1(n_6253),
.A2(n_503),
.B(n_501),
.C(n_502),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_6248),
.Y(n_6380)
);

NOR2xp33_ASAP7_75t_L g6381 ( 
.A(n_6204),
.B(n_502),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6211),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_6222),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_6226),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6188),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_6249),
.Y(n_6386)
);

OR2x2_ASAP7_75t_L g6387 ( 
.A(n_6191),
.B(n_502),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_6249),
.Y(n_6388)
);

OA21x2_ASAP7_75t_L g6389 ( 
.A1(n_6205),
.A2(n_503),
.B(n_504),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_6252),
.B(n_504),
.Y(n_6390)
);

OAI21x1_ASAP7_75t_L g6391 ( 
.A1(n_6242),
.A2(n_504),
.B(n_505),
.Y(n_6391)
);

BUFx12f_ASAP7_75t_L g6392 ( 
.A(n_6283),
.Y(n_6392)
);

INVx2_ASAP7_75t_L g6393 ( 
.A(n_6180),
.Y(n_6393)
);

INVx1_ASAP7_75t_L g6394 ( 
.A(n_6194),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_6235),
.Y(n_6395)
);

INVx2_ASAP7_75t_SL g6396 ( 
.A(n_6257),
.Y(n_6396)
);

BUFx3_ASAP7_75t_L g6397 ( 
.A(n_6241),
.Y(n_6397)
);

INVx2_ASAP7_75t_L g6398 ( 
.A(n_6201),
.Y(n_6398)
);

AND2x2_ASAP7_75t_L g6399 ( 
.A(n_6273),
.B(n_505),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6260),
.Y(n_6400)
);

NAND3xp33_ASAP7_75t_L g6401 ( 
.A(n_6292),
.B(n_506),
.C(n_507),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_6261),
.Y(n_6402)
);

BUFx2_ASAP7_75t_L g6403 ( 
.A(n_6300),
.Y(n_6403)
);

OR2x6_ASAP7_75t_L g6404 ( 
.A(n_6296),
.B(n_506),
.Y(n_6404)
);

CKINVDCx20_ASAP7_75t_R g6405 ( 
.A(n_6270),
.Y(n_6405)
);

BUFx3_ASAP7_75t_L g6406 ( 
.A(n_6302),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_6264),
.Y(n_6407)
);

BUFx2_ASAP7_75t_L g6408 ( 
.A(n_6294),
.Y(n_6408)
);

OAI21xp33_ASAP7_75t_L g6409 ( 
.A1(n_6259),
.A2(n_506),
.B(n_507),
.Y(n_6409)
);

INVx2_ASAP7_75t_L g6410 ( 
.A(n_6234),
.Y(n_6410)
);

INVx2_ASAP7_75t_L g6411 ( 
.A(n_6238),
.Y(n_6411)
);

CKINVDCx20_ASAP7_75t_R g6412 ( 
.A(n_6258),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_6265),
.Y(n_6413)
);

INVx2_ASAP7_75t_L g6414 ( 
.A(n_6278),
.Y(n_6414)
);

HB1xp67_ASAP7_75t_L g6415 ( 
.A(n_6232),
.Y(n_6415)
);

AND2x2_ASAP7_75t_L g6416 ( 
.A(n_6297),
.B(n_507),
.Y(n_6416)
);

BUFx3_ASAP7_75t_L g6417 ( 
.A(n_6302),
.Y(n_6417)
);

NAND2xp5_ASAP7_75t_L g6418 ( 
.A(n_6245),
.B(n_508),
.Y(n_6418)
);

HB1xp67_ASAP7_75t_L g6419 ( 
.A(n_6244),
.Y(n_6419)
);

NAND4xp25_ASAP7_75t_L g6420 ( 
.A(n_6251),
.B(n_510),
.C(n_508),
.D(n_509),
.Y(n_6420)
);

OAI211xp5_ASAP7_75t_L g6421 ( 
.A1(n_6182),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_6421)
);

OA21x2_ASAP7_75t_L g6422 ( 
.A1(n_6306),
.A2(n_511),
.B(n_512),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_6274),
.Y(n_6423)
);

INVx2_ASAP7_75t_SL g6424 ( 
.A(n_6316),
.Y(n_6424)
);

AOI21xp33_ASAP7_75t_L g6425 ( 
.A1(n_6299),
.A2(n_511),
.B(n_512),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6275),
.Y(n_6426)
);

INVx2_ASAP7_75t_L g6427 ( 
.A(n_6287),
.Y(n_6427)
);

OAI21xp33_ASAP7_75t_L g6428 ( 
.A1(n_6288),
.A2(n_512),
.B(n_513),
.Y(n_6428)
);

INVx4_ASAP7_75t_L g6429 ( 
.A(n_6262),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_6319),
.Y(n_6430)
);

INVx2_ASAP7_75t_L g6431 ( 
.A(n_6293),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6224),
.Y(n_6432)
);

HB1xp67_ASAP7_75t_L g6433 ( 
.A(n_6304),
.Y(n_6433)
);

NOR2xp33_ASAP7_75t_L g6434 ( 
.A(n_6281),
.B(n_513),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_6315),
.Y(n_6435)
);

INVx8_ASAP7_75t_L g6436 ( 
.A(n_6219),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_6215),
.Y(n_6437)
);

HB1xp67_ASAP7_75t_L g6438 ( 
.A(n_6220),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6197),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6317),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6225),
.Y(n_6441)
);

NOR2xp67_ASAP7_75t_L g6442 ( 
.A(n_6218),
.B(n_513),
.Y(n_6442)
);

AOI21xp5_ASAP7_75t_L g6443 ( 
.A1(n_6212),
.A2(n_514),
.B(n_515),
.Y(n_6443)
);

BUFx3_ASAP7_75t_L g6444 ( 
.A(n_6236),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_6308),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6303),
.Y(n_6446)
);

OR2x6_ASAP7_75t_SL g6447 ( 
.A(n_6239),
.B(n_6246),
.Y(n_6447)
);

AND2x2_ASAP7_75t_L g6448 ( 
.A(n_6305),
.B(n_514),
.Y(n_6448)
);

NOR3xp33_ASAP7_75t_L g6449 ( 
.A(n_6212),
.B(n_515),
.C(n_516),
.Y(n_6449)
);

INVx2_ASAP7_75t_L g6450 ( 
.A(n_6213),
.Y(n_6450)
);

INVx2_ASAP7_75t_L g6451 ( 
.A(n_6208),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_6280),
.Y(n_6452)
);

CKINVDCx20_ASAP7_75t_R g6453 ( 
.A(n_6309),
.Y(n_6453)
);

INVx2_ASAP7_75t_L g6454 ( 
.A(n_6247),
.Y(n_6454)
);

NAND2xp5_ASAP7_75t_L g6455 ( 
.A(n_6268),
.B(n_515),
.Y(n_6455)
);

AOI21xp5_ASAP7_75t_L g6456 ( 
.A1(n_6240),
.A2(n_516),
.B(n_517),
.Y(n_6456)
);

INVx3_ASAP7_75t_L g6457 ( 
.A(n_6243),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6256),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_6289),
.Y(n_6459)
);

AOI21xp5_ASAP7_75t_L g6460 ( 
.A1(n_6266),
.A2(n_516),
.B(n_517),
.Y(n_6460)
);

INVx1_ASAP7_75t_L g6461 ( 
.A(n_6250),
.Y(n_6461)
);

AND2x2_ASAP7_75t_L g6462 ( 
.A(n_6269),
.B(n_517),
.Y(n_6462)
);

INVx2_ASAP7_75t_SL g6463 ( 
.A(n_6311),
.Y(n_6463)
);

AOI21xp5_ASAP7_75t_L g6464 ( 
.A1(n_6295),
.A2(n_518),
.B(n_519),
.Y(n_6464)
);

HB1xp67_ASAP7_75t_L g6465 ( 
.A(n_6291),
.Y(n_6465)
);

OR2x2_ASAP7_75t_L g6466 ( 
.A(n_6282),
.B(n_519),
.Y(n_6466)
);

INVx2_ASAP7_75t_L g6467 ( 
.A(n_6272),
.Y(n_6467)
);

NAND2xp5_ASAP7_75t_L g6468 ( 
.A(n_6286),
.B(n_519),
.Y(n_6468)
);

NAND4xp25_ASAP7_75t_L g6469 ( 
.A(n_6313),
.B(n_522),
.C(n_520),
.D(n_521),
.Y(n_6469)
);

INVx2_ASAP7_75t_L g6470 ( 
.A(n_6314),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_6237),
.Y(n_6471)
);

A2O1A1Ixp33_ASAP7_75t_L g6472 ( 
.A1(n_6318),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_6472)
);

AND2x2_ASAP7_75t_L g6473 ( 
.A(n_6301),
.B(n_520),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_L g6474 ( 
.A(n_6310),
.B(n_521),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_6231),
.B(n_6267),
.Y(n_6475)
);

BUFx6f_ASAP7_75t_L g6476 ( 
.A(n_6241),
.Y(n_6476)
);

OA21x2_ASAP7_75t_L g6477 ( 
.A1(n_6189),
.A2(n_522),
.B(n_523),
.Y(n_6477)
);

INVx4_ASAP7_75t_SL g6478 ( 
.A(n_6216),
.Y(n_6478)
);

HB1xp67_ASAP7_75t_L g6479 ( 
.A(n_6179),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6193),
.Y(n_6480)
);

AND2x2_ASAP7_75t_L g6481 ( 
.A(n_6193),
.B(n_523),
.Y(n_6481)
);

INVx4_ASAP7_75t_L g6482 ( 
.A(n_6187),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6193),
.B(n_523),
.Y(n_6483)
);

NAND2xp5_ASAP7_75t_L g6484 ( 
.A(n_6189),
.B(n_524),
.Y(n_6484)
);

AND2x2_ASAP7_75t_L g6485 ( 
.A(n_6193),
.B(n_524),
.Y(n_6485)
);

NAND2xp5_ASAP7_75t_L g6486 ( 
.A(n_6189),
.B(n_524),
.Y(n_6486)
);

AND2x2_ASAP7_75t_L g6487 ( 
.A(n_6193),
.B(n_525),
.Y(n_6487)
);

OA21x2_ASAP7_75t_L g6488 ( 
.A1(n_6189),
.A2(n_525),
.B(n_526),
.Y(n_6488)
);

INVx3_ASAP7_75t_L g6489 ( 
.A(n_6193),
.Y(n_6489)
);

NAND2xp33_ASAP7_75t_L g6490 ( 
.A(n_6298),
.B(n_525),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6189),
.Y(n_6491)
);

NAND2xp5_ASAP7_75t_L g6492 ( 
.A(n_6189),
.B(n_526),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6189),
.B(n_526),
.Y(n_6493)
);

NAND2xp5_ASAP7_75t_L g6494 ( 
.A(n_6189),
.B(n_527),
.Y(n_6494)
);

INVx1_ASAP7_75t_L g6495 ( 
.A(n_6189),
.Y(n_6495)
);

O2A1O1Ixp33_ASAP7_75t_L g6496 ( 
.A1(n_6189),
.A2(n_529),
.B(n_527),
.C(n_528),
.Y(n_6496)
);

BUFx6f_ASAP7_75t_L g6497 ( 
.A(n_6241),
.Y(n_6497)
);

NAND2xp5_ASAP7_75t_L g6498 ( 
.A(n_6322),
.B(n_527),
.Y(n_6498)
);

OAI211xp5_ASAP7_75t_SL g6499 ( 
.A1(n_6338),
.A2(n_530),
.B(n_528),
.C(n_529),
.Y(n_6499)
);

NOR3xp33_ASAP7_75t_L g6500 ( 
.A(n_6482),
.B(n_531),
.C(n_530),
.Y(n_6500)
);

NAND3xp33_ASAP7_75t_L g6501 ( 
.A(n_6480),
.B(n_528),
.C(n_530),
.Y(n_6501)
);

NAND2xp5_ASAP7_75t_L g6502 ( 
.A(n_6489),
.B(n_531),
.Y(n_6502)
);

AOI22xp5_ASAP7_75t_L g6503 ( 
.A1(n_6392),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_6503)
);

INVxp67_ASAP7_75t_L g6504 ( 
.A(n_6336),
.Y(n_6504)
);

AOI22xp5_ASAP7_75t_L g6505 ( 
.A1(n_6377),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_6505)
);

OR2x2_ASAP7_75t_L g6506 ( 
.A(n_6491),
.B(n_6495),
.Y(n_6506)
);

OR2x2_ASAP7_75t_L g6507 ( 
.A(n_6484),
.B(n_533),
.Y(n_6507)
);

AND2x2_ASAP7_75t_L g6508 ( 
.A(n_6339),
.B(n_534),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_6346),
.B(n_534),
.Y(n_6509)
);

AND2x4_ASAP7_75t_SL g6510 ( 
.A(n_6429),
.B(n_535),
.Y(n_6510)
);

AOI22xp33_ASAP7_75t_L g6511 ( 
.A1(n_6396),
.A2(n_538),
.B1(n_535),
.B2(n_537),
.Y(n_6511)
);

AND2x4_ASAP7_75t_SL g6512 ( 
.A(n_6358),
.B(n_537),
.Y(n_6512)
);

NOR2xp33_ASAP7_75t_L g6513 ( 
.A(n_6329),
.B(n_537),
.Y(n_6513)
);

OR2x2_ASAP7_75t_L g6514 ( 
.A(n_6486),
.B(n_538),
.Y(n_6514)
);

INVx2_ASAP7_75t_L g6515 ( 
.A(n_6340),
.Y(n_6515)
);

AND2x2_ASAP7_75t_L g6516 ( 
.A(n_6424),
.B(n_539),
.Y(n_6516)
);

INVxp33_ASAP7_75t_SL g6517 ( 
.A(n_6481),
.Y(n_6517)
);

AO21x2_ASAP7_75t_L g6518 ( 
.A1(n_6386),
.A2(n_539),
.B(n_540),
.Y(n_6518)
);

AND2x4_ASAP7_75t_L g6519 ( 
.A(n_6478),
.B(n_540),
.Y(n_6519)
);

AND2x2_ASAP7_75t_L g6520 ( 
.A(n_6345),
.B(n_540),
.Y(n_6520)
);

AOI221xp5_ASAP7_75t_L g6521 ( 
.A1(n_6400),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.C(n_544),
.Y(n_6521)
);

AND2x2_ASAP7_75t_L g6522 ( 
.A(n_6403),
.B(n_541),
.Y(n_6522)
);

NAND3xp33_ASAP7_75t_L g6523 ( 
.A(n_6358),
.B(n_542),
.C(n_543),
.Y(n_6523)
);

NOR3xp33_ASAP7_75t_L g6524 ( 
.A(n_6348),
.B(n_545),
.C(n_544),
.Y(n_6524)
);

AND2x2_ASAP7_75t_L g6525 ( 
.A(n_6373),
.B(n_543),
.Y(n_6525)
);

NAND3xp33_ASAP7_75t_L g6526 ( 
.A(n_6476),
.B(n_6497),
.C(n_6325),
.Y(n_6526)
);

NOR3xp33_ASAP7_75t_L g6527 ( 
.A(n_6397),
.B(n_546),
.C(n_545),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_SL g6528 ( 
.A(n_6476),
.B(n_544),
.Y(n_6528)
);

NAND3xp33_ASAP7_75t_L g6529 ( 
.A(n_6497),
.B(n_545),
.C(n_547),
.Y(n_6529)
);

OAI211xp5_ASAP7_75t_SL g6530 ( 
.A1(n_6324),
.A2(n_550),
.B(n_548),
.C(n_549),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6483),
.Y(n_6531)
);

NOR2xp33_ASAP7_75t_L g6532 ( 
.A(n_6353),
.B(n_548),
.Y(n_6532)
);

AND2x2_ASAP7_75t_L g6533 ( 
.A(n_6378),
.B(n_548),
.Y(n_6533)
);

NAND4xp75_ASAP7_75t_L g6534 ( 
.A(n_6402),
.B(n_557),
.C(n_565),
.D(n_549),
.Y(n_6534)
);

NAND3xp33_ASAP7_75t_L g6535 ( 
.A(n_6337),
.B(n_550),
.C(n_551),
.Y(n_6535)
);

AND2x2_ASAP7_75t_L g6536 ( 
.A(n_6485),
.B(n_550),
.Y(n_6536)
);

OR2x2_ASAP7_75t_L g6537 ( 
.A(n_6492),
.B(n_551),
.Y(n_6537)
);

NAND3xp33_ASAP7_75t_L g6538 ( 
.A(n_6479),
.B(n_551),
.C(n_552),
.Y(n_6538)
);

BUFx3_ASAP7_75t_L g6539 ( 
.A(n_6351),
.Y(n_6539)
);

AND2x2_ASAP7_75t_L g6540 ( 
.A(n_6487),
.B(n_552),
.Y(n_6540)
);

OAI221xp5_ASAP7_75t_SL g6541 ( 
.A1(n_6362),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.C(n_556),
.Y(n_6541)
);

NAND3xp33_ASAP7_75t_L g6542 ( 
.A(n_6490),
.B(n_553),
.C(n_554),
.Y(n_6542)
);

AO21x1_ASAP7_75t_SL g6543 ( 
.A1(n_6327),
.A2(n_561),
.B(n_553),
.Y(n_6543)
);

CKINVDCx14_ASAP7_75t_R g6544 ( 
.A(n_6405),
.Y(n_6544)
);

NAND3xp33_ASAP7_75t_L g6545 ( 
.A(n_6364),
.B(n_554),
.C(n_555),
.Y(n_6545)
);

AND2x2_ASAP7_75t_L g6546 ( 
.A(n_6478),
.B(n_555),
.Y(n_6546)
);

BUFx3_ASAP7_75t_L g6547 ( 
.A(n_6357),
.Y(n_6547)
);

AND2x2_ASAP7_75t_L g6548 ( 
.A(n_6359),
.B(n_556),
.Y(n_6548)
);

INVx1_ASAP7_75t_L g6549 ( 
.A(n_6344),
.Y(n_6549)
);

AOI22xp33_ASAP7_75t_L g6550 ( 
.A1(n_6458),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_6550)
);

AND2x2_ASAP7_75t_SL g6551 ( 
.A(n_6449),
.B(n_557),
.Y(n_6551)
);

AOI22xp5_ASAP7_75t_L g6552 ( 
.A1(n_6412),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_6552)
);

OR2x6_ASAP7_75t_L g6553 ( 
.A(n_6361),
.B(n_558),
.Y(n_6553)
);

AO21x2_ASAP7_75t_L g6554 ( 
.A1(n_6388),
.A2(n_559),
.B(n_562),
.Y(n_6554)
);

NAND3xp33_ASAP7_75t_L g6555 ( 
.A(n_6334),
.B(n_562),
.C(n_563),
.Y(n_6555)
);

AOI22xp33_ASAP7_75t_L g6556 ( 
.A1(n_6471),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_6556)
);

OR2x2_ASAP7_75t_L g6557 ( 
.A(n_6493),
.B(n_563),
.Y(n_6557)
);

NOR3xp33_ASAP7_75t_L g6558 ( 
.A(n_6494),
.B(n_566),
.C(n_565),
.Y(n_6558)
);

NOR3xp33_ASAP7_75t_L g6559 ( 
.A(n_6496),
.B(n_566),
.C(n_565),
.Y(n_6559)
);

NAND4xp75_ASAP7_75t_L g6560 ( 
.A(n_6407),
.B(n_573),
.C(n_581),
.D(n_564),
.Y(n_6560)
);

AND2x2_ASAP7_75t_L g6561 ( 
.A(n_6462),
.B(n_564),
.Y(n_6561)
);

OR2x2_ASAP7_75t_L g6562 ( 
.A(n_6365),
.B(n_566),
.Y(n_6562)
);

OR2x2_ASAP7_75t_L g6563 ( 
.A(n_6387),
.B(n_567),
.Y(n_6563)
);

INVx1_ASAP7_75t_L g6564 ( 
.A(n_6408),
.Y(n_6564)
);

NOR3xp33_ASAP7_75t_L g6565 ( 
.A(n_6330),
.B(n_570),
.C(n_569),
.Y(n_6565)
);

INVx2_ASAP7_75t_L g6566 ( 
.A(n_6406),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_L g6567 ( 
.A(n_6381),
.B(n_568),
.Y(n_6567)
);

NOR3xp33_ASAP7_75t_L g6568 ( 
.A(n_6401),
.B(n_571),
.C(n_569),
.Y(n_6568)
);

AND2x4_ASAP7_75t_L g6569 ( 
.A(n_6333),
.B(n_568),
.Y(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_6433),
.B(n_568),
.Y(n_6570)
);

AND2x2_ASAP7_75t_L g6571 ( 
.A(n_6417),
.B(n_569),
.Y(n_6571)
);

BUFx2_ASAP7_75t_L g6572 ( 
.A(n_6360),
.Y(n_6572)
);

NAND3xp33_ASAP7_75t_L g6573 ( 
.A(n_6385),
.B(n_571),
.C(n_572),
.Y(n_6573)
);

INVxp67_ASAP7_75t_SL g6574 ( 
.A(n_6418),
.Y(n_6574)
);

NOR2xp33_ASAP7_75t_L g6575 ( 
.A(n_6367),
.B(n_572),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6335),
.B(n_573),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_6328),
.B(n_573),
.Y(n_6577)
);

NAND2xp5_ASAP7_75t_SL g6578 ( 
.A(n_6369),
.B(n_6371),
.Y(n_6578)
);

NAND3xp33_ASAP7_75t_L g6579 ( 
.A(n_6488),
.B(n_574),
.C(n_575),
.Y(n_6579)
);

INVx2_ASAP7_75t_L g6580 ( 
.A(n_6383),
.Y(n_6580)
);

AOI22xp33_ASAP7_75t_L g6581 ( 
.A1(n_6440),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_6581)
);

AOI22xp33_ASAP7_75t_L g6582 ( 
.A1(n_6445),
.A2(n_577),
.B1(n_574),
.B2(n_576),
.Y(n_6582)
);

OAI21xp5_ASAP7_75t_L g6583 ( 
.A1(n_6443),
.A2(n_577),
.B(n_578),
.Y(n_6583)
);

AND2x2_ASAP7_75t_L g6584 ( 
.A(n_6366),
.B(n_577),
.Y(n_6584)
);

NOR3xp33_ASAP7_75t_L g6585 ( 
.A(n_6421),
.B(n_580),
.C(n_579),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_6415),
.Y(n_6586)
);

AND2x2_ASAP7_75t_L g6587 ( 
.A(n_6473),
.B(n_578),
.Y(n_6587)
);

AND2x2_ASAP7_75t_L g6588 ( 
.A(n_6432),
.B(n_579),
.Y(n_6588)
);

OR2x2_ASAP7_75t_L g6589 ( 
.A(n_6468),
.B(n_579),
.Y(n_6589)
);

AOI22xp33_ASAP7_75t_L g6590 ( 
.A1(n_6430),
.A2(n_582),
.B1(n_580),
.B2(n_581),
.Y(n_6590)
);

AOI211xp5_ASAP7_75t_L g6591 ( 
.A1(n_6382),
.A2(n_583),
.B(n_581),
.C(n_582),
.Y(n_6591)
);

OR2x2_ASAP7_75t_L g6592 ( 
.A(n_6410),
.B(n_583),
.Y(n_6592)
);

AND2x4_ASAP7_75t_L g6593 ( 
.A(n_6444),
.B(n_583),
.Y(n_6593)
);

BUFx2_ASAP7_75t_L g6594 ( 
.A(n_6384),
.Y(n_6594)
);

NOR2x1_ASAP7_75t_SL g6595 ( 
.A(n_6331),
.B(n_584),
.Y(n_6595)
);

NAND2xp5_ASAP7_75t_L g6596 ( 
.A(n_6442),
.B(n_584),
.Y(n_6596)
);

AND2x2_ASAP7_75t_L g6597 ( 
.A(n_6347),
.B(n_584),
.Y(n_6597)
);

NAND2xp5_ASAP7_75t_L g6598 ( 
.A(n_6411),
.B(n_585),
.Y(n_6598)
);

NAND3xp33_ASAP7_75t_L g6599 ( 
.A(n_6488),
.B(n_585),
.C(n_586),
.Y(n_6599)
);

AND2x4_ASAP7_75t_L g6600 ( 
.A(n_6413),
.B(n_6414),
.Y(n_6600)
);

AND2x2_ASAP7_75t_L g6601 ( 
.A(n_6394),
.B(n_585),
.Y(n_6601)
);

AND2x2_ASAP7_75t_L g6602 ( 
.A(n_6341),
.B(n_6343),
.Y(n_6602)
);

AOI22xp5_ASAP7_75t_L g6603 ( 
.A1(n_6453),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_6603)
);

AND2x2_ASAP7_75t_L g6604 ( 
.A(n_6370),
.B(n_586),
.Y(n_6604)
);

INVx2_ASAP7_75t_L g6605 ( 
.A(n_6427),
.Y(n_6605)
);

INVx3_ASAP7_75t_L g6606 ( 
.A(n_6431),
.Y(n_6606)
);

NAND2xp5_ASAP7_75t_L g6607 ( 
.A(n_6435),
.B(n_587),
.Y(n_6607)
);

AOI22xp33_ASAP7_75t_L g6608 ( 
.A1(n_6439),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_6608)
);

AND2x2_ASAP7_75t_L g6609 ( 
.A(n_6356),
.B(n_6380),
.Y(n_6609)
);

NAND3xp33_ASAP7_75t_L g6610 ( 
.A(n_6477),
.B(n_588),
.C(n_589),
.Y(n_6610)
);

AND4x1_ASAP7_75t_L g6611 ( 
.A(n_6434),
.B(n_591),
.C(n_589),
.D(n_590),
.Y(n_6611)
);

NOR3xp33_ASAP7_75t_L g6612 ( 
.A(n_6428),
.B(n_590),
.C(n_591),
.Y(n_6612)
);

HB1xp67_ASAP7_75t_L g6613 ( 
.A(n_6419),
.Y(n_6613)
);

AND2x2_ASAP7_75t_L g6614 ( 
.A(n_6332),
.B(n_591),
.Y(n_6614)
);

OR2x2_ASAP7_75t_L g6615 ( 
.A(n_6395),
.B(n_592),
.Y(n_6615)
);

OA211x2_ASAP7_75t_L g6616 ( 
.A1(n_6475),
.A2(n_594),
.B(n_592),
.C(n_593),
.Y(n_6616)
);

NOR2x1_ASAP7_75t_L g6617 ( 
.A(n_6389),
.B(n_592),
.Y(n_6617)
);

AOI211xp5_ASAP7_75t_L g6618 ( 
.A1(n_6372),
.A2(n_595),
.B(n_593),
.C(n_594),
.Y(n_6618)
);

NOR3xp33_ASAP7_75t_L g6619 ( 
.A(n_6425),
.B(n_593),
.C(n_594),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6389),
.Y(n_6620)
);

NAND3xp33_ASAP7_75t_SL g6621 ( 
.A(n_6323),
.B(n_595),
.C(n_596),
.Y(n_6621)
);

AO21x2_ASAP7_75t_L g6622 ( 
.A1(n_6354),
.A2(n_595),
.B(n_596),
.Y(n_6622)
);

NAND3xp33_ASAP7_75t_L g6623 ( 
.A(n_6423),
.B(n_596),
.C(n_597),
.Y(n_6623)
);

NAND4xp75_ASAP7_75t_L g6624 ( 
.A(n_6426),
.B(n_599),
.C(n_597),
.D(n_598),
.Y(n_6624)
);

AOI22xp5_ASAP7_75t_L g6625 ( 
.A1(n_6463),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_6363),
.Y(n_6626)
);

NAND3xp33_ASAP7_75t_L g6627 ( 
.A(n_6393),
.B(n_598),
.C(n_599),
.Y(n_6627)
);

OR2x2_ASAP7_75t_L g6628 ( 
.A(n_6466),
.B(n_600),
.Y(n_6628)
);

AND2x2_ASAP7_75t_L g6629 ( 
.A(n_6452),
.B(n_600),
.Y(n_6629)
);

NAND3xp33_ASAP7_75t_L g6630 ( 
.A(n_6472),
.B(n_601),
.C(n_602),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_SL g6631 ( 
.A(n_6398),
.B(n_601),
.Y(n_6631)
);

NOR2xp33_ASAP7_75t_L g6632 ( 
.A(n_6436),
.B(n_602),
.Y(n_6632)
);

NOR3xp33_ASAP7_75t_SL g6633 ( 
.A(n_6420),
.B(n_603),
.C(n_604),
.Y(n_6633)
);

OR2x2_ASAP7_75t_L g6634 ( 
.A(n_6326),
.B(n_604),
.Y(n_6634)
);

NOR3xp33_ASAP7_75t_L g6635 ( 
.A(n_6409),
.B(n_6469),
.C(n_6474),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6391),
.Y(n_6636)
);

AND2x2_ASAP7_75t_L g6637 ( 
.A(n_6349),
.B(n_604),
.Y(n_6637)
);

AND2x2_ASAP7_75t_L g6638 ( 
.A(n_6352),
.B(n_605),
.Y(n_6638)
);

OR2x2_ASAP7_75t_L g6639 ( 
.A(n_6374),
.B(n_605),
.Y(n_6639)
);

NAND2xp5_ASAP7_75t_L g6640 ( 
.A(n_6460),
.B(n_605),
.Y(n_6640)
);

AND2x2_ASAP7_75t_L g6641 ( 
.A(n_6404),
.B(n_606),
.Y(n_6641)
);

NAND3xp33_ASAP7_75t_L g6642 ( 
.A(n_6437),
.B(n_606),
.C(n_607),
.Y(n_6642)
);

INVx4_ASAP7_75t_L g6643 ( 
.A(n_6539),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_6516),
.Y(n_6644)
);

AND2x2_ASAP7_75t_L g6645 ( 
.A(n_6544),
.B(n_6461),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6522),
.Y(n_6646)
);

NOR3xp33_ASAP7_75t_L g6647 ( 
.A(n_6526),
.B(n_6379),
.C(n_6464),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_6508),
.Y(n_6648)
);

INVx4_ASAP7_75t_L g6649 ( 
.A(n_6519),
.Y(n_6649)
);

AOI21xp5_ASAP7_75t_L g6650 ( 
.A1(n_6620),
.A2(n_6455),
.B(n_6456),
.Y(n_6650)
);

AND2x2_ASAP7_75t_L g6651 ( 
.A(n_6509),
.B(n_6404),
.Y(n_6651)
);

HB1xp67_ASAP7_75t_L g6652 ( 
.A(n_6547),
.Y(n_6652)
);

BUFx12f_ASAP7_75t_L g6653 ( 
.A(n_6519),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6520),
.Y(n_6654)
);

AND2x2_ASAP7_75t_L g6655 ( 
.A(n_6525),
.B(n_6454),
.Y(n_6655)
);

INVx2_ASAP7_75t_L g6656 ( 
.A(n_6566),
.Y(n_6656)
);

AND2x2_ASAP7_75t_L g6657 ( 
.A(n_6571),
.B(n_6467),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6546),
.Y(n_6658)
);

BUFx2_ASAP7_75t_L g6659 ( 
.A(n_6553),
.Y(n_6659)
);

AND2x2_ASAP7_75t_L g6660 ( 
.A(n_6548),
.B(n_6446),
.Y(n_6660)
);

OAI211xp5_ASAP7_75t_L g6661 ( 
.A1(n_6504),
.A2(n_6465),
.B(n_6321),
.C(n_6459),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_6502),
.Y(n_6662)
);

AND2x2_ASAP7_75t_L g6663 ( 
.A(n_6576),
.B(n_6399),
.Y(n_6663)
);

INVx2_ASAP7_75t_SL g6664 ( 
.A(n_6512),
.Y(n_6664)
);

AND2x2_ASAP7_75t_L g6665 ( 
.A(n_6604),
.B(n_6416),
.Y(n_6665)
);

INVx2_ASAP7_75t_L g6666 ( 
.A(n_6600),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_6498),
.Y(n_6667)
);

OAI21xp5_ASAP7_75t_L g6668 ( 
.A1(n_6499),
.A2(n_6438),
.B(n_6451),
.Y(n_6668)
);

INVx2_ASAP7_75t_L g6669 ( 
.A(n_6600),
.Y(n_6669)
);

AND2x2_ASAP7_75t_L g6670 ( 
.A(n_6588),
.B(n_6601),
.Y(n_6670)
);

OAI211xp5_ASAP7_75t_L g6671 ( 
.A1(n_6564),
.A2(n_6441),
.B(n_6457),
.C(n_6470),
.Y(n_6671)
);

AO31x2_ASAP7_75t_L g6672 ( 
.A1(n_6513),
.A2(n_6450),
.A3(n_6355),
.B(n_6368),
.Y(n_6672)
);

INVxp67_ASAP7_75t_SL g6673 ( 
.A(n_6570),
.Y(n_6673)
);

AOI32xp33_ASAP7_75t_L g6674 ( 
.A1(n_6618),
.A2(n_6375),
.A3(n_6390),
.B1(n_6448),
.B2(n_6342),
.Y(n_6674)
);

AOI22xp5_ASAP7_75t_L g6675 ( 
.A1(n_6517),
.A2(n_6436),
.B1(n_6422),
.B2(n_6350),
.Y(n_6675)
);

AND2x2_ASAP7_75t_L g6676 ( 
.A(n_6629),
.B(n_6447),
.Y(n_6676)
);

AND2x2_ASAP7_75t_L g6677 ( 
.A(n_6597),
.B(n_6637),
.Y(n_6677)
);

AND2x2_ASAP7_75t_L g6678 ( 
.A(n_6638),
.B(n_6376),
.Y(n_6678)
);

AND2x2_ASAP7_75t_L g6679 ( 
.A(n_6614),
.B(n_6584),
.Y(n_6679)
);

NAND3xp33_ASAP7_75t_L g6680 ( 
.A(n_6565),
.B(n_6376),
.C(n_607),
.Y(n_6680)
);

AND2x2_ASAP7_75t_L g6681 ( 
.A(n_6577),
.B(n_6543),
.Y(n_6681)
);

AND2x2_ASAP7_75t_L g6682 ( 
.A(n_6595),
.B(n_607),
.Y(n_6682)
);

INVx2_ASAP7_75t_L g6683 ( 
.A(n_6606),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6641),
.Y(n_6684)
);

NAND2xp5_ASAP7_75t_L g6685 ( 
.A(n_6510),
.B(n_608),
.Y(n_6685)
);

OAI22xp5_ASAP7_75t_L g6686 ( 
.A1(n_6506),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_6686)
);

NAND3xp33_ASAP7_75t_L g6687 ( 
.A(n_6579),
.B(n_608),
.C(n_609),
.Y(n_6687)
);

AND2x2_ASAP7_75t_L g6688 ( 
.A(n_6632),
.B(n_609),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6536),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6540),
.Y(n_6690)
);

CKINVDCx16_ASAP7_75t_R g6691 ( 
.A(n_6628),
.Y(n_6691)
);

HB1xp67_ASAP7_75t_L g6692 ( 
.A(n_6515),
.Y(n_6692)
);

INVx1_ASAP7_75t_SL g6693 ( 
.A(n_6594),
.Y(n_6693)
);

INVx2_ASAP7_75t_SL g6694 ( 
.A(n_6580),
.Y(n_6694)
);

OR2x2_ASAP7_75t_L g6695 ( 
.A(n_6553),
.B(n_610),
.Y(n_6695)
);

NOR2xp33_ASAP7_75t_L g6696 ( 
.A(n_6541),
.B(n_610),
.Y(n_6696)
);

HB1xp67_ASAP7_75t_L g6697 ( 
.A(n_6613),
.Y(n_6697)
);

INVx2_ASAP7_75t_SL g6698 ( 
.A(n_6605),
.Y(n_6698)
);

AND2x2_ASAP7_75t_L g6699 ( 
.A(n_6531),
.B(n_611),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6569),
.Y(n_6700)
);

INVx2_ASAP7_75t_SL g6701 ( 
.A(n_6569),
.Y(n_6701)
);

BUFx3_ASAP7_75t_L g6702 ( 
.A(n_6549),
.Y(n_6702)
);

AND2x2_ASAP7_75t_L g6703 ( 
.A(n_6533),
.B(n_6587),
.Y(n_6703)
);

AOI221xp5_ASAP7_75t_L g6704 ( 
.A1(n_6578),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.C(n_614),
.Y(n_6704)
);

INVx2_ASAP7_75t_SL g6705 ( 
.A(n_6593),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6572),
.Y(n_6706)
);

INVx2_ASAP7_75t_L g6707 ( 
.A(n_6593),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_6561),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6598),
.Y(n_6709)
);

NAND2xp5_ASAP7_75t_L g6710 ( 
.A(n_6622),
.B(n_611),
.Y(n_6710)
);

AND2x4_ASAP7_75t_L g6711 ( 
.A(n_6626),
.B(n_612),
.Y(n_6711)
);

INVx2_ASAP7_75t_L g6712 ( 
.A(n_6562),
.Y(n_6712)
);

NOR2x1_ASAP7_75t_L g6713 ( 
.A(n_6599),
.B(n_612),
.Y(n_6713)
);

OR2x2_ASAP7_75t_L g6714 ( 
.A(n_6563),
.B(n_613),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_6607),
.Y(n_6715)
);

INVx2_ASAP7_75t_L g6716 ( 
.A(n_6592),
.Y(n_6716)
);

NAND3xp33_ASAP7_75t_L g6717 ( 
.A(n_6610),
.B(n_613),
.C(n_614),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6636),
.Y(n_6718)
);

HB1xp67_ASAP7_75t_L g6719 ( 
.A(n_6586),
.Y(n_6719)
);

INVx2_ASAP7_75t_L g6720 ( 
.A(n_6534),
.Y(n_6720)
);

AOI22xp33_ASAP7_75t_SL g6721 ( 
.A1(n_6609),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_6721)
);

INVx1_ASAP7_75t_SL g6722 ( 
.A(n_6615),
.Y(n_6722)
);

OR2x2_ASAP7_75t_L g6723 ( 
.A(n_6589),
.B(n_615),
.Y(n_6723)
);

OAI33xp33_ASAP7_75t_L g6724 ( 
.A1(n_6631),
.A2(n_618),
.A3(n_620),
.B1(n_616),
.B2(n_617),
.B3(n_619),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_6617),
.Y(n_6725)
);

NAND3xp33_ASAP7_75t_L g6726 ( 
.A(n_6500),
.B(n_616),
.C(n_618),
.Y(n_6726)
);

BUFx3_ASAP7_75t_L g6727 ( 
.A(n_6567),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_6560),
.Y(n_6728)
);

INVx2_ASAP7_75t_L g6729 ( 
.A(n_6624),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_6518),
.Y(n_6730)
);

NAND2xp5_ASAP7_75t_L g6731 ( 
.A(n_6585),
.B(n_618),
.Y(n_6731)
);

INVx2_ASAP7_75t_SL g6732 ( 
.A(n_6507),
.Y(n_6732)
);

NAND2xp5_ASAP7_75t_L g6733 ( 
.A(n_6633),
.B(n_6527),
.Y(n_6733)
);

AND2x4_ASAP7_75t_SL g6734 ( 
.A(n_6635),
.B(n_619),
.Y(n_6734)
);

AND2x2_ASAP7_75t_L g6735 ( 
.A(n_6602),
.B(n_620),
.Y(n_6735)
);

NOR2xp33_ASAP7_75t_L g6736 ( 
.A(n_6621),
.B(n_621),
.Y(n_6736)
);

AOI22xp33_ASAP7_75t_SL g6737 ( 
.A1(n_6574),
.A2(n_623),
.B1(n_621),
.B2(n_622),
.Y(n_6737)
);

OR2x2_ASAP7_75t_L g6738 ( 
.A(n_6501),
.B(n_621),
.Y(n_6738)
);

NAND2xp5_ASAP7_75t_L g6739 ( 
.A(n_6524),
.B(n_622),
.Y(n_6739)
);

OR2x2_ASAP7_75t_L g6740 ( 
.A(n_6639),
.B(n_623),
.Y(n_6740)
);

INVxp67_ASAP7_75t_L g6741 ( 
.A(n_6575),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_6554),
.Y(n_6742)
);

AOI221xp5_ASAP7_75t_L g6743 ( 
.A1(n_6559),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.C(n_627),
.Y(n_6743)
);

AOI22xp33_ASAP7_75t_L g6744 ( 
.A1(n_6619),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_6744)
);

OR2x2_ASAP7_75t_L g6745 ( 
.A(n_6542),
.B(n_6634),
.Y(n_6745)
);

AND2x2_ASAP7_75t_L g6746 ( 
.A(n_6532),
.B(n_626),
.Y(n_6746)
);

AND2x2_ASAP7_75t_L g6747 ( 
.A(n_6558),
.B(n_627),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6514),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6537),
.Y(n_6749)
);

AND2x2_ASAP7_75t_L g6750 ( 
.A(n_6505),
.B(n_627),
.Y(n_6750)
);

OAI221xp5_ASAP7_75t_L g6751 ( 
.A1(n_6583),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.C(n_631),
.Y(n_6751)
);

AND2x2_ASAP7_75t_L g6752 ( 
.A(n_6551),
.B(n_628),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6590),
.B(n_628),
.Y(n_6753)
);

NAND3xp33_ASAP7_75t_L g6754 ( 
.A(n_6521),
.B(n_629),
.C(n_631),
.Y(n_6754)
);

AOI33xp33_ASAP7_75t_L g6755 ( 
.A1(n_6582),
.A2(n_633),
.A3(n_635),
.B1(n_629),
.B2(n_632),
.B3(n_634),
.Y(n_6755)
);

OAI22xp33_ASAP7_75t_L g6756 ( 
.A1(n_6625),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_6511),
.B(n_6591),
.Y(n_6757)
);

BUFx2_ASAP7_75t_L g6758 ( 
.A(n_6557),
.Y(n_6758)
);

AND2x2_ASAP7_75t_L g6759 ( 
.A(n_6611),
.B(n_632),
.Y(n_6759)
);

INVx1_ASAP7_75t_L g6760 ( 
.A(n_6627),
.Y(n_6760)
);

OAI22xp5_ASAP7_75t_L g6761 ( 
.A1(n_6555),
.A2(n_6535),
.B1(n_6538),
.B2(n_6608),
.Y(n_6761)
);

NAND3xp33_ASAP7_75t_L g6762 ( 
.A(n_6545),
.B(n_633),
.C(n_634),
.Y(n_6762)
);

NOR2xp33_ASAP7_75t_L g6763 ( 
.A(n_6596),
.B(n_635),
.Y(n_6763)
);

INVx6_ASAP7_75t_L g6764 ( 
.A(n_6616),
.Y(n_6764)
);

INVx3_ASAP7_75t_L g6765 ( 
.A(n_6640),
.Y(n_6765)
);

INVx2_ASAP7_75t_L g6766 ( 
.A(n_6528),
.Y(n_6766)
);

BUFx2_ASAP7_75t_L g6767 ( 
.A(n_6642),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6523),
.Y(n_6768)
);

AND2x2_ASAP7_75t_L g6769 ( 
.A(n_6612),
.B(n_636),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6529),
.Y(n_6770)
);

AND2x2_ASAP7_75t_L g6771 ( 
.A(n_6568),
.B(n_636),
.Y(n_6771)
);

NAND4xp25_ASAP7_75t_L g6772 ( 
.A(n_6630),
.B(n_639),
.C(n_637),
.D(n_638),
.Y(n_6772)
);

NAND2xp5_ASAP7_75t_L g6773 ( 
.A(n_6581),
.B(n_637),
.Y(n_6773)
);

INVx1_ASAP7_75t_L g6774 ( 
.A(n_6503),
.Y(n_6774)
);

AND2x4_ASAP7_75t_SL g6775 ( 
.A(n_6552),
.B(n_640),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6603),
.Y(n_6776)
);

AND2x2_ASAP7_75t_L g6777 ( 
.A(n_6550),
.B(n_641),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6623),
.Y(n_6778)
);

CKINVDCx5p33_ASAP7_75t_R g6779 ( 
.A(n_6556),
.Y(n_6779)
);

AOI221xp5_ASAP7_75t_L g6780 ( 
.A1(n_6573),
.A2(n_645),
.B1(n_642),
.B2(n_644),
.C(n_646),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_6530),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6516),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6516),
.Y(n_6783)
);

HB1xp67_ASAP7_75t_L g6784 ( 
.A(n_6516),
.Y(n_6784)
);

AND2x2_ASAP7_75t_L g6785 ( 
.A(n_6544),
.B(n_642),
.Y(n_6785)
);

AOI221x1_ASAP7_75t_SL g6786 ( 
.A1(n_6526),
.A2(n_645),
.B1(n_642),
.B2(n_644),
.C(n_646),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_6516),
.Y(n_6787)
);

INVx2_ASAP7_75t_L g6788 ( 
.A(n_6539),
.Y(n_6788)
);

AND2x2_ASAP7_75t_L g6789 ( 
.A(n_6544),
.B(n_644),
.Y(n_6789)
);

NAND4xp75_ASAP7_75t_L g6790 ( 
.A(n_6564),
.B(n_648),
.C(n_645),
.D(n_647),
.Y(n_6790)
);

NAND2xp5_ASAP7_75t_L g6791 ( 
.A(n_6546),
.B(n_647),
.Y(n_6791)
);

AND2x2_ASAP7_75t_L g6792 ( 
.A(n_6544),
.B(n_648),
.Y(n_6792)
);

AND2x2_ASAP7_75t_SL g6793 ( 
.A(n_6620),
.B(n_648),
.Y(n_6793)
);

XNOR2xp5_ASAP7_75t_L g6794 ( 
.A(n_6611),
.B(n_649),
.Y(n_6794)
);

OAI31xp33_ASAP7_75t_L g6795 ( 
.A1(n_6499),
.A2(n_651),
.A3(n_649),
.B(n_650),
.Y(n_6795)
);

NAND3xp33_ASAP7_75t_L g6796 ( 
.A(n_6544),
.B(n_649),
.C(n_650),
.Y(n_6796)
);

INVx6_ASAP7_75t_L g6797 ( 
.A(n_6519),
.Y(n_6797)
);

INVx5_ASAP7_75t_L g6798 ( 
.A(n_6519),
.Y(n_6798)
);

A2O1A1O1Ixp25_ASAP7_75t_L g6799 ( 
.A1(n_6661),
.A2(n_652),
.B(n_650),
.C(n_651),
.D(n_653),
.Y(n_6799)
);

NAND2xp5_ASAP7_75t_L g6800 ( 
.A(n_6643),
.B(n_651),
.Y(n_6800)
);

NAND2xp5_ASAP7_75t_L g6801 ( 
.A(n_6652),
.B(n_6788),
.Y(n_6801)
);

INVx1_ASAP7_75t_L g6802 ( 
.A(n_6785),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_6789),
.Y(n_6803)
);

OR2x2_ASAP7_75t_L g6804 ( 
.A(n_6656),
.B(n_652),
.Y(n_6804)
);

NOR2xp33_ASAP7_75t_L g6805 ( 
.A(n_6649),
.B(n_6653),
.Y(n_6805)
);

AOI22xp33_ASAP7_75t_L g6806 ( 
.A1(n_6647),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_6806)
);

OR2x2_ASAP7_75t_L g6807 ( 
.A(n_6693),
.B(n_653),
.Y(n_6807)
);

NOR2x1p5_ASAP7_75t_SL g6808 ( 
.A(n_6720),
.B(n_654),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6792),
.Y(n_6809)
);

NAND2xp5_ASAP7_75t_SL g6810 ( 
.A(n_6798),
.B(n_654),
.Y(n_6810)
);

INVx1_ASAP7_75t_L g6811 ( 
.A(n_6692),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_6645),
.Y(n_6812)
);

AND2x4_ASAP7_75t_L g6813 ( 
.A(n_6666),
.B(n_655),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_6791),
.Y(n_6814)
);

AOI22xp5_ASAP7_75t_L g6815 ( 
.A1(n_6764),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.Y(n_6815)
);

NAND3xp33_ASAP7_75t_SL g6816 ( 
.A(n_6779),
.B(n_655),
.C(n_656),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_6682),
.Y(n_6817)
);

AND2x2_ASAP7_75t_L g6818 ( 
.A(n_6735),
.B(n_657),
.Y(n_6818)
);

OR2x2_ASAP7_75t_L g6819 ( 
.A(n_6669),
.B(n_658),
.Y(n_6819)
);

HB1xp67_ASAP7_75t_L g6820 ( 
.A(n_6694),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6759),
.Y(n_6821)
);

NAND2xp5_ASAP7_75t_SL g6822 ( 
.A(n_6798),
.B(n_658),
.Y(n_6822)
);

OAI21xp33_ASAP7_75t_L g6823 ( 
.A1(n_6696),
.A2(n_659),
.B(n_660),
.Y(n_6823)
);

AOI22xp5_ASAP7_75t_L g6824 ( 
.A1(n_6764),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.Y(n_6824)
);

NAND2xp5_ASAP7_75t_L g6825 ( 
.A(n_6798),
.B(n_659),
.Y(n_6825)
);

INVx1_ASAP7_75t_SL g6826 ( 
.A(n_6797),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_6695),
.Y(n_6827)
);

AND2x4_ASAP7_75t_L g6828 ( 
.A(n_6698),
.B(n_661),
.Y(n_6828)
);

INVxp67_ASAP7_75t_L g6829 ( 
.A(n_6736),
.Y(n_6829)
);

AND2x2_ASAP7_75t_L g6830 ( 
.A(n_6681),
.B(n_661),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6685),
.Y(n_6831)
);

OAI211xp5_ASAP7_75t_L g6832 ( 
.A1(n_6733),
.A2(n_664),
.B(n_662),
.C(n_663),
.Y(n_6832)
);

AND2x2_ASAP7_75t_L g6833 ( 
.A(n_6676),
.B(n_662),
.Y(n_6833)
);

AO221x1_ASAP7_75t_L g6834 ( 
.A1(n_6728),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.C(n_666),
.Y(n_6834)
);

INVx1_ASAP7_75t_L g6835 ( 
.A(n_6793),
.Y(n_6835)
);

OR2x2_ASAP7_75t_L g6836 ( 
.A(n_6701),
.B(n_663),
.Y(n_6836)
);

NAND2xp5_ASAP7_75t_SL g6837 ( 
.A(n_6795),
.B(n_664),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6678),
.B(n_665),
.Y(n_6838)
);

INVx3_ASAP7_75t_L g6839 ( 
.A(n_6797),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_6697),
.Y(n_6840)
);

AOI22xp5_ASAP7_75t_L g6841 ( 
.A1(n_6781),
.A2(n_6729),
.B1(n_6774),
.B2(n_6769),
.Y(n_6841)
);

AND2x4_ASAP7_75t_L g6842 ( 
.A(n_6664),
.B(n_665),
.Y(n_6842)
);

OR2x2_ASAP7_75t_L g6843 ( 
.A(n_6738),
.B(n_666),
.Y(n_6843)
);

AND2x2_ASAP7_75t_L g6844 ( 
.A(n_6663),
.B(n_666),
.Y(n_6844)
);

INVx2_ASAP7_75t_L g6845 ( 
.A(n_6702),
.Y(n_6845)
);

INVxp67_ASAP7_75t_L g6846 ( 
.A(n_6790),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6659),
.Y(n_6847)
);

AOI32xp33_ASAP7_75t_L g6848 ( 
.A1(n_6767),
.A2(n_669),
.A3(n_667),
.B1(n_668),
.B2(n_670),
.Y(n_6848)
);

INVxp33_ASAP7_75t_L g6849 ( 
.A(n_6794),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_L g6850 ( 
.A(n_6786),
.B(n_667),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_6784),
.Y(n_6851)
);

INVx3_ASAP7_75t_L g6852 ( 
.A(n_6683),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6658),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6718),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_6665),
.B(n_668),
.Y(n_6855)
);

INVx4_ASAP7_75t_L g6856 ( 
.A(n_6734),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_6700),
.Y(n_6857)
);

NAND4xp25_ASAP7_75t_L g6858 ( 
.A(n_6674),
.B(n_671),
.C(n_669),
.D(n_670),
.Y(n_6858)
);

OR2x2_ASAP7_75t_L g6859 ( 
.A(n_6705),
.B(n_669),
.Y(n_6859)
);

OR2x2_ASAP7_75t_L g6860 ( 
.A(n_6796),
.B(n_670),
.Y(n_6860)
);

OR2x2_ASAP7_75t_L g6861 ( 
.A(n_6691),
.B(n_671),
.Y(n_6861)
);

NAND2xp5_ASAP7_75t_L g6862 ( 
.A(n_6721),
.B(n_671),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6688),
.Y(n_6863)
);

INVxp67_ASAP7_75t_L g6864 ( 
.A(n_6752),
.Y(n_6864)
);

NAND2xp5_ASAP7_75t_L g6865 ( 
.A(n_6737),
.B(n_672),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6655),
.Y(n_6866)
);

NAND2x1_ASAP7_75t_L g6867 ( 
.A(n_6707),
.B(n_672),
.Y(n_6867)
);

AND2x2_ASAP7_75t_L g6868 ( 
.A(n_6703),
.B(n_672),
.Y(n_6868)
);

NOR2x1_ASAP7_75t_L g6869 ( 
.A(n_6680),
.B(n_673),
.Y(n_6869)
);

INVx2_ASAP7_75t_L g6870 ( 
.A(n_6711),
.Y(n_6870)
);

AND2x2_ASAP7_75t_L g6871 ( 
.A(n_6670),
.B(n_673),
.Y(n_6871)
);

INVxp67_ASAP7_75t_SL g6872 ( 
.A(n_6719),
.Y(n_6872)
);

INVx1_ASAP7_75t_L g6873 ( 
.A(n_6657),
.Y(n_6873)
);

AND2x2_ASAP7_75t_L g6874 ( 
.A(n_6677),
.B(n_674),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6699),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6679),
.B(n_674),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6651),
.B(n_675),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_6714),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6723),
.Y(n_6879)
);

AND2x2_ASAP7_75t_L g6880 ( 
.A(n_6746),
.B(n_675),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_6650),
.B(n_676),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6706),
.Y(n_6882)
);

OAI21xp33_ASAP7_75t_L g6883 ( 
.A1(n_6757),
.A2(n_677),
.B(n_678),
.Y(n_6883)
);

INVxp67_ASAP7_75t_SL g6884 ( 
.A(n_6773),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_6644),
.Y(n_6885)
);

AND2x2_ASAP7_75t_L g6886 ( 
.A(n_6753),
.B(n_677),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_L g6887 ( 
.A(n_6675),
.B(n_6777),
.Y(n_6887)
);

INVx2_ASAP7_75t_L g6888 ( 
.A(n_6770),
.Y(n_6888)
);

AND2x4_ASAP7_75t_L g6889 ( 
.A(n_6768),
.B(n_6712),
.Y(n_6889)
);

NOR2x1p5_ASAP7_75t_L g6890 ( 
.A(n_6766),
.B(n_679),
.Y(n_6890)
);

NOR2xp33_ASAP7_75t_L g6891 ( 
.A(n_6710),
.B(n_679),
.Y(n_6891)
);

OR2x2_ASAP7_75t_L g6892 ( 
.A(n_6740),
.B(n_679),
.Y(n_6892)
);

INVx2_ASAP7_75t_L g6893 ( 
.A(n_6716),
.Y(n_6893)
);

INVx1_ASAP7_75t_L g6894 ( 
.A(n_6782),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_6783),
.Y(n_6895)
);

INVx1_ASAP7_75t_SL g6896 ( 
.A(n_6722),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6787),
.Y(n_6897)
);

NAND2xp5_ASAP7_75t_L g6898 ( 
.A(n_6771),
.B(n_680),
.Y(n_6898)
);

AND2x2_ASAP7_75t_L g6899 ( 
.A(n_6660),
.B(n_681),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6750),
.Y(n_6900)
);

OR2x2_ASAP7_75t_L g6901 ( 
.A(n_6772),
.B(n_682),
.Y(n_6901)
);

INVx1_ASAP7_75t_L g6902 ( 
.A(n_6755),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6648),
.Y(n_6903)
);

OAI21xp5_ASAP7_75t_L g6904 ( 
.A1(n_6713),
.A2(n_682),
.B(n_684),
.Y(n_6904)
);

OR2x2_ASAP7_75t_L g6905 ( 
.A(n_6731),
.B(n_682),
.Y(n_6905)
);

INVx1_ASAP7_75t_SL g6906 ( 
.A(n_6745),
.Y(n_6906)
);

INVx1_ASAP7_75t_L g6907 ( 
.A(n_6747),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_6686),
.Y(n_6908)
);

OR2x2_ASAP7_75t_L g6909 ( 
.A(n_6801),
.B(n_6725),
.Y(n_6909)
);

INVxp67_ASAP7_75t_SL g6910 ( 
.A(n_6805),
.Y(n_6910)
);

OAI22xp33_ASAP7_75t_L g6911 ( 
.A1(n_6815),
.A2(n_6824),
.B1(n_6799),
.B2(n_6856),
.Y(n_6911)
);

INVx2_ASAP7_75t_SL g6912 ( 
.A(n_6845),
.Y(n_6912)
);

OAI211xp5_ASAP7_75t_L g6913 ( 
.A1(n_6806),
.A2(n_6741),
.B(n_6744),
.C(n_6743),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6830),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6820),
.Y(n_6915)
);

INVx1_ASAP7_75t_SL g6916 ( 
.A(n_6826),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_6800),
.Y(n_6917)
);

INVx2_ASAP7_75t_SL g6918 ( 
.A(n_6839),
.Y(n_6918)
);

NAND2xp5_ASAP7_75t_SL g6919 ( 
.A(n_6828),
.B(n_6761),
.Y(n_6919)
);

INVx2_ASAP7_75t_SL g6920 ( 
.A(n_6852),
.Y(n_6920)
);

OAI21xp33_ASAP7_75t_L g6921 ( 
.A1(n_6849),
.A2(n_6776),
.B(n_6646),
.Y(n_6921)
);

OAI32xp33_ASAP7_75t_L g6922 ( 
.A1(n_6906),
.A2(n_6778),
.A3(n_6760),
.B1(n_6654),
.B2(n_6689),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6828),
.Y(n_6923)
);

OAI21xp33_ASAP7_75t_L g6924 ( 
.A1(n_6823),
.A2(n_6690),
.B(n_6668),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_6813),
.Y(n_6925)
);

INVx2_ASAP7_75t_L g6926 ( 
.A(n_6842),
.Y(n_6926)
);

OR2x2_ASAP7_75t_L g6927 ( 
.A(n_6812),
.B(n_6739),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6813),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6825),
.Y(n_6929)
);

OAI21xp5_ASAP7_75t_L g6930 ( 
.A1(n_6869),
.A2(n_6717),
.B(n_6687),
.Y(n_6930)
);

NAND2xp5_ASAP7_75t_L g6931 ( 
.A(n_6834),
.B(n_6704),
.Y(n_6931)
);

OAI32xp33_ASAP7_75t_L g6932 ( 
.A1(n_6887),
.A2(n_6708),
.A3(n_6684),
.B1(n_6667),
.B2(n_6749),
.Y(n_6932)
);

INVx1_ASAP7_75t_L g6933 ( 
.A(n_6877),
.Y(n_6933)
);

NAND2xp5_ASAP7_75t_L g6934 ( 
.A(n_6872),
.B(n_6780),
.Y(n_6934)
);

O2A1O1Ixp33_ASAP7_75t_L g6935 ( 
.A1(n_6810),
.A2(n_6742),
.B(n_6756),
.C(n_6751),
.Y(n_6935)
);

INVx2_ASAP7_75t_SL g6936 ( 
.A(n_6811),
.Y(n_6936)
);

OAI22xp33_ASAP7_75t_SL g6937 ( 
.A1(n_6867),
.A2(n_6822),
.B1(n_6838),
.B2(n_6837),
.Y(n_6937)
);

AOI32xp33_ASAP7_75t_L g6938 ( 
.A1(n_6902),
.A2(n_6767),
.A3(n_6765),
.B1(n_6758),
.B2(n_6775),
.Y(n_6938)
);

XNOR2xp5_ASAP7_75t_L g6939 ( 
.A(n_6858),
.B(n_6841),
.Y(n_6939)
);

NOR2xp67_ASAP7_75t_SL g6940 ( 
.A(n_6888),
.B(n_6840),
.Y(n_6940)
);

NAND3xp33_ASAP7_75t_L g6941 ( 
.A(n_6848),
.B(n_6726),
.C(n_6762),
.Y(n_6941)
);

OAI21xp5_ASAP7_75t_L g6942 ( 
.A1(n_6846),
.A2(n_6754),
.B(n_6671),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6859),
.Y(n_6943)
);

AND2x2_ASAP7_75t_L g6944 ( 
.A(n_6833),
.B(n_6748),
.Y(n_6944)
);

INVx1_ASAP7_75t_L g6945 ( 
.A(n_6861),
.Y(n_6945)
);

INVx2_ASAP7_75t_L g6946 ( 
.A(n_6893),
.Y(n_6946)
);

INVx1_ASAP7_75t_L g6947 ( 
.A(n_6836),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6807),
.Y(n_6948)
);

AOI22xp5_ASAP7_75t_L g6949 ( 
.A1(n_6816),
.A2(n_6763),
.B1(n_6732),
.B2(n_6673),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6819),
.Y(n_6950)
);

A2O1A1Ixp33_ASAP7_75t_L g6951 ( 
.A1(n_6808),
.A2(n_6883),
.B(n_6891),
.C(n_6832),
.Y(n_6951)
);

A2O1A1Ixp33_ASAP7_75t_L g6952 ( 
.A1(n_6847),
.A2(n_6727),
.B(n_6662),
.C(n_6715),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_6860),
.Y(n_6953)
);

INVx2_ASAP7_75t_L g6954 ( 
.A(n_6870),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6804),
.Y(n_6955)
);

INVx2_ASAP7_75t_L g6956 ( 
.A(n_6889),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6899),
.B(n_6730),
.Y(n_6957)
);

HB1xp67_ASAP7_75t_L g6958 ( 
.A(n_6873),
.Y(n_6958)
);

AND2x2_ASAP7_75t_L g6959 ( 
.A(n_6868),
.B(n_6709),
.Y(n_6959)
);

OAI21xp33_ASAP7_75t_L g6960 ( 
.A1(n_6821),
.A2(n_6672),
.B(n_6724),
.Y(n_6960)
);

INVx1_ASAP7_75t_L g6961 ( 
.A(n_6901),
.Y(n_6961)
);

NAND2xp5_ASAP7_75t_L g6962 ( 
.A(n_6871),
.B(n_6672),
.Y(n_6962)
);

AOI321xp33_ASAP7_75t_L g6963 ( 
.A1(n_6866),
.A2(n_6908),
.A3(n_6882),
.B1(n_6851),
.B2(n_6884),
.C(n_6857),
.Y(n_6963)
);

INVx2_ASAP7_75t_SL g6964 ( 
.A(n_6889),
.Y(n_6964)
);

NOR3xp33_ASAP7_75t_L g6965 ( 
.A(n_6881),
.B(n_684),
.C(n_685),
.Y(n_6965)
);

AND2x2_ASAP7_75t_L g6966 ( 
.A(n_6874),
.B(n_684),
.Y(n_6966)
);

NOR2xp33_ASAP7_75t_L g6967 ( 
.A(n_6850),
.B(n_685),
.Y(n_6967)
);

INVx2_ASAP7_75t_SL g6968 ( 
.A(n_6854),
.Y(n_6968)
);

AND2x2_ASAP7_75t_L g6969 ( 
.A(n_6855),
.B(n_685),
.Y(n_6969)
);

NAND2x2_ASAP7_75t_L g6970 ( 
.A(n_6890),
.B(n_686),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6876),
.Y(n_6971)
);

NAND2xp5_ASAP7_75t_L g6972 ( 
.A(n_6818),
.B(n_686),
.Y(n_6972)
);

OR2x2_ASAP7_75t_L g6973 ( 
.A(n_6898),
.B(n_686),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_6844),
.Y(n_6974)
);

OR2x6_ASAP7_75t_L g6975 ( 
.A(n_6904),
.B(n_687),
.Y(n_6975)
);

OAI32xp33_ASAP7_75t_L g6976 ( 
.A1(n_6896),
.A2(n_689),
.A3(n_687),
.B1(n_688),
.B2(n_690),
.Y(n_6976)
);

NAND2xp5_ASAP7_75t_L g6977 ( 
.A(n_6886),
.B(n_687),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6892),
.Y(n_6978)
);

AOI221xp5_ASAP7_75t_L g6979 ( 
.A1(n_6802),
.A2(n_690),
.B1(n_688),
.B2(n_689),
.C(n_691),
.Y(n_6979)
);

AOI32xp33_ASAP7_75t_L g6980 ( 
.A1(n_6835),
.A2(n_690),
.A3(n_688),
.B1(n_689),
.B2(n_691),
.Y(n_6980)
);

INVx1_ASAP7_75t_L g6981 ( 
.A(n_6880),
.Y(n_6981)
);

AND2x2_ASAP7_75t_L g6982 ( 
.A(n_6803),
.B(n_691),
.Y(n_6982)
);

AND2x4_ASAP7_75t_L g6983 ( 
.A(n_6817),
.B(n_692),
.Y(n_6983)
);

INVx1_ASAP7_75t_SL g6984 ( 
.A(n_6843),
.Y(n_6984)
);

INVx2_ASAP7_75t_L g6985 ( 
.A(n_6827),
.Y(n_6985)
);

INVx2_ASAP7_75t_L g6986 ( 
.A(n_6879),
.Y(n_6986)
);

OA22x2_ASAP7_75t_L g6987 ( 
.A1(n_6809),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_6987)
);

AOI22xp5_ASAP7_75t_L g6988 ( 
.A1(n_6900),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_6988)
);

AND2x2_ASAP7_75t_L g6989 ( 
.A(n_6863),
.B(n_693),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6865),
.Y(n_6990)
);

INVx1_ASAP7_75t_SL g6991 ( 
.A(n_6905),
.Y(n_6991)
);

NAND2xp5_ASAP7_75t_L g6992 ( 
.A(n_6907),
.B(n_694),
.Y(n_6992)
);

NAND2xp5_ASAP7_75t_L g6993 ( 
.A(n_6875),
.B(n_6878),
.Y(n_6993)
);

INVx2_ASAP7_75t_L g6994 ( 
.A(n_6853),
.Y(n_6994)
);

OR2x2_ASAP7_75t_L g6995 ( 
.A(n_6862),
.B(n_695),
.Y(n_6995)
);

AOI22xp33_ASAP7_75t_L g6996 ( 
.A1(n_6885),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.Y(n_6996)
);

NOR2xp33_ASAP7_75t_L g6997 ( 
.A(n_6864),
.B(n_696),
.Y(n_6997)
);

INVx1_ASAP7_75t_L g6998 ( 
.A(n_6894),
.Y(n_6998)
);

NAND2xp5_ASAP7_75t_L g6999 ( 
.A(n_6831),
.B(n_6814),
.Y(n_6999)
);

OR2x2_ASAP7_75t_L g7000 ( 
.A(n_6895),
.B(n_696),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6897),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6903),
.B(n_697),
.Y(n_7002)
);

OR2x2_ASAP7_75t_L g7003 ( 
.A(n_6829),
.B(n_697),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6801),
.Y(n_7004)
);

AND2x2_ASAP7_75t_L g7005 ( 
.A(n_6830),
.B(n_698),
.Y(n_7005)
);

NAND2xp5_ASAP7_75t_L g7006 ( 
.A(n_6828),
.B(n_698),
.Y(n_7006)
);

OR2x2_ASAP7_75t_L g7007 ( 
.A(n_6801),
.B(n_699),
.Y(n_7007)
);

AOI22xp5_ASAP7_75t_L g7008 ( 
.A1(n_6805),
.A2(n_701),
.B1(n_699),
.B2(n_700),
.Y(n_7008)
);

HB1xp67_ASAP7_75t_L g7009 ( 
.A(n_6828),
.Y(n_7009)
);

AO21x1_ASAP7_75t_L g7010 ( 
.A1(n_6805),
.A2(n_699),
.B(n_700),
.Y(n_7010)
);

BUFx2_ASAP7_75t_L g7011 ( 
.A(n_6828),
.Y(n_7011)
);

OR2x2_ASAP7_75t_L g7012 ( 
.A(n_6801),
.B(n_700),
.Y(n_7012)
);

INVx1_ASAP7_75t_SL g7013 ( 
.A(n_6801),
.Y(n_7013)
);

AOI21xp33_ASAP7_75t_L g7014 ( 
.A1(n_6849),
.A2(n_702),
.B(n_703),
.Y(n_7014)
);

OA21x2_ASAP7_75t_L g7015 ( 
.A1(n_6805),
.A2(n_702),
.B(n_703),
.Y(n_7015)
);

NAND2xp5_ASAP7_75t_L g7016 ( 
.A(n_6828),
.B(n_702),
.Y(n_7016)
);

OR2x2_ASAP7_75t_L g7017 ( 
.A(n_6801),
.B(n_703),
.Y(n_7017)
);

AOI31xp33_ASAP7_75t_L g7018 ( 
.A1(n_6805),
.A2(n_706),
.A3(n_704),
.B(n_705),
.Y(n_7018)
);

AND2x2_ASAP7_75t_L g7019 ( 
.A(n_6830),
.B(n_704),
.Y(n_7019)
);

XNOR2x2_ASAP7_75t_L g7020 ( 
.A(n_6805),
.B(n_706),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6801),
.Y(n_7021)
);

AND2x2_ASAP7_75t_L g7022 ( 
.A(n_6916),
.B(n_6910),
.Y(n_7022)
);

INVx1_ASAP7_75t_L g7023 ( 
.A(n_6964),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6956),
.Y(n_7024)
);

NAND2xp5_ASAP7_75t_L g7025 ( 
.A(n_6912),
.B(n_6918),
.Y(n_7025)
);

OR2x2_ASAP7_75t_L g7026 ( 
.A(n_7013),
.B(n_706),
.Y(n_7026)
);

INVx1_ASAP7_75t_SL g7027 ( 
.A(n_6946),
.Y(n_7027)
);

BUFx2_ASAP7_75t_L g7028 ( 
.A(n_6954),
.Y(n_7028)
);

HB1xp67_ASAP7_75t_L g7029 ( 
.A(n_7009),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_7005),
.B(n_707),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6987),
.Y(n_7031)
);

NOR2x1p5_ASAP7_75t_L g7032 ( 
.A(n_6931),
.B(n_707),
.Y(n_7032)
);

HB1xp67_ASAP7_75t_L g7033 ( 
.A(n_7015),
.Y(n_7033)
);

OR2x2_ASAP7_75t_L g7034 ( 
.A(n_7006),
.B(n_708),
.Y(n_7034)
);

INVx1_ASAP7_75t_SL g7035 ( 
.A(n_6909),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_6920),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_7019),
.B(n_708),
.Y(n_7037)
);

INVx1_ASAP7_75t_SL g7038 ( 
.A(n_6915),
.Y(n_7038)
);

HB1xp67_ASAP7_75t_L g7039 ( 
.A(n_7015),
.Y(n_7039)
);

AND2x2_ASAP7_75t_L g7040 ( 
.A(n_6966),
.B(n_708),
.Y(n_7040)
);

AOI22xp5_ASAP7_75t_L g7041 ( 
.A1(n_7004),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.Y(n_7041)
);

AND2x2_ASAP7_75t_L g7042 ( 
.A(n_6969),
.B(n_709),
.Y(n_7042)
);

OR2x2_ASAP7_75t_L g7043 ( 
.A(n_7016),
.B(n_709),
.Y(n_7043)
);

NAND2xp5_ASAP7_75t_L g7044 ( 
.A(n_6968),
.B(n_710),
.Y(n_7044)
);

AND2x4_ASAP7_75t_L g7045 ( 
.A(n_6926),
.B(n_711),
.Y(n_7045)
);

NAND2xp5_ASAP7_75t_L g7046 ( 
.A(n_6983),
.B(n_7011),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_L g7047 ( 
.A(n_6983),
.B(n_712),
.Y(n_7047)
);

AND2x4_ASAP7_75t_SL g7048 ( 
.A(n_7021),
.B(n_6944),
.Y(n_7048)
);

OR2x2_ASAP7_75t_L g7049 ( 
.A(n_7007),
.B(n_713),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6958),
.Y(n_7050)
);

INVx1_ASAP7_75t_SL g7051 ( 
.A(n_6925),
.Y(n_7051)
);

INVx3_ASAP7_75t_L g7052 ( 
.A(n_6985),
.Y(n_7052)
);

OR2x2_ASAP7_75t_L g7053 ( 
.A(n_7012),
.B(n_713),
.Y(n_7053)
);

CKINVDCx16_ASAP7_75t_R g7054 ( 
.A(n_7017),
.Y(n_7054)
);

INVx2_ASAP7_75t_L g7055 ( 
.A(n_6936),
.Y(n_7055)
);

OR2x2_ASAP7_75t_L g7056 ( 
.A(n_6923),
.B(n_713),
.Y(n_7056)
);

INVx1_ASAP7_75t_SL g7057 ( 
.A(n_6928),
.Y(n_7057)
);

INVx2_ASAP7_75t_L g7058 ( 
.A(n_6986),
.Y(n_7058)
);

NAND2xp5_ASAP7_75t_L g7059 ( 
.A(n_6982),
.B(n_714),
.Y(n_7059)
);

HB1xp67_ASAP7_75t_L g7060 ( 
.A(n_6945),
.Y(n_7060)
);

INVx1_ASAP7_75t_SL g7061 ( 
.A(n_6984),
.Y(n_7061)
);

AO21x2_ASAP7_75t_L g7062 ( 
.A1(n_6942),
.A2(n_714),
.B(n_715),
.Y(n_7062)
);

AOI22xp33_ASAP7_75t_L g7063 ( 
.A1(n_6965),
.A2(n_716),
.B1(n_714),
.B2(n_715),
.Y(n_7063)
);

INVx1_ASAP7_75t_L g7064 ( 
.A(n_7010),
.Y(n_7064)
);

INVx2_ASAP7_75t_L g7065 ( 
.A(n_6994),
.Y(n_7065)
);

NAND2xp5_ASAP7_75t_L g7066 ( 
.A(n_6989),
.B(n_716),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6940),
.Y(n_7067)
);

AND2x4_ASAP7_75t_SL g7068 ( 
.A(n_6961),
.B(n_716),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_7018),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_7002),
.Y(n_7070)
);

AND2x2_ASAP7_75t_L g7071 ( 
.A(n_6914),
.B(n_6959),
.Y(n_7071)
);

OAI22xp5_ASAP7_75t_SL g7072 ( 
.A1(n_6941),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_7000),
.Y(n_7073)
);

INVx1_ASAP7_75t_SL g7074 ( 
.A(n_6991),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6972),
.Y(n_7075)
);

OR2x2_ASAP7_75t_L g7076 ( 
.A(n_7003),
.B(n_717),
.Y(n_7076)
);

INVx2_ASAP7_75t_L g7077 ( 
.A(n_6950),
.Y(n_7077)
);

AOI22xp33_ASAP7_75t_L g7078 ( 
.A1(n_6970),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_7078)
);

INVx2_ASAP7_75t_L g7079 ( 
.A(n_6955),
.Y(n_7079)
);

NOR2xp33_ASAP7_75t_L g7080 ( 
.A(n_6911),
.B(n_718),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_6996),
.B(n_719),
.Y(n_7081)
);

OR2x2_ASAP7_75t_L g7082 ( 
.A(n_6977),
.B(n_720),
.Y(n_7082)
);

OR2x2_ASAP7_75t_L g7083 ( 
.A(n_6973),
.B(n_721),
.Y(n_7083)
);

HB1xp67_ASAP7_75t_L g7084 ( 
.A(n_6943),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_7020),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6980),
.B(n_721),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6976),
.Y(n_7087)
);

AND2x2_ASAP7_75t_SL g7088 ( 
.A(n_7045),
.B(n_6967),
.Y(n_7088)
);

OAI321xp33_ASAP7_75t_L g7089 ( 
.A1(n_7025),
.A2(n_6963),
.A3(n_6938),
.B1(n_6921),
.B2(n_6934),
.C(n_6924),
.Y(n_7089)
);

OAI32xp33_ASAP7_75t_L g7090 ( 
.A1(n_7027),
.A2(n_6962),
.A3(n_6995),
.B1(n_6927),
.B2(n_6957),
.Y(n_7090)
);

INVx1_ASAP7_75t_L g7091 ( 
.A(n_7022),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_7023),
.Y(n_7092)
);

AOI21xp33_ASAP7_75t_L g7093 ( 
.A1(n_7080),
.A2(n_6939),
.B(n_6997),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_7028),
.Y(n_7094)
);

AND2x2_ASAP7_75t_L g7095 ( 
.A(n_7035),
.B(n_6933),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_7024),
.B(n_6971),
.Y(n_7096)
);

OR2x2_ASAP7_75t_L g7097 ( 
.A(n_7036),
.B(n_6919),
.Y(n_7097)
);

AND2x2_ASAP7_75t_L g7098 ( 
.A(n_7048),
.B(n_6974),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_7029),
.Y(n_7099)
);

INVx1_ASAP7_75t_L g7100 ( 
.A(n_7072),
.Y(n_7100)
);

AOI222xp33_ASAP7_75t_L g7101 ( 
.A1(n_7067),
.A2(n_6960),
.B1(n_6930),
.B2(n_7001),
.C1(n_6998),
.C2(n_6947),
.Y(n_7101)
);

AOI22xp5_ASAP7_75t_L g7102 ( 
.A1(n_7038),
.A2(n_6913),
.B1(n_6948),
.B2(n_6953),
.Y(n_7102)
);

NAND2xp5_ASAP7_75t_SL g7103 ( 
.A(n_7045),
.B(n_6937),
.Y(n_7103)
);

INVxp67_ASAP7_75t_L g7104 ( 
.A(n_7047),
.Y(n_7104)
);

INVx2_ASAP7_75t_L g7105 ( 
.A(n_7058),
.Y(n_7105)
);

OAI22xp5_ASAP7_75t_L g7106 ( 
.A1(n_7078),
.A2(n_6949),
.B1(n_6951),
.B2(n_6992),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_7056),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_7031),
.Y(n_7108)
);

AND2x2_ASAP7_75t_L g7109 ( 
.A(n_7030),
.B(n_6981),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_7068),
.Y(n_7110)
);

INVxp67_ASAP7_75t_L g7111 ( 
.A(n_7046),
.Y(n_7111)
);

AOI21xp33_ASAP7_75t_SL g7112 ( 
.A1(n_7085),
.A2(n_7014),
.B(n_6935),
.Y(n_7112)
);

AOI21xp33_ASAP7_75t_SL g7113 ( 
.A1(n_7086),
.A2(n_6993),
.B(n_6990),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_7055),
.Y(n_7114)
);

AOI332xp33_ASAP7_75t_L g7115 ( 
.A1(n_7050),
.A2(n_6929),
.A3(n_6917),
.B1(n_6978),
.B2(n_6999),
.B3(n_6922),
.C1(n_6988),
.C2(n_7008),
.Y(n_7115)
);

AOI21xp5_ASAP7_75t_L g7116 ( 
.A1(n_7059),
.A2(n_6952),
.B(n_6932),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_7026),
.Y(n_7117)
);

NOR2xp33_ASAP7_75t_R g7118 ( 
.A(n_7052),
.B(n_721),
.Y(n_7118)
);

O2A1O1Ixp33_ASAP7_75t_L g7119 ( 
.A1(n_7033),
.A2(n_6979),
.B(n_6975),
.C(n_725),
.Y(n_7119)
);

INVx1_ASAP7_75t_L g7120 ( 
.A(n_7071),
.Y(n_7120)
);

O2A1O1Ixp33_ASAP7_75t_L g7121 ( 
.A1(n_7039),
.A2(n_6975),
.B(n_725),
.C(n_723),
.Y(n_7121)
);

AOI222xp33_ASAP7_75t_L g7122 ( 
.A1(n_7061),
.A2(n_725),
.B1(n_727),
.B2(n_723),
.C1(n_724),
.C2(n_726),
.Y(n_7122)
);

INVx1_ASAP7_75t_L g7123 ( 
.A(n_7044),
.Y(n_7123)
);

NAND2xp5_ASAP7_75t_L g7124 ( 
.A(n_7052),
.B(n_723),
.Y(n_7124)
);

AND2x2_ASAP7_75t_L g7125 ( 
.A(n_7040),
.B(n_724),
.Y(n_7125)
);

NOR2x1_ASAP7_75t_L g7126 ( 
.A(n_7032),
.B(n_724),
.Y(n_7126)
);

INVx2_ASAP7_75t_L g7127 ( 
.A(n_7065),
.Y(n_7127)
);

AOI22xp5_ASAP7_75t_L g7128 ( 
.A1(n_7074),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_7060),
.Y(n_7129)
);

NAND2xp5_ASAP7_75t_L g7130 ( 
.A(n_7042),
.B(n_726),
.Y(n_7130)
);

INVx1_ASAP7_75t_L g7131 ( 
.A(n_7049),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_SL g7132 ( 
.A(n_7087),
.B(n_728),
.Y(n_7132)
);

INVx2_ASAP7_75t_L g7133 ( 
.A(n_7077),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_7053),
.Y(n_7134)
);

INVxp67_ASAP7_75t_L g7135 ( 
.A(n_7062),
.Y(n_7135)
);

A2O1A1Ixp33_ASAP7_75t_L g7136 ( 
.A1(n_7041),
.A2(n_731),
.B(n_729),
.C(n_730),
.Y(n_7136)
);

INVx2_ASAP7_75t_L g7137 ( 
.A(n_7079),
.Y(n_7137)
);

AOI22xp5_ASAP7_75t_L g7138 ( 
.A1(n_7051),
.A2(n_731),
.B1(n_729),
.B2(n_730),
.Y(n_7138)
);

NAND2xp5_ASAP7_75t_L g7139 ( 
.A(n_7057),
.B(n_729),
.Y(n_7139)
);

AND2x2_ASAP7_75t_L g7140 ( 
.A(n_7069),
.B(n_731),
.Y(n_7140)
);

NAND2xp5_ASAP7_75t_L g7141 ( 
.A(n_7064),
.B(n_732),
.Y(n_7141)
);

INVxp67_ASAP7_75t_L g7142 ( 
.A(n_7084),
.Y(n_7142)
);

INVxp67_ASAP7_75t_L g7143 ( 
.A(n_7037),
.Y(n_7143)
);

AOI22xp33_ASAP7_75t_L g7144 ( 
.A1(n_7070),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.Y(n_7144)
);

NOR2xp67_ASAP7_75t_SL g7145 ( 
.A(n_7034),
.B(n_7043),
.Y(n_7145)
);

OAI321xp33_ASAP7_75t_L g7146 ( 
.A1(n_7073),
.A2(n_734),
.A3(n_736),
.B1(n_732),
.B2(n_733),
.C(n_735),
.Y(n_7146)
);

NAND2xp5_ASAP7_75t_SL g7147 ( 
.A(n_7054),
.B(n_734),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_7063),
.B(n_735),
.Y(n_7148)
);

NOR2xp67_ASAP7_75t_L g7149 ( 
.A(n_7083),
.B(n_7082),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_7066),
.B(n_735),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_7076),
.Y(n_7151)
);

INVx2_ASAP7_75t_L g7152 ( 
.A(n_7075),
.Y(n_7152)
);

INVxp67_ASAP7_75t_L g7153 ( 
.A(n_7081),
.Y(n_7153)
);

NAND2xp5_ASAP7_75t_L g7154 ( 
.A(n_7022),
.B(n_736),
.Y(n_7154)
);

OAI221xp5_ASAP7_75t_L g7155 ( 
.A1(n_7078),
.A2(n_738),
.B1(n_736),
.B2(n_737),
.C(n_739),
.Y(n_7155)
);

AOI221xp5_ASAP7_75t_L g7156 ( 
.A1(n_7080),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.C(n_740),
.Y(n_7156)
);

OAI21xp33_ASAP7_75t_SL g7157 ( 
.A1(n_7080),
.A2(n_738),
.B(n_739),
.Y(n_7157)
);

A2O1A1Ixp33_ASAP7_75t_L g7158 ( 
.A1(n_7080),
.A2(n_743),
.B(n_741),
.C(n_742),
.Y(n_7158)
);

INVx1_ASAP7_75t_L g7159 ( 
.A(n_7022),
.Y(n_7159)
);

OR2x2_ASAP7_75t_L g7160 ( 
.A(n_7025),
.B(n_741),
.Y(n_7160)
);

INVxp67_ASAP7_75t_L g7161 ( 
.A(n_7022),
.Y(n_7161)
);

INVxp67_ASAP7_75t_L g7162 ( 
.A(n_7022),
.Y(n_7162)
);

AND2x2_ASAP7_75t_L g7163 ( 
.A(n_7022),
.B(n_742),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_7022),
.Y(n_7164)
);

AOI222xp33_ASAP7_75t_L g7165 ( 
.A1(n_7027),
.A2(n_746),
.B1(n_748),
.B2(n_743),
.C1(n_744),
.C2(n_747),
.Y(n_7165)
);

OAI32xp33_ASAP7_75t_L g7166 ( 
.A1(n_7027),
.A2(n_746),
.A3(n_743),
.B1(n_744),
.B2(n_747),
.Y(n_7166)
);

AOI222xp33_ASAP7_75t_L g7167 ( 
.A1(n_7027),
.A2(n_747),
.B1(n_749),
.B2(n_744),
.C1(n_746),
.C2(n_748),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_7022),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_7022),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_7022),
.B(n_748),
.Y(n_7170)
);

NAND2xp5_ASAP7_75t_L g7171 ( 
.A(n_7105),
.B(n_749),
.Y(n_7171)
);

NAND2xp5_ASAP7_75t_L g7172 ( 
.A(n_7127),
.B(n_749),
.Y(n_7172)
);

INVx1_ASAP7_75t_L g7173 ( 
.A(n_7097),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_7163),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_7154),
.Y(n_7175)
);

HB1xp67_ASAP7_75t_L g7176 ( 
.A(n_7161),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_7170),
.Y(n_7177)
);

AND2x2_ASAP7_75t_L g7178 ( 
.A(n_7162),
.B(n_750),
.Y(n_7178)
);

NAND2xp5_ASAP7_75t_L g7179 ( 
.A(n_7114),
.B(n_750),
.Y(n_7179)
);

OAI21xp33_ASAP7_75t_L g7180 ( 
.A1(n_7091),
.A2(n_750),
.B(n_751),
.Y(n_7180)
);

OAI32xp33_ASAP7_75t_L g7181 ( 
.A1(n_7092),
.A2(n_753),
.A3(n_751),
.B1(n_752),
.B2(n_754),
.Y(n_7181)
);

A2O1A1Ixp33_ASAP7_75t_L g7182 ( 
.A1(n_7121),
.A2(n_7119),
.B(n_7116),
.C(n_7112),
.Y(n_7182)
);

AOI22xp5_ASAP7_75t_L g7183 ( 
.A1(n_7108),
.A2(n_755),
.B1(n_753),
.B2(n_754),
.Y(n_7183)
);

OAI221xp5_ASAP7_75t_L g7184 ( 
.A1(n_7144),
.A2(n_7128),
.B1(n_7138),
.B2(n_7102),
.C(n_7156),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_7096),
.Y(n_7185)
);

AND2x2_ASAP7_75t_L g7186 ( 
.A(n_7159),
.B(n_753),
.Y(n_7186)
);

OAI22xp33_ASAP7_75t_L g7187 ( 
.A1(n_7133),
.A2(n_758),
.B1(n_755),
.B2(n_756),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_L g7188 ( 
.A(n_7164),
.B(n_755),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_7098),
.Y(n_7189)
);

AOI221xp5_ASAP7_75t_L g7190 ( 
.A1(n_7166),
.A2(n_759),
.B1(n_756),
.B2(n_758),
.C(n_760),
.Y(n_7190)
);

AOI22xp33_ASAP7_75t_L g7191 ( 
.A1(n_7137),
.A2(n_760),
.B1(n_756),
.B2(n_759),
.Y(n_7191)
);

NAND2xp5_ASAP7_75t_L g7192 ( 
.A(n_7168),
.B(n_762),
.Y(n_7192)
);

OR2x2_ASAP7_75t_L g7193 ( 
.A(n_7169),
.B(n_762),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_7140),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_7124),
.Y(n_7195)
);

O2A1O1Ixp5_ASAP7_75t_L g7196 ( 
.A1(n_7132),
.A2(n_764),
.B(n_762),
.C(n_763),
.Y(n_7196)
);

AOI21xp5_ASAP7_75t_L g7197 ( 
.A1(n_7089),
.A2(n_7103),
.B(n_7130),
.Y(n_7197)
);

NOR2xp33_ASAP7_75t_L g7198 ( 
.A(n_7120),
.B(n_7099),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_7095),
.Y(n_7199)
);

AOI21xp5_ASAP7_75t_L g7200 ( 
.A1(n_7141),
.A2(n_763),
.B(n_765),
.Y(n_7200)
);

AND2x2_ASAP7_75t_L g7201 ( 
.A(n_7125),
.B(n_765),
.Y(n_7201)
);

OAI221xp5_ASAP7_75t_L g7202 ( 
.A1(n_7111),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.C(n_769),
.Y(n_7202)
);

INVx2_ASAP7_75t_L g7203 ( 
.A(n_7094),
.Y(n_7203)
);

OAI21xp5_ASAP7_75t_L g7204 ( 
.A1(n_7158),
.A2(n_767),
.B(n_768),
.Y(n_7204)
);

AND2x2_ASAP7_75t_L g7205 ( 
.A(n_7109),
.B(n_7129),
.Y(n_7205)
);

NAND3xp33_ASAP7_75t_L g7206 ( 
.A(n_7165),
.B(n_768),
.C(n_769),
.Y(n_7206)
);

INVx1_ASAP7_75t_L g7207 ( 
.A(n_7139),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_7160),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_7150),
.Y(n_7209)
);

OR2x2_ASAP7_75t_L g7210 ( 
.A(n_7189),
.B(n_7142),
.Y(n_7210)
);

NAND2xp5_ASAP7_75t_L g7211 ( 
.A(n_7173),
.B(n_7167),
.Y(n_7211)
);

OAI21xp5_ASAP7_75t_L g7212 ( 
.A1(n_7197),
.A2(n_7157),
.B(n_7106),
.Y(n_7212)
);

HB1xp67_ASAP7_75t_L g7213 ( 
.A(n_7176),
.Y(n_7213)
);

NAND3xp33_ASAP7_75t_L g7214 ( 
.A(n_7191),
.B(n_7122),
.C(n_7101),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_7178),
.Y(n_7215)
);

INVx1_ASAP7_75t_L g7216 ( 
.A(n_7186),
.Y(n_7216)
);

AND2x2_ASAP7_75t_L g7217 ( 
.A(n_7205),
.B(n_7110),
.Y(n_7217)
);

NOR2xp33_ASAP7_75t_L g7218 ( 
.A(n_7199),
.B(n_7090),
.Y(n_7218)
);

INVx3_ASAP7_75t_SL g7219 ( 
.A(n_7203),
.Y(n_7219)
);

INVx1_ASAP7_75t_L g7220 ( 
.A(n_7179),
.Y(n_7220)
);

AND2x2_ASAP7_75t_L g7221 ( 
.A(n_7201),
.B(n_7088),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_7171),
.Y(n_7222)
);

OR2x2_ASAP7_75t_L g7223 ( 
.A(n_7185),
.B(n_7100),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_7172),
.Y(n_7224)
);

INVx1_ASAP7_75t_SL g7225 ( 
.A(n_7193),
.Y(n_7225)
);

AND2x2_ASAP7_75t_L g7226 ( 
.A(n_7174),
.B(n_7107),
.Y(n_7226)
);

AND2x2_ASAP7_75t_L g7227 ( 
.A(n_7198),
.B(n_7131),
.Y(n_7227)
);

INVx2_ASAP7_75t_L g7228 ( 
.A(n_7208),
.Y(n_7228)
);

INVx1_ASAP7_75t_SL g7229 ( 
.A(n_7188),
.Y(n_7229)
);

OR2x6_ASAP7_75t_L g7230 ( 
.A(n_7200),
.B(n_7152),
.Y(n_7230)
);

NOR2xp33_ASAP7_75t_L g7231 ( 
.A(n_7180),
.B(n_7093),
.Y(n_7231)
);

NOR2xp33_ASAP7_75t_L g7232 ( 
.A(n_7192),
.B(n_7147),
.Y(n_7232)
);

NAND2xp5_ASAP7_75t_L g7233 ( 
.A(n_7183),
.B(n_7117),
.Y(n_7233)
);

INVx1_ASAP7_75t_L g7234 ( 
.A(n_7183),
.Y(n_7234)
);

NOR2xp33_ASAP7_75t_L g7235 ( 
.A(n_7184),
.B(n_7151),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_7181),
.Y(n_7236)
);

INVx2_ASAP7_75t_L g7237 ( 
.A(n_7209),
.Y(n_7237)
);

OR2x2_ASAP7_75t_L g7238 ( 
.A(n_7182),
.B(n_7134),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7194),
.B(n_7149),
.Y(n_7239)
);

NAND2xp5_ASAP7_75t_L g7240 ( 
.A(n_7190),
.B(n_7187),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_7202),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_7175),
.B(n_7126),
.Y(n_7242)
);

NOR2x1_ASAP7_75t_L g7243 ( 
.A(n_7206),
.B(n_7123),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_7196),
.Y(n_7244)
);

NOR2xp33_ASAP7_75t_L g7245 ( 
.A(n_7177),
.B(n_7113),
.Y(n_7245)
);

NAND2xp5_ASAP7_75t_L g7246 ( 
.A(n_7207),
.B(n_7126),
.Y(n_7246)
);

OR2x2_ASAP7_75t_L g7247 ( 
.A(n_7204),
.B(n_7148),
.Y(n_7247)
);

HB1xp67_ASAP7_75t_L g7248 ( 
.A(n_7195),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_7189),
.Y(n_7249)
);

NAND2xp5_ASAP7_75t_L g7250 ( 
.A(n_7189),
.B(n_7136),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_L g7251 ( 
.A(n_7189),
.B(n_7145),
.Y(n_7251)
);

NAND2xp5_ASAP7_75t_L g7252 ( 
.A(n_7189),
.B(n_7118),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_7189),
.Y(n_7253)
);

AND2x2_ASAP7_75t_L g7254 ( 
.A(n_7189),
.B(n_7143),
.Y(n_7254)
);

AND2x2_ASAP7_75t_L g7255 ( 
.A(n_7217),
.B(n_7104),
.Y(n_7255)
);

NAND3xp33_ASAP7_75t_L g7256 ( 
.A(n_7218),
.B(n_7153),
.C(n_7155),
.Y(n_7256)
);

AOI21xp33_ASAP7_75t_L g7257 ( 
.A1(n_7210),
.A2(n_7146),
.B(n_7135),
.Y(n_7257)
);

NOR2xp67_ASAP7_75t_L g7258 ( 
.A(n_7214),
.B(n_7115),
.Y(n_7258)
);

A2O1A1Ixp33_ASAP7_75t_L g7259 ( 
.A1(n_7235),
.A2(n_771),
.B(n_769),
.C(n_770),
.Y(n_7259)
);

INVx1_ASAP7_75t_L g7260 ( 
.A(n_7213),
.Y(n_7260)
);

NAND4xp25_ASAP7_75t_L g7261 ( 
.A(n_7251),
.B(n_772),
.C(n_770),
.D(n_771),
.Y(n_7261)
);

NAND4xp25_ASAP7_75t_L g7262 ( 
.A(n_7231),
.B(n_772),
.C(n_770),
.D(n_771),
.Y(n_7262)
);

NAND3xp33_ASAP7_75t_SL g7263 ( 
.A(n_7212),
.B(n_772),
.C(n_773),
.Y(n_7263)
);

NOR3xp33_ASAP7_75t_L g7264 ( 
.A(n_7249),
.B(n_773),
.C(n_774),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_7253),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_7238),
.Y(n_7266)
);

AOI21xp33_ASAP7_75t_L g7267 ( 
.A1(n_7223),
.A2(n_773),
.B(n_774),
.Y(n_7267)
);

INVx1_ASAP7_75t_L g7268 ( 
.A(n_7227),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7252),
.Y(n_7269)
);

AO22x1_ASAP7_75t_SL g7270 ( 
.A1(n_7219),
.A2(n_777),
.B1(n_775),
.B2(n_776),
.Y(n_7270)
);

NOR2xp67_ASAP7_75t_L g7271 ( 
.A(n_7244),
.B(n_775),
.Y(n_7271)
);

NAND2xp5_ASAP7_75t_L g7272 ( 
.A(n_7236),
.B(n_775),
.Y(n_7272)
);

INVx1_ASAP7_75t_L g7273 ( 
.A(n_7211),
.Y(n_7273)
);

NAND3xp33_ASAP7_75t_L g7274 ( 
.A(n_7241),
.B(n_776),
.C(n_777),
.Y(n_7274)
);

INVx1_ASAP7_75t_L g7275 ( 
.A(n_7254),
.Y(n_7275)
);

NAND2xp5_ASAP7_75t_L g7276 ( 
.A(n_7234),
.B(n_776),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_SL g7277 ( 
.A(n_7228),
.B(n_7250),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_7226),
.Y(n_7278)
);

NOR4xp25_ASAP7_75t_L g7279 ( 
.A(n_7225),
.B(n_779),
.C(n_777),
.D(n_778),
.Y(n_7279)
);

NAND2xp5_ASAP7_75t_SL g7280 ( 
.A(n_7237),
.B(n_778),
.Y(n_7280)
);

NAND4xp75_ASAP7_75t_L g7281 ( 
.A(n_7243),
.B(n_7233),
.C(n_7239),
.D(n_7221),
.Y(n_7281)
);

NAND2xp5_ASAP7_75t_L g7282 ( 
.A(n_7215),
.B(n_779),
.Y(n_7282)
);

NAND3xp33_ASAP7_75t_L g7283 ( 
.A(n_7245),
.B(n_779),
.C(n_780),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_7230),
.Y(n_7284)
);

NAND5xp2_ASAP7_75t_L g7285 ( 
.A(n_7232),
.B(n_782),
.C(n_780),
.D(n_781),
.E(n_783),
.Y(n_7285)
);

NOR2xp33_ASAP7_75t_L g7286 ( 
.A(n_7260),
.B(n_7216),
.Y(n_7286)
);

AOI21xp5_ASAP7_75t_L g7287 ( 
.A1(n_7272),
.A2(n_7240),
.B(n_7242),
.Y(n_7287)
);

INVx1_ASAP7_75t_SL g7288 ( 
.A(n_7255),
.Y(n_7288)
);

AOI211xp5_ASAP7_75t_L g7289 ( 
.A1(n_7267),
.A2(n_7229),
.B(n_7248),
.C(n_7222),
.Y(n_7289)
);

NOR2x1_ASAP7_75t_L g7290 ( 
.A(n_7274),
.B(n_7230),
.Y(n_7290)
);

NAND2xp5_ASAP7_75t_L g7291 ( 
.A(n_7258),
.B(n_7220),
.Y(n_7291)
);

INVx1_ASAP7_75t_L g7292 ( 
.A(n_7270),
.Y(n_7292)
);

INVx1_ASAP7_75t_L g7293 ( 
.A(n_7276),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_7271),
.Y(n_7294)
);

BUFx2_ASAP7_75t_L g7295 ( 
.A(n_7275),
.Y(n_7295)
);

OAI211xp5_ASAP7_75t_SL g7296 ( 
.A1(n_7257),
.A2(n_7246),
.B(n_7224),
.C(n_7247),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_7282),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_7278),
.Y(n_7298)
);

OR2x2_ASAP7_75t_L g7299 ( 
.A(n_7261),
.B(n_780),
.Y(n_7299)
);

AND3x1_ASAP7_75t_L g7300 ( 
.A(n_7285),
.B(n_781),
.C(n_782),
.Y(n_7300)
);

BUFx2_ASAP7_75t_L g7301 ( 
.A(n_7268),
.Y(n_7301)
);

AND3x1_ASAP7_75t_L g7302 ( 
.A(n_7264),
.B(n_781),
.C(n_782),
.Y(n_7302)
);

NAND2xp5_ASAP7_75t_SL g7303 ( 
.A(n_7266),
.B(n_783),
.Y(n_7303)
);

NOR3xp33_ASAP7_75t_L g7304 ( 
.A(n_7263),
.B(n_783),
.C(n_784),
.Y(n_7304)
);

AND2x2_ASAP7_75t_L g7305 ( 
.A(n_7265),
.B(n_785),
.Y(n_7305)
);

NAND2xp5_ASAP7_75t_L g7306 ( 
.A(n_7259),
.B(n_785),
.Y(n_7306)
);

NAND2xp5_ASAP7_75t_L g7307 ( 
.A(n_7279),
.B(n_785),
.Y(n_7307)
);

NAND2xp5_ASAP7_75t_L g7308 ( 
.A(n_7284),
.B(n_786),
.Y(n_7308)
);

NOR2xp33_ASAP7_75t_L g7309 ( 
.A(n_7281),
.B(n_786),
.Y(n_7309)
);

AOI22xp5_ASAP7_75t_L g7310 ( 
.A1(n_7273),
.A2(n_788),
.B1(n_786),
.B2(n_787),
.Y(n_7310)
);

INVx3_ASAP7_75t_L g7311 ( 
.A(n_7269),
.Y(n_7311)
);

NAND4xp75_ASAP7_75t_L g7312 ( 
.A(n_7277),
.B(n_789),
.C(n_787),
.D(n_788),
.Y(n_7312)
);

OAI22xp5_ASAP7_75t_L g7313 ( 
.A1(n_7256),
.A2(n_792),
.B1(n_789),
.B2(n_790),
.Y(n_7313)
);

NOR2x1_ASAP7_75t_L g7314 ( 
.A(n_7280),
.B(n_789),
.Y(n_7314)
);

OAI22xp5_ASAP7_75t_L g7315 ( 
.A1(n_7283),
.A2(n_793),
.B1(n_790),
.B2(n_792),
.Y(n_7315)
);

AOI21xp5_ASAP7_75t_L g7316 ( 
.A1(n_7262),
.A2(n_792),
.B(n_793),
.Y(n_7316)
);

AOI221xp5_ASAP7_75t_L g7317 ( 
.A1(n_7267),
.A2(n_795),
.B1(n_793),
.B2(n_794),
.C(n_796),
.Y(n_7317)
);

NAND3xp33_ASAP7_75t_SL g7318 ( 
.A(n_7264),
.B(n_794),
.C(n_795),
.Y(n_7318)
);

NAND4xp25_ASAP7_75t_L g7319 ( 
.A(n_7258),
.B(n_797),
.C(n_794),
.D(n_796),
.Y(n_7319)
);

INVx2_ASAP7_75t_L g7320 ( 
.A(n_7255),
.Y(n_7320)
);

INVx2_ASAP7_75t_L g7321 ( 
.A(n_7255),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_7270),
.Y(n_7322)
);

OAI211xp5_ASAP7_75t_SL g7323 ( 
.A1(n_7267),
.A2(n_799),
.B(n_797),
.C(n_798),
.Y(n_7323)
);

AND2x2_ASAP7_75t_L g7324 ( 
.A(n_7255),
.B(n_797),
.Y(n_7324)
);

OAI31xp33_ASAP7_75t_L g7325 ( 
.A1(n_7313),
.A2(n_800),
.A3(n_798),
.B(n_799),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_7311),
.Y(n_7326)
);

INVx2_ASAP7_75t_L g7327 ( 
.A(n_7311),
.Y(n_7327)
);

NOR3xp33_ASAP7_75t_L g7328 ( 
.A(n_7296),
.B(n_798),
.C(n_799),
.Y(n_7328)
);

XOR2xp5_ASAP7_75t_L g7329 ( 
.A(n_7320),
.B(n_800),
.Y(n_7329)
);

AOI22xp33_ASAP7_75t_L g7330 ( 
.A1(n_7309),
.A2(n_802),
.B1(n_800),
.B2(n_801),
.Y(n_7330)
);

NOR3x1_ASAP7_75t_L g7331 ( 
.A(n_7295),
.B(n_801),
.C(n_802),
.Y(n_7331)
);

AOI22xp5_ASAP7_75t_SL g7332 ( 
.A1(n_7305),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_7332)
);

NAND3xp33_ASAP7_75t_L g7333 ( 
.A(n_7317),
.B(n_7304),
.C(n_7319),
.Y(n_7333)
);

AOI22xp33_ASAP7_75t_SL g7334 ( 
.A1(n_7288),
.A2(n_805),
.B1(n_803),
.B2(n_804),
.Y(n_7334)
);

NAND2xp5_ASAP7_75t_L g7335 ( 
.A(n_7321),
.B(n_803),
.Y(n_7335)
);

OAI21xp33_ASAP7_75t_L g7336 ( 
.A1(n_7286),
.A2(n_804),
.B(n_805),
.Y(n_7336)
);

AOI22xp5_ASAP7_75t_L g7337 ( 
.A1(n_7298),
.A2(n_807),
.B1(n_805),
.B2(n_806),
.Y(n_7337)
);

NAND2xp5_ASAP7_75t_SL g7338 ( 
.A(n_7308),
.B(n_806),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_7324),
.Y(n_7339)
);

OAI221xp5_ASAP7_75t_L g7340 ( 
.A1(n_7310),
.A2(n_7307),
.B1(n_7299),
.B2(n_7316),
.C(n_7306),
.Y(n_7340)
);

INVxp67_ASAP7_75t_L g7341 ( 
.A(n_7301),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7312),
.B(n_7315),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_7300),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_7303),
.Y(n_7344)
);

NAND2xp5_ASAP7_75t_L g7345 ( 
.A(n_7287),
.B(n_806),
.Y(n_7345)
);

AO22x2_ASAP7_75t_L g7346 ( 
.A1(n_7292),
.A2(n_809),
.B1(n_807),
.B2(n_808),
.Y(n_7346)
);

BUFx24_ASAP7_75t_SL g7347 ( 
.A(n_7289),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_7302),
.Y(n_7348)
);

AOI32xp33_ASAP7_75t_L g7349 ( 
.A1(n_7323),
.A2(n_809),
.A3(n_807),
.B1(n_808),
.B2(n_810),
.Y(n_7349)
);

AOI322xp5_ASAP7_75t_L g7350 ( 
.A1(n_7290),
.A2(n_809),
.A3(n_810),
.B1(n_811),
.B2(n_812),
.C1(n_813),
.C2(n_814),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_L g7351 ( 
.A(n_7322),
.B(n_810),
.Y(n_7351)
);

AOI211xp5_ASAP7_75t_L g7352 ( 
.A1(n_7318),
.A2(n_813),
.B(n_811),
.C(n_812),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_7291),
.Y(n_7353)
);

INVxp67_ASAP7_75t_L g7354 ( 
.A(n_7314),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_L g7355 ( 
.A(n_7293),
.B(n_811),
.Y(n_7355)
);

NAND2xp5_ASAP7_75t_L g7356 ( 
.A(n_7350),
.B(n_7297),
.Y(n_7356)
);

AO22x2_ASAP7_75t_L g7357 ( 
.A1(n_7347),
.A2(n_7294),
.B1(n_814),
.B2(n_812),
.Y(n_7357)
);

NAND4xp25_ASAP7_75t_L g7358 ( 
.A(n_7353),
.B(n_815),
.C(n_813),
.D(n_814),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_7346),
.Y(n_7359)
);

NAND3xp33_ASAP7_75t_L g7360 ( 
.A(n_7328),
.B(n_815),
.C(n_816),
.Y(n_7360)
);

OAI22xp5_ASAP7_75t_SL g7361 ( 
.A1(n_7329),
.A2(n_819),
.B1(n_817),
.B2(n_818),
.Y(n_7361)
);

INVx2_ASAP7_75t_L g7362 ( 
.A(n_7326),
.Y(n_7362)
);

A2O1A1Ixp33_ASAP7_75t_SL g7363 ( 
.A1(n_7341),
.A2(n_819),
.B(n_817),
.C(n_818),
.Y(n_7363)
);

O2A1O1Ixp33_ASAP7_75t_L g7364 ( 
.A1(n_7351),
.A2(n_819),
.B(n_817),
.C(n_818),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_7346),
.Y(n_7365)
);

NAND2xp5_ASAP7_75t_L g7366 ( 
.A(n_7334),
.B(n_7327),
.Y(n_7366)
);

AOI221xp5_ASAP7_75t_L g7367 ( 
.A1(n_7336),
.A2(n_823),
.B1(n_820),
.B2(n_822),
.C(n_824),
.Y(n_7367)
);

AOI22xp5_ASAP7_75t_L g7368 ( 
.A1(n_7343),
.A2(n_823),
.B1(n_820),
.B2(n_822),
.Y(n_7368)
);

OA22x2_ASAP7_75t_L g7369 ( 
.A1(n_7335),
.A2(n_824),
.B1(n_822),
.B2(n_823),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_7337),
.Y(n_7370)
);

OAI22xp33_ASAP7_75t_SL g7371 ( 
.A1(n_7355),
.A2(n_826),
.B1(n_824),
.B2(n_825),
.Y(n_7371)
);

NAND2xp5_ASAP7_75t_SL g7372 ( 
.A(n_7345),
.B(n_825),
.Y(n_7372)
);

BUFx2_ASAP7_75t_L g7373 ( 
.A(n_7339),
.Y(n_7373)
);

AOI22xp5_ASAP7_75t_L g7374 ( 
.A1(n_7348),
.A2(n_828),
.B1(n_826),
.B2(n_827),
.Y(n_7374)
);

AOI22xp5_ASAP7_75t_L g7375 ( 
.A1(n_7333),
.A2(n_829),
.B1(n_826),
.B2(n_828),
.Y(n_7375)
);

OAI22xp5_ASAP7_75t_L g7376 ( 
.A1(n_7340),
.A2(n_831),
.B1(n_829),
.B2(n_830),
.Y(n_7376)
);

NAND2xp5_ASAP7_75t_SL g7377 ( 
.A(n_7325),
.B(n_829),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_7332),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_7330),
.B(n_7352),
.Y(n_7379)
);

INVx1_ASAP7_75t_L g7380 ( 
.A(n_7331),
.Y(n_7380)
);

NOR2xp33_ASAP7_75t_L g7381 ( 
.A(n_7373),
.B(n_7354),
.Y(n_7381)
);

OAI221xp5_ASAP7_75t_L g7382 ( 
.A1(n_7362),
.A2(n_7349),
.B1(n_7342),
.B2(n_7338),
.C(n_7344),
.Y(n_7382)
);

INVx2_ASAP7_75t_L g7383 ( 
.A(n_7369),
.Y(n_7383)
);

NAND2xp5_ASAP7_75t_L g7384 ( 
.A(n_7375),
.B(n_7368),
.Y(n_7384)
);

NOR2x1_ASAP7_75t_L g7385 ( 
.A(n_7359),
.B(n_830),
.Y(n_7385)
);

NOR2x1_ASAP7_75t_L g7386 ( 
.A(n_7365),
.B(n_830),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_7357),
.Y(n_7387)
);

INVxp67_ASAP7_75t_L g7388 ( 
.A(n_7357),
.Y(n_7388)
);

AND2x2_ASAP7_75t_L g7389 ( 
.A(n_7380),
.B(n_831),
.Y(n_7389)
);

OAI22xp5_ASAP7_75t_L g7390 ( 
.A1(n_7378),
.A2(n_833),
.B1(n_831),
.B2(n_832),
.Y(n_7390)
);

NOR2x1_ASAP7_75t_L g7391 ( 
.A(n_7360),
.B(n_832),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_7361),
.Y(n_7392)
);

NAND2xp5_ASAP7_75t_L g7393 ( 
.A(n_7374),
.B(n_833),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_7376),
.B(n_834),
.Y(n_7394)
);

NOR2x1_ASAP7_75t_L g7395 ( 
.A(n_7356),
.B(n_834),
.Y(n_7395)
);

NAND3x1_ASAP7_75t_SL g7396 ( 
.A(n_7367),
.B(n_835),
.C(n_836),
.Y(n_7396)
);

XNOR2xp5_ASAP7_75t_L g7397 ( 
.A(n_7358),
.B(n_835),
.Y(n_7397)
);

NAND3xp33_ASAP7_75t_L g7398 ( 
.A(n_7364),
.B(n_835),
.C(n_837),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_7371),
.Y(n_7399)
);

NOR3xp33_ASAP7_75t_SL g7400 ( 
.A(n_7382),
.B(n_7381),
.C(n_7366),
.Y(n_7400)
);

NOR3xp33_ASAP7_75t_L g7401 ( 
.A(n_7399),
.B(n_7379),
.C(n_7377),
.Y(n_7401)
);

NAND3xp33_ASAP7_75t_SL g7402 ( 
.A(n_7384),
.B(n_7370),
.C(n_7372),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_7385),
.Y(n_7403)
);

NAND3xp33_ASAP7_75t_SL g7404 ( 
.A(n_7389),
.B(n_7363),
.C(n_837),
.Y(n_7404)
);

NOR2x1_ASAP7_75t_L g7405 ( 
.A(n_7395),
.B(n_970),
.Y(n_7405)
);

NAND3xp33_ASAP7_75t_L g7406 ( 
.A(n_7397),
.B(n_837),
.C(n_838),
.Y(n_7406)
);

INVx2_ASAP7_75t_SL g7407 ( 
.A(n_7383),
.Y(n_7407)
);

NOR3xp33_ASAP7_75t_L g7408 ( 
.A(n_7392),
.B(n_972),
.C(n_971),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_L g7409 ( 
.A(n_7400),
.B(n_7388),
.Y(n_7409)
);

NOR2xp67_ASAP7_75t_L g7410 ( 
.A(n_7402),
.B(n_7387),
.Y(n_7410)
);

NOR2xp33_ASAP7_75t_L g7411 ( 
.A(n_7404),
.B(n_7394),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_7409),
.Y(n_7412)
);

INVx2_ASAP7_75t_L g7413 ( 
.A(n_7411),
.Y(n_7413)
);

OR3x1_ASAP7_75t_L g7414 ( 
.A(n_7412),
.B(n_7403),
.C(n_7401),
.Y(n_7414)
);

BUFx2_ASAP7_75t_L g7415 ( 
.A(n_7413),
.Y(n_7415)
);

AOI22xp5_ASAP7_75t_L g7416 ( 
.A1(n_7414),
.A2(n_7407),
.B1(n_7410),
.B2(n_7393),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7415),
.Y(n_7417)
);

NAND2xp5_ASAP7_75t_L g7418 ( 
.A(n_7417),
.B(n_7386),
.Y(n_7418)
);

HB1xp67_ASAP7_75t_L g7419 ( 
.A(n_7416),
.Y(n_7419)
);

INVxp67_ASAP7_75t_SL g7420 ( 
.A(n_7419),
.Y(n_7420)
);

INVx2_ASAP7_75t_L g7421 ( 
.A(n_7420),
.Y(n_7421)
);

OAI21xp5_ASAP7_75t_L g7422 ( 
.A1(n_7421),
.A2(n_7418),
.B(n_7391),
.Y(n_7422)
);

BUFx2_ASAP7_75t_L g7423 ( 
.A(n_7422),
.Y(n_7423)
);

AOI22xp5_ASAP7_75t_L g7424 ( 
.A1(n_7423),
.A2(n_7405),
.B1(n_7406),
.B2(n_7408),
.Y(n_7424)
);

OAI222xp33_ASAP7_75t_L g7425 ( 
.A1(n_7424),
.A2(n_7390),
.B1(n_7396),
.B2(n_7398),
.C1(n_1031),
.C2(n_1030),
.Y(n_7425)
);

BUFx24_ASAP7_75t_SL g7426 ( 
.A(n_7425),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_7426),
.Y(n_7427)
);

OAI221xp5_ASAP7_75t_L g7428 ( 
.A1(n_7427),
.A2(n_974),
.B1(n_975),
.B2(n_972),
.C(n_971),
.Y(n_7428)
);

AOI22xp5_ASAP7_75t_L g7429 ( 
.A1(n_7428),
.A2(n_840),
.B1(n_838),
.B2(n_839),
.Y(n_7429)
);

AOI211xp5_ASAP7_75t_L g7430 ( 
.A1(n_7429),
.A2(n_841),
.B(n_839),
.C(n_840),
.Y(n_7430)
);


endmodule