module fake_jpeg_1232_n_535 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_50),
.B(n_95),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_57),
.Y(n_137)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_13),
.B(n_12),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_59),
.A2(n_44),
.B(n_29),
.C(n_26),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_61),
.Y(n_140)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_83),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_SL g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_80),
.A2(n_32),
.B1(n_21),
.B2(n_36),
.Y(n_153)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_34),
.B(n_11),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_43),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_16),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

BUFx12f_ASAP7_75t_SL g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_20),
.Y(n_94)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_22),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_102),
.B(n_119),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_107),
.A2(n_114),
.B1(n_108),
.B2(n_110),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_108),
.A2(n_110),
.B1(n_114),
.B2(n_134),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_28),
.B1(n_45),
.B2(n_33),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_109),
.A2(n_153),
.B1(n_17),
.B2(n_64),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_44),
.B1(n_45),
.B2(n_22),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_132),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_33),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_70),
.A2(n_38),
.B1(n_32),
.B2(n_21),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_38),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_42),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_80),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_58),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_85),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_52),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_180),
.Y(n_218)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_92),
.C(n_91),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_190),
.C(n_127),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_77),
.B1(n_53),
.B2(n_66),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_186),
.B1(n_196),
.B2(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_57),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_185),
.Y(n_211)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_183),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_184),
.A2(n_195),
.B(n_145),
.Y(n_237)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_105),
.A2(n_96),
.B1(n_75),
.B2(n_79),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_73),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_191),
.Y(n_234)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_65),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_123),
.B(n_42),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_134),
.A2(n_78),
.B1(n_86),
.B2(n_60),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_192),
.A2(n_201),
.B1(n_204),
.B2(n_118),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_39),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_197),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_54),
.B1(n_72),
.B2(n_88),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_152),
.A2(n_39),
.B1(n_17),
.B2(n_36),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_156),
.Y(n_197)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_140),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_101),
.A2(n_63),
.B1(n_56),
.B2(n_55),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_135),
.A2(n_17),
.B1(n_76),
.B2(n_71),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_138),
.B1(n_125),
.B2(n_144),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_157),
.B1(n_118),
.B2(n_124),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_210),
.A2(n_225),
.B1(n_183),
.B2(n_170),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_163),
.C(n_165),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_226),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_136),
.B1(n_157),
.B2(n_122),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_150),
.B1(n_125),
.B2(n_144),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_101),
.B1(n_147),
.B2(n_143),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_206),
.B1(n_159),
.B2(n_168),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_155),
.B1(n_99),
.B2(n_121),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx11_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_251),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_237),
.B(n_205),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_212),
.B(n_219),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_198),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_202),
.B1(n_191),
.B2(n_195),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_253),
.A2(n_259),
.B1(n_274),
.B2(n_239),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_180),
.B(n_187),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_254),
.A2(n_171),
.B(n_215),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_225),
.B1(n_214),
.B2(n_240),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_178),
.B1(n_190),
.B2(n_161),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_212),
.B1(n_226),
.B2(n_241),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_124),
.B1(n_122),
.B2(n_136),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_189),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_262),
.Y(n_296)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_175),
.Y(n_262)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_210),
.B1(n_221),
.B2(n_236),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_264),
.A2(n_176),
.B(n_209),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_209),
.Y(n_266)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_177),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_276),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_234),
.B(n_181),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_275),
.Y(n_293)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_218),
.A2(n_208),
.B1(n_173),
.B2(n_190),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_213),
.B(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_230),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_228),
.B1(n_226),
.B2(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_282),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_283),
.A2(n_290),
.B1(n_300),
.B2(n_307),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_268),
.B(n_250),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_226),
.C(n_242),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_289),
.C(n_292),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_242),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_216),
.B1(n_244),
.B2(n_235),
.Y(n_290)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_241),
.A3(n_229),
.B1(n_232),
.B2(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_185),
.C(n_220),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_159),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_220),
.C(n_188),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_258),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_265),
.A2(n_216),
.B(n_200),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_262),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_251),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_265),
.A2(n_227),
.B1(n_160),
.B2(n_167),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_215),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_278),
.Y(n_312)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_315),
.A2(n_319),
.B(n_335),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_318),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_260),
.Y(n_317)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_294),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_268),
.B(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_247),
.Y(n_320)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_299),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_324),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_286),
.A2(n_252),
.B(n_268),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_325),
.A2(n_319),
.B(n_315),
.Y(n_377)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_282),
.A2(n_257),
.B1(n_269),
.B2(n_270),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_327),
.A2(n_344),
.B1(n_266),
.B2(n_209),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_SL g328 ( 
.A(n_290),
.B(n_253),
.C(n_270),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_328),
.B(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_254),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_333),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_332),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_310),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_264),
.B(n_270),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_254),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_272),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_302),
.A2(n_258),
.B1(n_256),
.B2(n_248),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_287),
.B1(n_289),
.B2(n_303),
.Y(n_349)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_341),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_276),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_339),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_279),
.B(n_246),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_279),
.A2(n_256),
.B1(n_267),
.B2(n_259),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_349),
.A2(n_350),
.B1(n_359),
.B2(n_367),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_311),
.A2(n_300),
.B1(n_302),
.B2(n_307),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_341),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_352),
.B(n_329),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_353),
.A2(n_231),
.B(n_174),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_284),
.C(n_292),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_323),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_309),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_366),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_335),
.A2(n_297),
.B1(n_300),
.B2(n_284),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_358),
.A2(n_365),
.B1(n_339),
.B2(n_325),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_311),
.A2(n_297),
.B1(n_263),
.B2(n_291),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_363),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_285),
.B1(n_305),
.B2(n_299),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_337),
.B(n_274),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_314),
.A2(n_285),
.B1(n_305),
.B2(n_266),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_266),
.B1(n_261),
.B2(n_277),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_369),
.A2(n_376),
.B1(n_324),
.B2(n_332),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_371),
.A2(n_377),
.B(n_312),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_326),
.B(n_232),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_372),
.B(n_150),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_231),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_314),
.A2(n_277),
.B1(n_261),
.B2(n_227),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_374),
.A2(n_321),
.B1(n_340),
.B2(n_313),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_338),
.Y(n_375)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_334),
.A2(n_227),
.B1(n_217),
.B2(n_222),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_378),
.A2(n_403),
.B1(n_374),
.B2(n_364),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_345),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_397),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_380),
.B(n_364),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_336),
.B1(n_317),
.B2(n_320),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_387),
.B1(n_394),
.B2(n_399),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_333),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_384),
.B(n_393),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_357),
.C(n_373),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_402),
.C(n_366),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_331),
.Y(n_388)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g389 ( 
.A(n_358),
.B(n_328),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_389),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_346),
.Y(n_391)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_316),
.Y(n_393)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_396),
.Y(n_435)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_351),
.B(n_332),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_405),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_359),
.A2(n_329),
.B1(n_199),
.B2(n_166),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_406),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_117),
.C(n_126),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_360),
.B1(n_367),
.B2(n_351),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_404),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_355),
.B(n_0),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_377),
.A2(n_231),
.B(n_174),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_362),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_356),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_433),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_427),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_SL g412 ( 
.A(n_380),
.B(n_360),
.Y(n_412)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_354),
.C(n_365),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_421),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_386),
.A2(n_354),
.B1(n_371),
.B2(n_350),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_419),
.A2(n_429),
.B1(n_401),
.B2(n_398),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_408),
.B(n_370),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_423),
.B(n_426),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_388),
.B(n_362),
.CI(n_347),
.CON(n_426),
.SN(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_382),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_431),
.B(n_395),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_89),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_97),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_378),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_411),
.A2(n_386),
.B1(n_403),
.B2(n_399),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_437),
.A2(n_440),
.B1(n_138),
.B2(n_87),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_435),
.B(n_408),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_442),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_451),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_428),
.A2(n_379),
.B1(n_401),
.B2(n_392),
.Y(n_440)
);

AOI21xp33_ASAP7_75t_L g442 ( 
.A1(n_416),
.A2(n_406),
.B(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_445),
.Y(n_476)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_389),
.C(n_387),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_391),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_448),
.B(n_455),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_415),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_456),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_431),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_25),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_453),
.A2(n_429),
.B1(n_430),
.B2(n_433),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_432),
.A2(n_389),
.B(n_381),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_426),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_404),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_417),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_405),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_459),
.Y(n_474)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_458),
.B(n_428),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_397),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_469),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_472),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_443),
.B(n_414),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_464),
.B(n_465),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_409),
.C(n_425),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_454),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_446),
.B(n_426),
.CI(n_413),
.CON(n_469),
.SN(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_420),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_470),
.B(n_478),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_441),
.A2(n_423),
.B(n_419),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_471),
.B(n_475),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_434),
.C(n_138),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_477),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_437),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_481),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_457),
.Y(n_481)
);

AOI221xp5_ASAP7_75t_L g482 ( 
.A1(n_468),
.A2(n_450),
.B1(n_440),
.B2(n_451),
.C(n_459),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_472),
.B1(n_466),
.B2(n_469),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_450),
.Y(n_483)
);

AOI21x1_ASAP7_75t_L g506 ( 
.A1(n_483),
.A2(n_478),
.B(n_5),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_439),
.C(n_447),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_495),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_447),
.B1(n_25),
.B2(n_3),
.Y(n_485)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_473),
.B(n_1),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_486),
.B(n_488),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_463),
.A2(n_25),
.B(n_2),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_491),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_474),
.B(n_1),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_3),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_479),
.A2(n_469),
.B(n_470),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_497),
.A2(n_500),
.B(n_505),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_499),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_475),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_466),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_507),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_490),
.B(n_494),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_506),
.A2(n_491),
.B(n_6),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_484),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_4),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_508),
.B(n_5),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_493),
.B(n_4),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_509),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_493),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_516),
.Y(n_522)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_512),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_507),
.A2(n_5),
.B(n_6),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_513),
.A2(n_517),
.B(n_518),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_496),
.B(n_5),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_500),
.B(n_5),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_498),
.C(n_501),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_6),
.Y(n_530)
);

O2A1O1Ixp33_ASAP7_75t_SL g523 ( 
.A1(n_519),
.A2(n_515),
.B(n_514),
.C(n_501),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_523),
.A2(n_524),
.B(n_526),
.Y(n_527)
);

A2O1A1O1Ixp25_ASAP7_75t_L g524 ( 
.A1(n_519),
.A2(n_502),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_511),
.A2(n_10),
.B(n_7),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_522),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_529),
.B(n_530),
.Y(n_531)
);

OAI21xp33_ASAP7_75t_SL g529 ( 
.A1(n_525),
.A2(n_6),
.B(n_7),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_527),
.A2(n_520),
.B(n_8),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_7),
.C(n_9),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_531),
.B(n_10),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_10),
.Y(n_535)
);


endmodule