module fake_jpeg_8137_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.C(n_1),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_37),
.B1(n_44),
.B2(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_92)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_23),
.B1(n_32),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_28),
.B1(n_34),
.B2(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_20),
.B1(n_18),
.B2(n_25),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_44),
.B1(n_35),
.B2(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_62),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_32),
.B1(n_20),
.B2(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_68),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_42),
.B1(n_26),
.B2(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_75),
.B1(n_79),
.B2(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_31),
.B1(n_27),
.B2(n_33),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_17),
.B(n_24),
.C(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_27),
.B1(n_31),
.B2(n_26),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_45),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_69),
.B1(n_67),
.B2(n_53),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_65),
.B1(n_30),
.B2(n_24),
.Y(n_114)
);

NAND2x1_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_41),
.Y(n_85)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_65),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_33),
.B1(n_19),
.B2(n_2),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_46),
.B1(n_52),
.B2(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_68),
.Y(n_99)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_103),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_96),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_100),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_59),
.B1(n_64),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_54),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_110),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_73),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_54),
.C(n_48),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_19),
.B1(n_56),
.B2(n_30),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_24),
.B1(n_9),
.B2(n_2),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_84),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_119),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_85),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_82),
.B(n_86),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_135),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_80),
.B(n_76),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_130),
.B(n_143),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_76),
.B(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_119),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_103),
.B(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_108),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_108),
.B(n_97),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_158),
.B(n_164),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_107),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_152),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_169),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_114),
.B1(n_96),
.B2(n_109),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_167),
.B1(n_128),
.B2(n_135),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_100),
.B(n_112),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_125),
.B1(n_142),
.B2(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_163),
.B1(n_166),
.B2(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_157),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_115),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_104),
.B1(n_79),
.B2(n_75),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_128),
.B(n_123),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_74),
.B1(n_132),
.B2(n_83),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_90),
.B1(n_88),
.B2(n_87),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_168),
.B(n_130),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_88),
.B1(n_87),
.B2(n_91),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_94),
.B1(n_74),
.B2(n_82),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_91),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_86),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_178),
.B(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_124),
.C(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_3),
.C(n_4),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_162),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_124),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_191),
.C(n_196),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_189),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_136),
.B(n_139),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_122),
.B(n_123),
.Y(n_190)
);

NOR4xp25_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_164),
.C(n_157),
.D(n_150),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_146),
.A2(n_132),
.B(n_83),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_165),
.B1(n_159),
.B2(n_167),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_0),
.C(n_1),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_1),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_148),
.C(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_212),
.C(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_206),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_153),
.B1(n_172),
.B2(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_180),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_219),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_147),
.C(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_147),
.C(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_166),
.B1(n_154),
.B2(n_162),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_16),
.C(n_4),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_225),
.Y(n_249)
);

OAI322xp33_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_173),
.A3(n_182),
.B1(n_185),
.B2(n_188),
.C1(n_186),
.C2(n_176),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_193),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_228),
.C(n_235),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_176),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_185),
.B1(n_178),
.B2(n_175),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_204),
.B1(n_218),
.B2(n_205),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_196),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_195),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.C(n_220),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_3),
.C(n_5),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_241),
.Y(n_258)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_209),
.B1(n_207),
.B2(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_233),
.B1(n_210),
.B2(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_219),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_212),
.C(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_3),
.C(n_5),
.Y(n_257)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_253),
.B1(n_6),
.B2(n_7),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_222),
.B(n_216),
.CI(n_214),
.CON(n_253),
.SN(n_253)
);

AOI322xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_230),
.A3(n_235),
.B1(n_234),
.B2(n_228),
.C1(n_238),
.C2(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_254),
.B(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_5),
.C(n_6),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_240),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_263),
.B(n_262),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_249),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_241),
.B1(n_244),
.B2(n_247),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_259),
.B1(n_266),
.B2(n_264),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_281),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_263),
.A3(n_266),
.B1(n_246),
.B2(n_261),
.C1(n_257),
.C2(n_252),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_250),
.B(n_242),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_253),
.C(n_10),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_11),
.B(n_12),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_272),
.B1(n_273),
.B2(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_7),
.C(n_11),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_290),
.A2(n_13),
.B(n_14),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

NOR2x1p5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_15),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_289),
.B(n_286),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_294),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_296),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_16),
.Y(n_299)
);


endmodule