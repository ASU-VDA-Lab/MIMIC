module fake_netlist_5_598_n_2001 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_598, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2001);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_598;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2001;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_1508;
wire n_785;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_1007;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_933;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_1696;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_1230;
wire n_668;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_1016;
wire n_1243;
wire n_1280;
wire n_1845;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_926;
wire n_1218;
wire n_1931;
wire n_1070;
wire n_777;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_1796;
wire n_1473;
wire n_680;
wire n_1587;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_889;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_1819;
wire n_1527;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_832;
wire n_857;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_1775;
wire n_1368;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_1609;
wire n_1989;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_1591;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_860;
wire n_1805;
wire n_1816;
wire n_948;
wire n_1217;
wire n_628;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_602;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_1645;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_885;
wire n_1432;
wire n_1357;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_618;
wire n_896;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_681;
wire n_1638;
wire n_1786;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_1457;
wire n_766;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1999;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_1235;
wire n_703;
wire n_980;
wire n_1115;
wire n_698;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_812;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1995;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_751;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_1842;
wire n_871;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_1937;
wire n_1739;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_401),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_294),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_553),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_555),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_138),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_213),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_306),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_447),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_537),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_551),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_517),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_564),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_122),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_539),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_220),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_503),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_361),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_532),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_336),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_591),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_371),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_593),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_96),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_238),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_421),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_481),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_203),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_24),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_93),
.Y(n_627)
);

CKINVDCx14_ASAP7_75t_R g628 ( 
.A(n_146),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_468),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_171),
.Y(n_630)
);

CKINVDCx16_ASAP7_75t_R g631 ( 
.A(n_262),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_419),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_304),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_31),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_368),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_445),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_406),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_516),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_496),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_183),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_565),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_216),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_256),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_549),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_326),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_563),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_594),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_446),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_206),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_221),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_55),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_330),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_433),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_247),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_103),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_64),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_531),
.Y(n_658)
);

BUFx8_ASAP7_75t_SL g659 ( 
.A(n_126),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_597),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_243),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_75),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_585),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_550),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_509),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_554),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_325),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_515),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_216),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_129),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_530),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_583),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_459),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_106),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_577),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_512),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_274),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_568),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_347),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_561),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_572),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_383),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_289),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_139),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_580),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_359),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_88),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_139),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_470),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_289),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_290),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_535),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_587),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_588),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_558),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_569),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_544),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_584),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_570),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_245),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_430),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_534),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_452),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_356),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_417),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_592),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_510),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_44),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_21),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_525),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_309),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_283),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_183),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_548),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_598),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_483),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_526),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_426),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_76),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_199),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_311),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_76),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_559),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_574),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_61),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_248),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_302),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_414),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_457),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_79),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_533),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_511),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_21),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_536),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_132),
.Y(n_735)
);

BUFx5_ASAP7_75t_L g736 ( 
.A(n_186),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_541),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_78),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_323),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_527),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_519),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_233),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_311),
.Y(n_743)
);

CKINVDCx14_ASAP7_75t_R g744 ( 
.A(n_250),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_10),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_444),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_161),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_478),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_187),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_596),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_384),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_405),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_524),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_477),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_582),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_11),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_514),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_68),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_557),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_165),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_579),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_327),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_199),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_540),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_236),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_365),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_442),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_529),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_408),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_578),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_545),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_239),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_595),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_507),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_538),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_518),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_395),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_364),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_546),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_566),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_175),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_179),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_432),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_390),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_171),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_522),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_571),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_102),
.Y(n_788)
);

INVxp33_ASAP7_75t_R g789 ( 
.A(n_376),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_581),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_355),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_575),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_191),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_294),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_351),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_320),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_590),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_267),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_261),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_145),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_169),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_508),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_12),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_165),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_513),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_521),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_586),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_428),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_450),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_560),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_528),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_181),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_576),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_449),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_486),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_556),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_144),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_11),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_542),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_153),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_475),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_155),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_337),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_523),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_448),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_429),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_543),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_431),
.Y(n_828)
);

BUFx10_ASAP7_75t_L g829 ( 
.A(n_167),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_340),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_275),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_520),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_118),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_562),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_235),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_246),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_257),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_16),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_415),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_480),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_573),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_69),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_552),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_230),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_77),
.Y(n_845)
);

BUFx8_ASAP7_75t_SL g846 ( 
.A(n_332),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_58),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_112),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_505),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_423),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_110),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_589),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_472),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_547),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_17),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_143),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_69),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_285),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_220),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_659),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_749),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_628),
.B(n_0),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_674),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_668),
.B(n_0),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_749),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_736),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_749),
.Y(n_867)
);

INVx5_ASAP7_75t_L g868 ( 
.A(n_676),
.Y(n_868)
);

INVx5_ASAP7_75t_L g869 ( 
.A(n_676),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_744),
.B(n_1),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_724),
.B(n_2),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_781),
.Y(n_872)
);

INVx5_ASAP7_75t_L g873 ( 
.A(n_676),
.Y(n_873)
);

BUFx8_ASAP7_75t_SL g874 ( 
.A(n_846),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_701),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_706),
.B(n_1),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_781),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_631),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_643),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_677),
.B(n_2),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_764),
.B(n_3),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_736),
.Y(n_882)
);

INVx6_ASAP7_75t_L g883 ( 
.A(n_643),
.Y(n_883)
);

BUFx8_ASAP7_75t_SL g884 ( 
.A(n_605),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_599),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_781),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_715),
.B(n_3),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_736),
.B(n_4),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_683),
.Y(n_889)
);

AO22x2_ASAP7_75t_L g890 ( 
.A1(n_864),
.A2(n_798),
.B1(n_604),
.B2(n_634),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_881),
.A2(n_722),
.B1(n_623),
.B2(n_652),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_861),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_871),
.A2(n_666),
.B1(n_689),
.B2(n_620),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_885),
.B(n_639),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_863),
.B(n_644),
.Y(n_895)
);

OAI22xp33_ASAP7_75t_L g896 ( 
.A1(n_862),
.A2(n_837),
.B1(n_649),
.B2(n_711),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_861),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_878),
.A2(n_820),
.B1(n_611),
.B2(n_621),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_870),
.B(n_789),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_879),
.B(n_662),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_880),
.B(n_729),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_865),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_889),
.B(n_821),
.Y(n_903)
);

OAI22xp33_ASAP7_75t_L g904 ( 
.A1(n_876),
.A2(n_735),
.B1(n_738),
.B2(n_733),
.Y(n_904)
);

OAI22xp33_ASAP7_75t_SL g905 ( 
.A1(n_887),
.A2(n_625),
.B1(n_626),
.B2(n_600),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_868),
.B(n_821),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_865),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_868),
.B(n_614),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_860),
.A2(n_704),
.B1(n_826),
.B2(n_697),
.Y(n_909)
);

OAI22xp33_ASAP7_75t_R g910 ( 
.A1(n_884),
.A2(n_848),
.B1(n_613),
.B2(n_657),
.Y(n_910)
);

OAI22xp33_ASAP7_75t_L g911 ( 
.A1(n_888),
.A2(n_630),
.B1(n_633),
.B2(n_627),
.Y(n_911)
);

OAI22xp33_ASAP7_75t_L g912 ( 
.A1(n_883),
.A2(n_642),
.B1(n_651),
.B2(n_640),
.Y(n_912)
);

OA22x2_ASAP7_75t_L g913 ( 
.A1(n_882),
.A2(n_661),
.B1(n_669),
.B2(n_655),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_869),
.B(n_658),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_867),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_873),
.B(n_660),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_875),
.B(n_703),
.Y(n_917)
);

AO22x2_ASAP7_75t_L g918 ( 
.A1(n_866),
.A2(n_690),
.B1(n_700),
.B2(n_687),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_867),
.A2(n_654),
.B1(n_684),
.B2(n_670),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_895),
.B(n_872),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_897),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_908),
.B(n_872),
.Y(n_922)
);

BUFx6f_ASAP7_75t_SL g923 ( 
.A(n_899),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_902),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_907),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_915),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_892),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_913),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_918),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_918),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_901),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_901),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_914),
.B(n_877),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_894),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_916),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_917),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_909),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_SL g938 ( 
.A(n_904),
.B(n_650),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_890),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_906),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_903),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_900),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_893),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_919),
.B(n_886),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_898),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_905),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_911),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_912),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_891),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_896),
.B(n_875),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_910),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_897),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_897),
.Y(n_953)
);

CKINVDCx16_ASAP7_75t_R g954 ( 
.A(n_909),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_899),
.B(n_688),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_908),
.B(n_784),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_895),
.B(n_877),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_897),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_897),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_894),
.A2(n_705),
.B(n_665),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_935),
.B(n_608),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_920),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_922),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_926),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_956),
.B(n_609),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_931),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_933),
.Y(n_968)
);

AND2x2_ASAP7_75t_SL g969 ( 
.A(n_955),
.B(n_859),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_934),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_960),
.B(n_617),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_921),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_936),
.B(n_619),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_942),
.B(n_941),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_932),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_928),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_944),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_940),
.B(n_683),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_924),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_927),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_939),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_947),
.B(n_632),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_949),
.B(n_760),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_948),
.B(n_637),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_925),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_952),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_929),
.A2(n_667),
.B(n_664),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_946),
.B(n_708),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_953),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_938),
.B(n_760),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_930),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_R g992 ( 
.A(n_945),
.B(n_951),
.Y(n_992)
);

AND2x6_ASAP7_75t_L g993 ( 
.A(n_958),
.B(n_641),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_950),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_937),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_923),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_923),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_955),
.B(n_829),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_943),
.B(n_646),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_954),
.B(n_648),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_954),
.A2(n_797),
.B(n_714),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_922),
.B(n_886),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_920),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_922),
.B(n_709),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_922),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_922),
.B(n_742),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_923),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_922),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_920),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_920),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_922),
.B(n_756),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_959),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_922),
.B(n_793),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_942),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_955),
.B(n_859),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_922),
.B(n_691),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_920),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_959),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_922),
.B(n_720),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_922),
.B(n_725),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_931),
.B(n_656),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_946),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_922),
.B(n_726),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_922),
.B(n_743),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_959),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_942),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_920),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_935),
.B(n_671),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_934),
.B(n_832),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_934),
.B(n_815),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_922),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_920),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_922),
.B(n_745),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_922),
.B(n_758),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_931),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_922),
.B(n_763),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_922),
.B(n_765),
.Y(n_1037)
);

BUFx2_ASAP7_75t_SL g1038 ( 
.A(n_934),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_920),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_935),
.B(n_692),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_920),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_959),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_920),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_922),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_935),
.B(n_710),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_920),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_922),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_997),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_997),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_1038),
.B(n_712),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_1007),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_967),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_997),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_971),
.B(n_717),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_983),
.B(n_772),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_966),
.B(n_734),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_1004),
.Y(n_1057)
);

CKINVDCx8_ASAP7_75t_R g1058 ( 
.A(n_1038),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_976),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_975),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_1035),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1002),
.B(n_713),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_1035),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_995),
.B(n_874),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_990),
.B(n_751),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_1000),
.B(n_785),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_994),
.B(n_847),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_964),
.B(n_719),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_984),
.B(n_754),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_974),
.B(n_794),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1014),
.B(n_799),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_981),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_982),
.B(n_757),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1026),
.B(n_801),
.Y(n_1074)
);

BUFx4f_ASAP7_75t_SL g1075 ( 
.A(n_1022),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_991),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_977),
.B(n_803),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_962),
.Y(n_1078)
);

INVx6_ASAP7_75t_L g1079 ( 
.A(n_999),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_1044),
.B(n_721),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_970),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1005),
.B(n_727),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_963),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_969),
.B(n_804),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1035),
.B(n_762),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_1006),
.B(n_817),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1015),
.B(n_822),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_970),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_1022),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1016),
.B(n_768),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1009),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1008),
.B(n_730),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1010),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1003),
.B(n_601),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1011),
.B(n_851),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1013),
.B(n_831),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1019),
.B(n_771),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_1003),
.B(n_701),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1027),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_996),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1017),
.B(n_747),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1032),
.Y(n_1102)
);

CKINVDCx16_ASAP7_75t_R g1103 ( 
.A(n_998),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_988),
.B(n_782),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_986),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1021),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1020),
.B(n_833),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1039),
.Y(n_1108)
);

BUFx2_ASAP7_75t_SL g1109 ( 
.A(n_1017),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1021),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1012),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_988),
.Y(n_1112)
);

AND2x6_ASAP7_75t_L g1113 ( 
.A(n_1041),
.B(n_773),
.Y(n_1113)
);

BUFx8_ASAP7_75t_SL g1114 ( 
.A(n_999),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1043),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_968),
.Y(n_1116)
);

BUFx8_ASAP7_75t_SL g1117 ( 
.A(n_978),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1046),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_985),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1001),
.B(n_836),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_1031),
.B(n_788),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1047),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1033),
.B(n_778),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1034),
.B(n_842),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1036),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1018),
.Y(n_1127)
);

AND2x6_ASAP7_75t_SL g1128 ( 
.A(n_973),
.B(n_858),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1037),
.B(n_855),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1029),
.B(n_856),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_980),
.B(n_796),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1030),
.B(n_857),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1025),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_979),
.B(n_800),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_989),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_961),
.B(n_783),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1042),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1028),
.B(n_795),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1040),
.B(n_602),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1045),
.B(n_818),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_965),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_987),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_972),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_992),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_993),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_993),
.B(n_835),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_967),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_976),
.Y(n_1148)
);

INVx6_ASAP7_75t_L g1149 ( 
.A(n_997),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1002),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1002),
.B(n_838),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_1038),
.B(n_844),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1002),
.B(n_845),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1000),
.B(n_603),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1038),
.B(n_622),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_967),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1002),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1002),
.B(n_812),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_995),
.B(n_606),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_997),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_976),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_967),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_983),
.B(n_607),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_967),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_967),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_969),
.B(n_610),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1000),
.B(n_802),
.Y(n_1167)
);

NAND2x1_ASAP7_75t_L g1168 ( 
.A(n_1035),
.B(n_702),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_967),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_971),
.B(n_807),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1004),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_971),
.B(n_811),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_983),
.B(n_612),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_1038),
.B(n_859),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1002),
.B(n_813),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_971),
.B(n_827),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_983),
.B(n_615),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_SL g1178 ( 
.A(n_969),
.B(n_616),
.Y(n_1178)
);

NAND2x1_ASAP7_75t_L g1179 ( 
.A(n_1035),
.B(n_702),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_967),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1103),
.B(n_834),
.Y(n_1181)
);

BUFx5_ASAP7_75t_L g1182 ( 
.A(n_1060),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1049),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_1053),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_1149),
.Y(n_1185)
);

BUFx2_ASAP7_75t_SL g1186 ( 
.A(n_1049),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1048),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1156),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1164),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1160),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1119),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1148),
.Y(n_1192)
);

BUFx2_ASAP7_75t_SL g1193 ( 
.A(n_1058),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1148),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1161),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1120),
.B(n_618),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1122),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1100),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1070),
.B(n_624),
.Y(n_1199)
);

BUFx4_ASAP7_75t_SL g1200 ( 
.A(n_1051),
.Y(n_1200)
);

INVx3_ASAP7_75t_SL g1201 ( 
.A(n_1116),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1161),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_1089),
.Y(n_1203)
);

INVx6_ASAP7_75t_SL g1204 ( 
.A(n_1104),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1123),
.B(n_841),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1079),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1061),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1106),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_1114),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1075),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1078),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1169),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1057),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1117),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1066),
.B(n_854),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1171),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1061),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1063),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1106),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1109),
.B(n_775),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1083),
.Y(n_1221)
);

BUFx8_ASAP7_75t_L g1222 ( 
.A(n_1112),
.Y(n_1222)
);

INVx5_ASAP7_75t_SL g1223 ( 
.A(n_1155),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1091),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1063),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1050),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1105),
.B(n_779),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1068),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1128),
.Y(n_1229)
);

BUFx4f_ASAP7_75t_SL g1230 ( 
.A(n_1101),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1110),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_SL g1232 ( 
.A(n_1080),
.Y(n_1232)
);

INVx6_ASAP7_75t_SL g1233 ( 
.A(n_1152),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1064),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1084),
.B(n_1087),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1093),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1076),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1067),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1121),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1052),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1110),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1059),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1062),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1151),
.Y(n_1244)
);

BUFx12f_ASAP7_75t_L g1245 ( 
.A(n_1153),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1134),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1147),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1162),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1158),
.Y(n_1249)
);

CKINVDCx11_ASAP7_75t_R g1250 ( 
.A(n_1174),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1099),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1081),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1082),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1092),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1102),
.Y(n_1255)
);

INVx6_ASAP7_75t_SL g1256 ( 
.A(n_1131),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1165),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1141),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1088),
.B(n_808),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1108),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1140),
.B(n_629),
.Y(n_1261)
);

BUFx2_ASAP7_75t_SL g1262 ( 
.A(n_1126),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1150),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1144),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1135),
.Y(n_1265)
);

NOR2x1_ASAP7_75t_SL g1266 ( 
.A(n_1085),
.B(n_1180),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1175),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_SL g1268 ( 
.A(n_1065),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1115),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1159),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1055),
.B(n_635),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1086),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1145),
.B(n_840),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1118),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1065),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1143),
.B(n_636),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1095),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1072),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1111),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1127),
.Y(n_1281)
);

CKINVDCx16_ASAP7_75t_R g1282 ( 
.A(n_1166),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1178),
.A2(n_850),
.B1(n_736),
.B2(n_645),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1113),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1191),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1235),
.A2(n_1065),
.B1(n_1132),
.B2(n_1130),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1196),
.A2(n_1173),
.B1(n_1177),
.B2(n_1163),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1270),
.A2(n_1090),
.B1(n_1124),
.B2(n_1097),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1184),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1185),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1283),
.A2(n_1096),
.B1(n_1113),
.B2(n_1107),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1211),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1201),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1198),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1221),
.Y(n_1295)
);

INVx6_ASAP7_75t_L g1296 ( 
.A(n_1192),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1238),
.B(n_1125),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1240),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1260),
.A2(n_1113),
.B1(n_1129),
.B2(n_1077),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1224),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1236),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1199),
.B(n_1154),
.Y(n_1302)
);

CKINVDCx6p67_ASAP7_75t_R g1303 ( 
.A(n_1209),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1282),
.A2(n_1167),
.B1(n_1054),
.B2(n_1170),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1275),
.A2(n_1071),
.B1(n_1074),
.B2(n_1146),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1251),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1255),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1247),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1273),
.A2(n_1176),
.B1(n_1172),
.B2(n_1069),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1269),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1248),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1213),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1200),
.Y(n_1313)
);

CKINVDCx6p67_ASAP7_75t_R g1314 ( 
.A(n_1209),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1278),
.A2(n_1073),
.B1(n_1056),
.B2(n_1098),
.Y(n_1315)
);

BUFx12f_ASAP7_75t_L g1316 ( 
.A(n_1250),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1242),
.A2(n_1137),
.B1(n_1133),
.B2(n_1094),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1195),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1194),
.B(n_1142),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1272),
.A2(n_1139),
.B1(n_1136),
.B2(n_1138),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1284),
.A2(n_736),
.B1(n_1179),
.B2(n_1168),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1234),
.A2(n_647),
.B1(n_653),
.B2(n_638),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1257),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1281),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1188),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1189),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1212),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1203),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1268),
.A2(n_672),
.B1(n_673),
.B2(n_663),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1229),
.A2(n_678),
.B1(n_679),
.B2(n_675),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1202),
.Y(n_1332)
);

CKINVDCx11_ASAP7_75t_R g1333 ( 
.A(n_1243),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1226),
.A2(n_681),
.B1(n_682),
.B2(n_680),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1181),
.A2(n_723),
.B1(n_746),
.B2(n_698),
.Y(n_1335)
);

INVx8_ASAP7_75t_L g1336 ( 
.A(n_1202),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1216),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1280),
.Y(n_1338)
);

BUFx2_ASAP7_75t_SL g1339 ( 
.A(n_1187),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1237),
.B(n_685),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1182),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1222),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1182),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1264),
.A2(n_693),
.B1(n_694),
.B2(n_686),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1215),
.A2(n_4),
.B(n_5),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1279),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1226),
.A2(n_696),
.B1(n_699),
.B2(n_695),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1214),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1230),
.Y(n_1349)
);

CKINVDCx14_ASAP7_75t_R g1350 ( 
.A(n_1214),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1279),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1254),
.B(n_707),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1190),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1249),
.A2(n_1267),
.B(n_1239),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1271),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1266),
.Y(n_1356)
);

INVx6_ASAP7_75t_L g1357 ( 
.A(n_1245),
.Y(n_1357)
);

INVx5_ASAP7_75t_L g1358 ( 
.A(n_1241),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1246),
.A2(n_718),
.B1(n_728),
.B2(n_716),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1241),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1197),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1183),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1205),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1265),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1253),
.A2(n_732),
.B1(n_737),
.B2(n_731),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1204),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1258),
.Y(n_1367)
);

INVx11_ASAP7_75t_L g1368 ( 
.A(n_1186),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1246),
.A2(n_769),
.B1(n_790),
.B2(n_755),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1262),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1261),
.A2(n_740),
.B1(n_741),
.B2(n_739),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1276),
.A2(n_750),
.B1(n_752),
.B2(n_748),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1193),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1277),
.A2(n_759),
.B1(n_761),
.B2(n_753),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_L g1375 ( 
.A(n_1208),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1210),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1219),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1232),
.A2(n_824),
.B1(n_825),
.B2(n_823),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1231),
.B(n_766),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1217),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1218),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1220),
.A2(n_770),
.B1(n_774),
.B2(n_767),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1228),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1244),
.A2(n_777),
.B1(n_780),
.B2(n_776),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1244),
.A2(n_810),
.B1(n_814),
.B2(n_809),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1263),
.B(n_786),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1227),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1207),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1274),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1225),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1206),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1252),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1233),
.A2(n_791),
.B1(n_792),
.B2(n_787),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1259),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1223),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1297),
.B(n_805),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1288),
.A2(n_1304),
.B1(n_1286),
.B2(n_1363),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1287),
.A2(n_1256),
.B1(n_843),
.B2(n_816),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1298),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1302),
.B(n_1379),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1305),
.B(n_806),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1299),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1308),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1293),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1309),
.A2(n_819),
.B1(n_830),
.B2(n_828),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1291),
.A2(n_849),
.B1(n_853),
.B2(n_852),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1313),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1321),
.A2(n_839),
.B1(n_8),
.B2(n_6),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1342),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1315),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1285),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1337),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1345),
.A2(n_13),
.B(n_12),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1331),
.A2(n_22),
.B1(n_30),
.B2(n_9),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1312),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1340),
.B(n_14),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1344),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1292),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1323),
.A2(n_18),
.B(n_17),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1356),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_1420)
);

BUFx4f_ASAP7_75t_SL g1421 ( 
.A(n_1303),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1295),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1300),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1336),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1335),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1330),
.A2(n_1393),
.B(n_1359),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1350),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1318),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1311),
.B(n_27),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1371),
.A2(n_1374),
.B1(n_1329),
.B2(n_1394),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1301),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1306),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1370),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1355),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1307),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1310),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1325),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1368),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1384),
.A2(n_1334),
.B1(n_1347),
.B2(n_1395),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1320),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1346),
.B(n_32),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1382),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1389),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1443)
);

CKINVDCx14_ASAP7_75t_R g1444 ( 
.A(n_1289),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1387),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1324),
.B(n_38),
.Y(n_1446)
);

INVx5_ASAP7_75t_L g1447 ( 
.A(n_1336),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1354),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1326),
.Y(n_1449)
);

NOR2x1_ASAP7_75t_R g1450 ( 
.A(n_1333),
.B(n_324),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1353),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1316),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1327),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1328),
.B(n_1352),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1341),
.A2(n_329),
.B(n_328),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1365),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1378),
.A2(n_1386),
.B(n_1369),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1357),
.A2(n_53),
.B1(n_62),
.B2(n_45),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1317),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1372),
.A2(n_1338),
.B1(n_1361),
.B2(n_1364),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1358),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_SL g1462 ( 
.A1(n_1385),
.A2(n_48),
.B(n_47),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1376),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1317),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1408),
.A2(n_1348),
.B1(n_1314),
.B2(n_1351),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1397),
.A2(n_1373),
.B1(n_1290),
.B2(n_1339),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1400),
.B(n_1380),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1417),
.A2(n_1343),
.B1(n_1290),
.B2(n_1322),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1462),
.B(n_1391),
.C(n_1381),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1456),
.A2(n_1367),
.B1(n_1294),
.B2(n_1366),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1427),
.A2(n_1349),
.B1(n_1358),
.B2(n_1362),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1457),
.A2(n_1383),
.B1(n_1388),
.B2(n_1392),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1440),
.B(n_1360),
.Y(n_1473)
);

OAI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1413),
.A2(n_1426),
.B1(n_1398),
.B2(n_1419),
.C(n_1414),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1399),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1411),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1448),
.A2(n_1391),
.B1(n_1377),
.B2(n_1360),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1415),
.B(n_1332),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1412),
.B(n_1454),
.Y(n_1479)
);

OAI222xp33_ASAP7_75t_L g1480 ( 
.A1(n_1410),
.A2(n_1390),
.B1(n_49),
.B2(n_51),
.C1(n_46),
.C2(n_48),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1425),
.A2(n_1375),
.B1(n_1319),
.B2(n_1296),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1428),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1405),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1459),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1442),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1433),
.A2(n_1401),
.B1(n_1416),
.B2(n_1444),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1403),
.B(n_56),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_SL g1488 ( 
.A(n_1443),
.B(n_57),
.C(n_58),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1402),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1420),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.Y(n_1490)
);

AOI222xp33_ASAP7_75t_L g1491 ( 
.A1(n_1434),
.A2(n_66),
.B1(n_68),
.B2(n_64),
.C1(n_65),
.C2(n_67),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1446),
.B(n_331),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1445),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1440),
.B(n_70),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1453),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1458),
.B(n_73),
.C(n_74),
.Y(n_1496)
);

OAI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1439),
.A2(n_77),
.B1(n_74),
.B2(n_75),
.C(n_78),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1449),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1430),
.A2(n_1396),
.B1(n_1460),
.B2(n_1406),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1441),
.B(n_333),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1429),
.B(n_334),
.Y(n_1501)
);

OAI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1418),
.A2(n_82),
.B1(n_84),
.B2(n_80),
.C1(n_81),
.C2(n_83),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1451),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1422),
.B(n_85),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1474),
.A2(n_1461),
.B(n_1450),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1499),
.A2(n_1447),
.B1(n_1431),
.B2(n_1432),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1467),
.B(n_1423),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1498),
.B(n_1435),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1475),
.B(n_1436),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1476),
.B(n_1437),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1469),
.A2(n_1497),
.B(n_1483),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1491),
.B(n_1455),
.C(n_1447),
.Y(n_1512)
);

OAI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1496),
.A2(n_1463),
.B1(n_1404),
.B2(n_1421),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1501),
.B(n_1464),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1486),
.A2(n_1424),
.B1(n_1438),
.B2(n_1447),
.C(n_1407),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1479),
.B(n_1464),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1466),
.B(n_1438),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_SL g1518 ( 
.A(n_1480),
.B(n_1409),
.Y(n_1518)
);

NAND4xp25_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_88),
.C(n_86),
.D(n_87),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1503),
.B(n_1452),
.C(n_90),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_89),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1478),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_L g1523 ( 
.A(n_1488),
.B(n_91),
.C(n_92),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1504),
.B(n_92),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1489),
.A2(n_1482),
.B(n_1477),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_93),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1487),
.B(n_94),
.Y(n_1527)
);

OAI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1471),
.A2(n_98),
.B1(n_95),
.B2(n_97),
.C(n_99),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1473),
.B(n_97),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1472),
.B(n_98),
.Y(n_1530)
);

AOI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1502),
.A2(n_103),
.B1(n_100),
.B2(n_101),
.C(n_104),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1485),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1495),
.A2(n_338),
.B(n_335),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1494),
.B(n_105),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1473),
.B(n_107),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1484),
.B(n_107),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1493),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1470),
.B(n_108),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1465),
.B(n_111),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1468),
.B(n_339),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_SL g1541 ( 
.A1(n_1490),
.A2(n_113),
.B(n_112),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1481),
.B(n_111),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1474),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1474),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1519),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1508),
.B(n_119),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1507),
.B(n_120),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_121),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_121),
.Y(n_1549)
);

OAI211xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1530),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_L g1551 ( 
.A(n_1543),
.B(n_124),
.C(n_125),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_127),
.C(n_128),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1514),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1534),
.Y(n_1554)
);

NOR3xp33_ASAP7_75t_L g1555 ( 
.A(n_1520),
.B(n_129),
.C(n_130),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1506),
.B(n_1524),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1520),
.A2(n_1532),
.B1(n_1531),
.B2(n_1525),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.B(n_1526),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_131),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1535),
.B(n_131),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_132),
.C(n_133),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1536),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1544),
.B(n_134),
.C(n_135),
.Y(n_1563)
);

AOI211x1_ASAP7_75t_L g1564 ( 
.A1(n_1513),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1521),
.B(n_140),
.Y(n_1565)
);

AND4x1_ASAP7_75t_L g1566 ( 
.A(n_1512),
.B(n_143),
.C(n_141),
.D(n_142),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1517),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1538),
.B(n_141),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1539),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1505),
.B(n_142),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1571)
);

AOI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1541),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.C(n_150),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1540),
.B(n_1533),
.Y(n_1573)
);

NOR3xp33_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_149),
.C(n_150),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1510),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1522),
.B(n_151),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1523),
.B(n_151),
.C(n_152),
.Y(n_1577)
);

NOR3xp33_ASAP7_75t_L g1578 ( 
.A(n_1520),
.B(n_152),
.C(n_153),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1519),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1579)
);

NOR3xp33_ASAP7_75t_L g1580 ( 
.A(n_1520),
.B(n_154),
.C(n_156),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1520),
.B(n_157),
.C(n_158),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1510),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1523),
.B(n_157),
.C(n_158),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1523),
.B(n_159),
.C(n_160),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1522),
.B(n_162),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1516),
.B(n_162),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1510),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1522),
.B(n_163),
.Y(n_1588)
);

OAI211xp5_ASAP7_75t_L g1589 ( 
.A1(n_1519),
.A2(n_172),
.B(n_181),
.C(n_163),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1510),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1522),
.B(n_164),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1510),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1510),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1518),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1519),
.A2(n_168),
.B(n_169),
.Y(n_1595)
);

AOI31xp33_ASAP7_75t_L g1596 ( 
.A1(n_1520),
.A2(n_173),
.A3(n_170),
.B(n_172),
.Y(n_1596)
);

OAI211xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1530),
.A2(n_174),
.B(n_170),
.C(n_173),
.Y(n_1597)
);

NAND4xp75_ASAP7_75t_SL g1598 ( 
.A(n_1576),
.B(n_177),
.C(n_174),
.D(n_176),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1575),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1567),
.B(n_176),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1590),
.B(n_178),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1593),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1582),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1593),
.B(n_1553),
.Y(n_1604)
);

XOR2x2_ASAP7_75t_L g1605 ( 
.A(n_1558),
.B(n_180),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1587),
.Y(n_1606)
);

XOR2x2_ASAP7_75t_L g1607 ( 
.A(n_1594),
.B(n_1557),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1554),
.B(n_182),
.Y(n_1608)
);

NAND4xp75_ASAP7_75t_L g1609 ( 
.A(n_1595),
.B(n_185),
.C(n_182),
.D(n_184),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1569),
.B(n_187),
.Y(n_1610)
);

NOR4xp25_ASAP7_75t_L g1611 ( 
.A(n_1550),
.B(n_190),
.C(n_188),
.D(n_189),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1592),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_188),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1546),
.B(n_189),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1556),
.B(n_191),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1585),
.B(n_192),
.Y(n_1616)
);

NAND4xp75_ASAP7_75t_L g1617 ( 
.A(n_1572),
.B(n_194),
.C(n_192),
.D(n_193),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1588),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1548),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1591),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1549),
.B(n_1586),
.Y(n_1621)
);

NAND4xp75_ASAP7_75t_L g1622 ( 
.A(n_1570),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_1622)
);

XOR2x2_ASAP7_75t_L g1623 ( 
.A(n_1566),
.B(n_196),
.Y(n_1623)
);

NAND4xp75_ASAP7_75t_SL g1624 ( 
.A(n_1596),
.B(n_200),
.C(n_197),
.D(n_198),
.Y(n_1624)
);

XOR2x2_ASAP7_75t_L g1625 ( 
.A(n_1555),
.B(n_198),
.Y(n_1625)
);

NAND4xp75_ASAP7_75t_SL g1626 ( 
.A(n_1561),
.B(n_1580),
.C(n_1581),
.D(n_1578),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1571),
.Y(n_1627)
);

XNOR2xp5_ASAP7_75t_L g1628 ( 
.A(n_1565),
.B(n_200),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1547),
.B(n_201),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1560),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1559),
.B(n_202),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1568),
.B(n_202),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1573),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1597),
.B(n_204),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1577),
.B(n_205),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1583),
.Y(n_1636)
);

NAND4xp75_ASAP7_75t_SL g1637 ( 
.A(n_1589),
.B(n_1551),
.C(n_1584),
.D(n_1579),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1563),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1574),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1545),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1575),
.Y(n_1641)
);

XOR2xp5_ASAP7_75t_L g1642 ( 
.A(n_1571),
.B(n_341),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1575),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1575),
.Y(n_1644)
);

NAND4xp75_ASAP7_75t_SL g1645 ( 
.A(n_1576),
.B(n_209),
.C(n_207),
.D(n_208),
.Y(n_1645)
);

XNOR2x2_ASAP7_75t_L g1646 ( 
.A(n_1552),
.B(n_210),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1575),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1554),
.Y(n_1648)
);

OAI21xp33_ASAP7_75t_L g1649 ( 
.A1(n_1557),
.A2(n_211),
.B(n_212),
.Y(n_1649)
);

XOR2x2_ASAP7_75t_L g1650 ( 
.A(n_1558),
.B(n_211),
.Y(n_1650)
);

XNOR2xp5_ASAP7_75t_L g1651 ( 
.A(n_1558),
.B(n_212),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1575),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1554),
.B(n_214),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1575),
.B(n_215),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1575),
.B(n_215),
.Y(n_1655)
);

XOR2x2_ASAP7_75t_L g1656 ( 
.A(n_1558),
.B(n_217),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1575),
.B(n_218),
.Y(n_1657)
);

NAND4xp75_ASAP7_75t_SL g1658 ( 
.A(n_1576),
.B(n_221),
.C(n_218),
.D(n_219),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1575),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1575),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1575),
.Y(n_1661)
);

NAND4xp75_ASAP7_75t_L g1662 ( 
.A(n_1564),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1627),
.B(n_222),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1614),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1641),
.Y(n_1665)
);

XNOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1650),
.B(n_226),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1604),
.Y(n_1667)
);

XOR2x2_ASAP7_75t_L g1668 ( 
.A(n_1656),
.B(n_1607),
.Y(n_1668)
);

XOR2x2_ASAP7_75t_L g1669 ( 
.A(n_1651),
.B(n_225),
.Y(n_1669)
);

AO22x2_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_227),
.B1(n_228),
.B2(n_226),
.Y(n_1670)
);

XOR2x2_ASAP7_75t_L g1671 ( 
.A(n_1623),
.B(n_1628),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1599),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1643),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1633),
.B(n_227),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1644),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1619),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1647),
.Y(n_1677)
);

XNOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1625),
.B(n_230),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1652),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1602),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1659),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1630),
.B(n_229),
.Y(n_1682)
);

XOR2xp5_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_231),
.Y(n_1683)
);

OA22x2_ASAP7_75t_L g1684 ( 
.A1(n_1636),
.A2(n_234),
.B1(n_231),
.B2(n_232),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1660),
.B(n_232),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1621),
.Y(n_1686)
);

XOR2x2_ASAP7_75t_L g1687 ( 
.A(n_1637),
.B(n_234),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1661),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1618),
.B(n_237),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1648),
.B(n_240),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1620),
.Y(n_1691)
);

AND2x6_ASAP7_75t_L g1692 ( 
.A(n_1639),
.B(n_242),
.Y(n_1692)
);

XOR2x2_ASAP7_75t_L g1693 ( 
.A(n_1646),
.B(n_241),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1603),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1612),
.Y(n_1695)
);

XOR2x2_ASAP7_75t_L g1696 ( 
.A(n_1624),
.B(n_241),
.Y(n_1696)
);

INVxp67_ASAP7_75t_SL g1697 ( 
.A(n_1608),
.Y(n_1697)
);

XNOR2x2_ASAP7_75t_L g1698 ( 
.A(n_1622),
.B(n_243),
.Y(n_1698)
);

XNOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1631),
.B(n_245),
.Y(n_1699)
);

AOI22x1_ASAP7_75t_SL g1700 ( 
.A1(n_1638),
.A2(n_247),
.B1(n_244),
.B2(n_246),
.Y(n_1700)
);

XNOR2xp5_ASAP7_75t_L g1701 ( 
.A(n_1598),
.B(n_1645),
.Y(n_1701)
);

XOR2x2_ASAP7_75t_L g1702 ( 
.A(n_1617),
.B(n_244),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1601),
.Y(n_1703)
);

XOR2x2_ASAP7_75t_L g1704 ( 
.A(n_1609),
.B(n_249),
.Y(n_1704)
);

XOR2x2_ASAP7_75t_L g1705 ( 
.A(n_1658),
.B(n_251),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1654),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1655),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1613),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1657),
.B(n_251),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1632),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1653),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1615),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1635),
.Y(n_1713)
);

CKINVDCx8_ASAP7_75t_R g1714 ( 
.A(n_1610),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1629),
.B(n_252),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1640),
.B(n_253),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1616),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1600),
.B(n_254),
.Y(n_1718)
);

CKINVDCx16_ASAP7_75t_R g1719 ( 
.A(n_1634),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1611),
.B(n_255),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1649),
.Y(n_1721)
);

XOR2xp5_ASAP7_75t_L g1722 ( 
.A(n_1662),
.B(n_255),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1641),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1641),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1641),
.Y(n_1725)
);

XNOR2x1_ASAP7_75t_L g1726 ( 
.A(n_1605),
.B(n_259),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1606),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1602),
.Y(n_1728)
);

XNOR2x2_ASAP7_75t_L g1729 ( 
.A(n_1646),
.B(n_258),
.Y(n_1729)
);

XOR2x2_ASAP7_75t_L g1730 ( 
.A(n_1605),
.B(n_259),
.Y(n_1730)
);

INVxp33_ASAP7_75t_L g1731 ( 
.A(n_1642),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1641),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1641),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1691),
.Y(n_1734)
);

XNOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1668),
.B(n_260),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1694),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1727),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1695),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1720),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1676),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1672),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1682),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1729),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1670),
.A2(n_269),
.B1(n_266),
.B2(n_268),
.Y(n_1744)
);

XNOR2x1_ASAP7_75t_L g1745 ( 
.A(n_1678),
.B(n_270),
.Y(n_1745)
);

AO22x2_ASAP7_75t_L g1746 ( 
.A1(n_1703),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1663),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1665),
.Y(n_1748)
);

OA22x2_ASAP7_75t_L g1749 ( 
.A1(n_1721),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1673),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1675),
.Y(n_1751)
);

OA22x2_ASAP7_75t_L g1752 ( 
.A1(n_1701),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_1752)
);

OA22x2_ASAP7_75t_L g1753 ( 
.A1(n_1686),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_1753)
);

OA22x2_ASAP7_75t_L g1754 ( 
.A1(n_1664),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1677),
.Y(n_1755)
);

OAI22x1_ASAP7_75t_L g1756 ( 
.A1(n_1697),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1710),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1679),
.Y(n_1758)
);

OA22x2_ASAP7_75t_L g1759 ( 
.A1(n_1683),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1687),
.A2(n_291),
.B1(n_288),
.B2(n_290),
.Y(n_1760)
);

AO22x1_ASAP7_75t_L g1761 ( 
.A1(n_1692),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.Y(n_1761)
);

AOI22x1_ASAP7_75t_L g1762 ( 
.A1(n_1712),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1680),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1728),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1692),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1681),
.Y(n_1766)
);

OA22x2_ASAP7_75t_L g1767 ( 
.A1(n_1711),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_1767)
);

XNOR2xp5_ASAP7_75t_L g1768 ( 
.A(n_1730),
.B(n_299),
.Y(n_1768)
);

CKINVDCx16_ASAP7_75t_R g1769 ( 
.A(n_1700),
.Y(n_1769)
);

OA22x2_ASAP7_75t_L g1770 ( 
.A1(n_1708),
.A2(n_1717),
.B1(n_1667),
.B2(n_1723),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1714),
.A2(n_1726),
.B1(n_1666),
.B2(n_1684),
.Y(n_1771)
);

OA22x2_ASAP7_75t_L g1772 ( 
.A1(n_1724),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_1772)
);

OA22x2_ASAP7_75t_L g1773 ( 
.A1(n_1725),
.A2(n_303),
.B1(n_300),
.B2(n_301),
.Y(n_1773)
);

XNOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1669),
.B(n_303),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1688),
.Y(n_1775)
);

OA22x2_ASAP7_75t_L g1776 ( 
.A1(n_1732),
.A2(n_1733),
.B1(n_1706),
.B2(n_1707),
.Y(n_1776)
);

XOR2x2_ASAP7_75t_L g1777 ( 
.A(n_1699),
.B(n_1702),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1685),
.Y(n_1778)
);

XOR2x2_ASAP7_75t_L g1779 ( 
.A(n_1704),
.B(n_305),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1689),
.Y(n_1780)
);

BUFx12f_ASAP7_75t_L g1781 ( 
.A(n_1715),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1674),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1716),
.Y(n_1783)
);

XOR2x2_ASAP7_75t_L g1784 ( 
.A(n_1698),
.B(n_307),
.Y(n_1784)
);

AO22x2_ASAP7_75t_L g1785 ( 
.A1(n_1690),
.A2(n_312),
.B1(n_308),
.B2(n_310),
.Y(n_1785)
);

OA22x2_ASAP7_75t_L g1786 ( 
.A1(n_1709),
.A2(n_313),
.B1(n_310),
.B2(n_312),
.Y(n_1786)
);

XOR2x2_ASAP7_75t_L g1787 ( 
.A(n_1696),
.B(n_313),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1705),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1718),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1731),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1691),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1691),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1719),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_1793)
);

XOR2x2_ASAP7_75t_L g1794 ( 
.A(n_1668),
.B(n_314),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1691),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1676),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1719),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1691),
.Y(n_1798)
);

XNOR2x1_ASAP7_75t_L g1799 ( 
.A(n_1668),
.B(n_317),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1713),
.B(n_318),
.Y(n_1800)
);

XOR2x2_ASAP7_75t_L g1801 ( 
.A(n_1668),
.B(n_319),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1719),
.B(n_321),
.Y(n_1802)
);

INVx8_ASAP7_75t_L g1803 ( 
.A(n_1692),
.Y(n_1803)
);

INVx4_ASAP7_75t_L g1804 ( 
.A(n_1692),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1719),
.A2(n_322),
.B1(n_343),
.B2(n_342),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1727),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1719),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_1807)
);

OA22x2_ASAP7_75t_L g1808 ( 
.A1(n_1722),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_1808)
);

OA22x2_ASAP7_75t_L g1809 ( 
.A1(n_1722),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_1809)
);

OA22x2_ASAP7_75t_L g1810 ( 
.A1(n_1722),
.A2(n_360),
.B1(n_357),
.B2(n_358),
.Y(n_1810)
);

OA22x2_ASAP7_75t_L g1811 ( 
.A1(n_1722),
.A2(n_366),
.B1(n_362),
.B2(n_363),
.Y(n_1811)
);

INVx3_ASAP7_75t_SL g1812 ( 
.A(n_1693),
.Y(n_1812)
);

OA22x2_ASAP7_75t_L g1813 ( 
.A1(n_1722),
.A2(n_370),
.B1(n_367),
.B2(n_369),
.Y(n_1813)
);

OA22x2_ASAP7_75t_L g1814 ( 
.A1(n_1722),
.A2(n_374),
.B1(n_372),
.B2(n_373),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1719),
.A2(n_378),
.B1(n_375),
.B2(n_377),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1719),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_1816)
);

OAI22x1_ASAP7_75t_L g1817 ( 
.A1(n_1713),
.A2(n_386),
.B1(n_382),
.B2(n_385),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1719),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1691),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1682),
.Y(n_1820)
);

XNOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1668),
.B(n_391),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1691),
.Y(n_1822)
);

OA22x2_ASAP7_75t_L g1823 ( 
.A1(n_1722),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1727),
.Y(n_1824)
);

XNOR2xp5_ASAP7_75t_L g1825 ( 
.A(n_1671),
.B(n_396),
.Y(n_1825)
);

XNOR2xp5_ASAP7_75t_L g1826 ( 
.A(n_1671),
.B(n_397),
.Y(n_1826)
);

AO22x1_ASAP7_75t_L g1827 ( 
.A1(n_1663),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_1827)
);

OA22x2_ASAP7_75t_L g1828 ( 
.A1(n_1722),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1727),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1727),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1727),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1719),
.A2(n_410),
.B1(n_407),
.B2(n_409),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1727),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1736),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1738),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1741),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1750),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1803),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1751),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1755),
.Y(n_1840)
);

BUFx4_ASAP7_75t_SL g1841 ( 
.A(n_1735),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1758),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1766),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1757),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1769),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_1845)
);

INVx8_ASAP7_75t_L g1846 ( 
.A(n_1803),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1775),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1783),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1812),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1740),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1804),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1747),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1780),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1796),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1782),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1742),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1764),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1734),
.Y(n_1858)
);

OAI322xp33_ASAP7_75t_L g1859 ( 
.A1(n_1739),
.A2(n_425),
.A3(n_424),
.B1(n_420),
.B2(n_416),
.C1(n_418),
.C2(n_422),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1791),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1820),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1792),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1795),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1798),
.Y(n_1864)
);

INVx5_ASAP7_75t_L g1865 ( 
.A(n_1784),
.Y(n_1865)
);

XOR2x2_ASAP7_75t_L g1866 ( 
.A(n_1794),
.B(n_427),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1776),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1778),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1781),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1819),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1748),
.Y(n_1871)
);

XOR2x2_ASAP7_75t_L g1872 ( 
.A(n_1801),
.B(n_1777),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1822),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1737),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1763),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1806),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1800),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1790),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1824),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1785),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1770),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1746),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1789),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1753),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1829),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1754),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1830),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1831),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1833),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1744),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1772),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1773),
.Y(n_1892)
);

INVxp33_ASAP7_75t_SL g1893 ( 
.A(n_1771),
.Y(n_1893)
);

OAI322xp33_ASAP7_75t_L g1894 ( 
.A1(n_1749),
.A2(n_434),
.A3(n_435),
.B1(n_436),
.B2(n_437),
.C1(n_438),
.C2(n_439),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1743),
.A2(n_443),
.B1(n_440),
.B2(n_441),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1767),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1799),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1802),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1756),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1788),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1752),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1786),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1745),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1761),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1762),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1765),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1850),
.Y(n_1907)
);

OAI322xp33_ASAP7_75t_L g1908 ( 
.A1(n_1880),
.A2(n_1760),
.A3(n_1793),
.B1(n_1797),
.B2(n_1759),
.C1(n_1774),
.C2(n_1768),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1838),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1854),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1873),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1871),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1834),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1835),
.Y(n_1914)
);

AO22x2_ASAP7_75t_L g1915 ( 
.A1(n_1852),
.A2(n_1821),
.B1(n_1779),
.B2(n_1787),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1869),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1851),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1836),
.Y(n_1918)
);

NAND4xp75_ASAP7_75t_L g1919 ( 
.A(n_1904),
.B(n_1815),
.C(n_1832),
.D(n_1816),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1837),
.Y(n_1920)
);

OAI322xp33_ASAP7_75t_L g1921 ( 
.A1(n_1882),
.A2(n_1828),
.A3(n_1808),
.B1(n_1809),
.B2(n_1810),
.C1(n_1823),
.C2(n_1811),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1839),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1840),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1842),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1843),
.Y(n_1925)
);

OAI322xp33_ASAP7_75t_L g1926 ( 
.A1(n_1884),
.A2(n_1814),
.A3(n_1813),
.B1(n_1825),
.B2(n_1826),
.C1(n_1805),
.C2(n_1807),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1893),
.A2(n_1818),
.B1(n_1827),
.B2(n_1817),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_1846),
.Y(n_1928)
);

BUFx4f_ASAP7_75t_SL g1929 ( 
.A(n_1878),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1847),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1883),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1849),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1844),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1865),
.A2(n_454),
.B1(n_451),
.B2(n_453),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1881),
.A2(n_458),
.B1(n_455),
.B2(n_456),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1901),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1875),
.Y(n_1937)
);

NOR2x1_ASAP7_75t_L g1938 ( 
.A(n_1900),
.B(n_1886),
.Y(n_1938)
);

OA22x2_ASAP7_75t_L g1939 ( 
.A1(n_1867),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_1939)
);

AOI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1865),
.A2(n_469),
.B1(n_466),
.B2(n_467),
.C(n_471),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1890),
.A2(n_476),
.B1(n_473),
.B2(n_474),
.Y(n_1941)
);

OAI322xp33_ASAP7_75t_L g1942 ( 
.A1(n_1891),
.A2(n_479),
.A3(n_482),
.B1(n_484),
.B2(n_485),
.C1(n_487),
.C2(n_488),
.Y(n_1942)
);

AO22x2_ASAP7_75t_L g1943 ( 
.A1(n_1861),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1853),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1872),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_1945)
);

OA22x2_ASAP7_75t_SL g1946 ( 
.A1(n_1899),
.A2(n_498),
.B1(n_495),
.B2(n_497),
.Y(n_1946)
);

OAI322xp33_ASAP7_75t_L g1947 ( 
.A1(n_1892),
.A2(n_499),
.A3(n_500),
.B1(n_501),
.B2(n_502),
.C1(n_504),
.C2(n_506),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1907),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1910),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1927),
.A2(n_1896),
.B1(n_1902),
.B2(n_1906),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1911),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1929),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1915),
.A2(n_1919),
.B1(n_1932),
.B2(n_1938),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_SL g1954 ( 
.A1(n_1916),
.A2(n_1845),
.B(n_1898),
.C(n_1905),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1912),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1935),
.A2(n_1856),
.B1(n_1897),
.B2(n_1868),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1913),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1939),
.A2(n_1877),
.B1(n_1857),
.B2(n_1876),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1909),
.A2(n_1888),
.B1(n_1889),
.B2(n_1887),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1914),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1918),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1920),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1945),
.A2(n_1879),
.B1(n_1885),
.B2(n_1874),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1922),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1923),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1924),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1925),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1933),
.A2(n_1903),
.B1(n_1848),
.B2(n_1860),
.Y(n_1968)
);

AO22x1_ASAP7_75t_SL g1969 ( 
.A1(n_1928),
.A2(n_1841),
.B1(n_1855),
.B2(n_1858),
.Y(n_1969)
);

O2A1O1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1908),
.A2(n_1863),
.B(n_1864),
.C(n_1862),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1955),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1948),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1949),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1951),
.Y(n_1974)
);

NAND2x1_ASAP7_75t_L g1975 ( 
.A(n_1952),
.B(n_1917),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1953),
.A2(n_1940),
.B1(n_1934),
.B2(n_1870),
.Y(n_1976)
);

AO22x1_ASAP7_75t_L g1977 ( 
.A1(n_1950),
.A2(n_1946),
.B1(n_1931),
.B2(n_1944),
.Y(n_1977)
);

NOR4xp25_ASAP7_75t_L g1978 ( 
.A(n_1970),
.B(n_1926),
.C(n_1930),
.D(n_1937),
.Y(n_1978)
);

AOI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1956),
.A2(n_1958),
.B1(n_1968),
.B2(n_1963),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1959),
.A2(n_1866),
.B1(n_1941),
.B2(n_1936),
.Y(n_1980)
);

NOR2x1_ASAP7_75t_L g1981 ( 
.A(n_1975),
.B(n_1957),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1971),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1972),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1978),
.B(n_1969),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1973),
.Y(n_1985)
);

AND4x1_ASAP7_75t_L g1986 ( 
.A(n_1981),
.B(n_1979),
.C(n_1976),
.D(n_1980),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1982),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1984),
.A2(n_1954),
.B(n_1977),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1983),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1985),
.Y(n_1990)
);

O2A1O1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1988),
.A2(n_1974),
.B(n_1960),
.C(n_1962),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1989),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1987),
.Y(n_1993)
);

AO22x2_ASAP7_75t_L g1994 ( 
.A1(n_1992),
.A2(n_1990),
.B1(n_1964),
.B2(n_1965),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1994),
.Y(n_1995)
);

AO22x2_ASAP7_75t_L g1996 ( 
.A1(n_1995),
.A2(n_1993),
.B1(n_1961),
.B2(n_1967),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1996),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1997),
.A2(n_1966),
.B1(n_1986),
.B2(n_1943),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1998),
.Y(n_1999)
);

AOI221xp5_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1991),
.B1(n_1921),
.B2(n_1942),
.C(n_1947),
.Y(n_2000)
);

AOI211xp5_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1894),
.B(n_1859),
.C(n_1895),
.Y(n_2001)
);


endmodule