module fake_jpeg_26330_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_32),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_22),
.B1(n_25),
.B2(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_22),
.B1(n_21),
.B2(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_59),
.Y(n_94)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_89),
.B1(n_38),
.B2(n_35),
.Y(n_104)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_22),
.B1(n_16),
.B2(n_17),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_86),
.B1(n_21),
.B2(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_17),
.B1(n_40),
.B2(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_85),
.B1(n_40),
.B2(n_35),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_41),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_17),
.B1(n_40),
.B2(n_38),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_21),
.B1(n_19),
.B2(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_36),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_19),
.B1(n_21),
.B2(n_35),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_101),
.B1(n_79),
.B2(n_85),
.Y(n_129)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_34),
.C(n_36),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_83),
.C(n_34),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_114),
.B1(n_82),
.B2(n_67),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_69),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_39),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_84),
.Y(n_140)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_88),
.B(n_61),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_120),
.A2(n_133),
.B(n_137),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_126),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_92),
.B1(n_90),
.B2(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_61),
.B1(n_80),
.B2(n_65),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_134),
.B1(n_139),
.B2(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_29),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_131),
.B(n_132),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_18),
.B1(n_27),
.B2(n_75),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_87),
.B1(n_70),
.B2(n_71),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_27),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_145),
.C(n_13),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_62),
.B1(n_81),
.B2(n_77),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_144),
.B1(n_23),
.B2(n_28),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_30),
.B1(n_28),
.B2(n_31),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_105),
.B1(n_114),
.B2(n_102),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_62),
.B1(n_67),
.B2(n_34),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_18),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_103),
.A2(n_78),
.B1(n_68),
.B2(n_59),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_113),
.B1(n_95),
.B2(n_36),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_147),
.B(n_154),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_149),
.B1(n_163),
.B2(n_165),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_109),
.B1(n_117),
.B2(n_106),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_32),
.B(n_113),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_9),
.B(n_14),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_28),
.B(n_30),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_169),
.B(n_170),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_121),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_39),
.C(n_33),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_168),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_121),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_172),
.B1(n_0),
.B2(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_11),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_95),
.B1(n_36),
.B2(n_39),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_116),
.C(n_24),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_127),
.C(n_1),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_178),
.B1(n_135),
.B2(n_1),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_167)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_30),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_116),
.B(n_1),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_142),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_122),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_128),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_186),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_185),
.B(n_203),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_118),
.B(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_9),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_6),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_213),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_157),
.B1(n_175),
.B2(n_165),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_180),
.B1(n_172),
.B2(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_223),
.B1(n_157),
.B2(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_234),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_182),
.C(n_164),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_229),
.C(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_179),
.C(n_198),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_186),
.B(n_196),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_237),
.B1(n_209),
.B2(n_174),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_179),
.C(n_150),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_205),
.C(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_203),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_151),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_168),
.C(n_190),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_190),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_180),
.B1(n_212),
.B2(n_181),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_237),
.A2(n_223),
.B1(n_211),
.B2(n_218),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_206),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_252),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_220),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_255),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_195),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_253),
.A2(n_241),
.B1(n_228),
.B2(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_156),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_256),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_173),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_212),
.B1(n_178),
.B2(n_219),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_250),
.B1(n_248),
.B2(n_253),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_221),
.B(n_210),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_268),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_193),
.C(n_189),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_163),
.C(n_166),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_159),
.C(n_170),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_260),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_248),
.B1(n_159),
.B2(n_2),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_275),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_4),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_281),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_267),
.B1(n_268),
.B2(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_5),
.Y(n_284)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_270),
.C(n_281),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_290),
.B(n_287),
.Y(n_291)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_277),
.C(n_283),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_287),
.B(n_285),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_272),
.C(n_271),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_6),
.B(n_10),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_11),
.C(n_12),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_11),
.B(n_12),
.Y(n_296)
);


endmodule