module fake_jpeg_19464_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_4),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_7),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_26),
.B(n_12),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_11),
.B(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_32),
.B(n_3),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_26),
.B1(n_21),
.B2(n_22),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_41)
);

AOI31xp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_12),
.A3(n_15),
.B(n_16),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_16),
.C(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_18),
.B1(n_4),
.B2(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_30),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_31),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_28),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_46),
.C(n_32),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_34),
.C(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_46),
.C(n_44),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_42),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_31),
.B(n_3),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

AO221x1_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_6),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.Y(n_60)
);


endmodule