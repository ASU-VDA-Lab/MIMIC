module fake_ariane_70_n_1703 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1703);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1703;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_17),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_43),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_74),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_52),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_59),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_41),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_34),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_35),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_82),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_66),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_22),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_95),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_58),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_90),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_39),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_51),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_40),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_44),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_57),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_89),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_41),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_15),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_105),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_107),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_18),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_47),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_119),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_28),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_20),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_56),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_53),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_48),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_0),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_68),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_65),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_72),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_13),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_24),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_35),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_20),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_34),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_153),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_93),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_106),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_64),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_137),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_103),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_27),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_7),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_11),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_39),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_99),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_127),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_108),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_4),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_122),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_30),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_83),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_70),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_32),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_146),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_12),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_22),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_100),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_15),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_152),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_102),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_85),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_61),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_126),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_50),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_71),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_11),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_139),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_10),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_117),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_26),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_8),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_9),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_79),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_44),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_1),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_128),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_76),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_37),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_46),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_135),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_18),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_148),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_88),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_150),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_3),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_91),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_4),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_55),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_125),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_104),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_21),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_45),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_33),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_10),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_145),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_33),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_84),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_157),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_168),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_305),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_157),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_164),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_176),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_259),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_216),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_159),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_267),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_163),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_273),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_159),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_304),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_198),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_189),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_164),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_190),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_191),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_190),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_193),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_259),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_193),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_163),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_167),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_167),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_239),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_239),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_178),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_181),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_201),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_202),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_194),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_215),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_225),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_169),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_207),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_194),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_226),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_257),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_210),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_212),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_277),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_281),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_283),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_286),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_165),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_218),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_296),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_228),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_299),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_229),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_236),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_253),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_230),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_158),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_172),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_232),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_242),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_179),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_268),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_171),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_217),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_315),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_332),
.B(n_206),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_339),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_319),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_217),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_325),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_326),
.A2(n_169),
.B1(n_285),
.B2(n_306),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_301),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_301),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_316),
.B(n_180),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_263),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_342),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_317),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_321),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_375),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_337),
.B(n_192),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_314),
.B(n_196),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

CKINVDCx8_ASAP7_75t_R g421 ( 
.A(n_374),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_320),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_348),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_346),
.B(n_171),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_334),
.B(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_351),
.Y(n_430)
);

NAND2x1_ASAP7_75t_L g431 ( 
.A(n_377),
.B(n_291),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_314),
.B(n_200),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_245),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_360),
.B(n_171),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_220),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_381),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_310),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_310),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_233),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_362),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_383),
.B(n_291),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_311),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

BUFx8_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_368),
.B(n_291),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_371),
.B(n_213),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_313),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_374),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_389),
.A2(n_424),
.B1(n_452),
.B2(n_436),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_385),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_409),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_439),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

INVx8_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_439),
.B(n_451),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_439),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_424),
.B(n_436),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_452),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_409),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_445),
.B(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_372),
.Y(n_474)
);

INVxp67_ASAP7_75t_R g475 ( 
.A(n_399),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_416),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_394),
.B(n_384),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_446),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_356),
.B1(n_322),
.B2(n_344),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_379),
.C(n_376),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_409),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_208),
.Y(n_482)
);

CKINVDCx6p67_ASAP7_75t_R g483 ( 
.A(n_448),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_394),
.B(n_380),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_419),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_429),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_429),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_446),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_442),
.B(n_223),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_411),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_352),
.Y(n_491)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_450),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_394),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_352),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_429),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_407),
.B(n_208),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_394),
.B(n_354),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_429),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_429),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_404),
.B(n_224),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_404),
.B(n_227),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_449),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_404),
.B(n_407),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_418),
.B(n_237),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_388),
.B(n_354),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_398),
.B(n_208),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_395),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_413),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_393),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_401),
.B(n_355),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_401),
.A2(n_244),
.B1(n_231),
.B2(n_213),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_396),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_393),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_435),
.A2(n_276),
.B1(n_252),
.B2(n_254),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_400),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_399),
.B(n_373),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_405),
.A2(n_188),
.B1(n_289),
.B2(n_282),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_400),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_402),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_401),
.B(n_238),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_400),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_422),
.B(n_177),
.C(n_175),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_406),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_401),
.B(n_248),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_406),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_408),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_440),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_438),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_398),
.B(n_426),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_408),
.Y(n_542)
);

BUFx6f_ASAP7_75t_SL g543 ( 
.A(n_421),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_410),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_410),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_386),
.A2(n_175),
.B1(n_306),
.B2(n_303),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_412),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_398),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_450),
.B(n_355),
.Y(n_552)
);

NOR2x1p5_ASAP7_75t_L g553 ( 
.A(n_421),
.B(n_177),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_386),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_450),
.A2(n_213),
.B1(n_293),
.B2(n_231),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_426),
.B(n_208),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_412),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_450),
.B(n_256),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_414),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_387),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_390),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_417),
.B(n_359),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_390),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_425),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_426),
.B(n_359),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_414),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_415),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_415),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_441),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_431),
.A2(n_278),
.B1(n_292),
.B2(n_289),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_420),
.B(n_265),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_434),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_431),
.A2(n_278),
.B1(n_188),
.B2(n_186),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_423),
.Y(n_578)
);

CKINVDCx6p67_ASAP7_75t_R g579 ( 
.A(n_437),
.Y(n_579)
);

AND3x1_ASAP7_75t_L g580 ( 
.A(n_453),
.B(n_373),
.C(n_369),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_423),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_387),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_428),
.B(n_269),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_428),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_453),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_392),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_392),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_403),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_403),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_432),
.B(n_363),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_432),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_409),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_447),
.B(n_363),
.Y(n_593)
);

BUFx16f_ASAP7_75t_R g594 ( 
.A(n_421),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_409),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_444),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_409),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_451),
.B(n_364),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_409),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_409),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_593),
.B(n_270),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_541),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_566),
.B(n_183),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_454),
.B(n_183),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_541),
.B(n_271),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_554),
.B(n_466),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_472),
.B(n_285),
.C(n_282),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_468),
.B(n_186),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_469),
.A2(n_231),
.B1(n_293),
.B2(n_233),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_469),
.B(n_160),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_457),
.B(n_293),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_460),
.A2(n_240),
.B(n_162),
.C(n_272),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_456),
.B(n_160),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_476),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_460),
.B(n_161),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_484),
.B(n_292),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_463),
.A2(n_369),
.B(n_366),
.C(n_365),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_507),
.B(n_303),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_457),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_463),
.A2(n_467),
.B1(n_493),
.B2(n_508),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_485),
.B(n_294),
.Y(n_622)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_479),
.A2(n_274),
.B1(n_264),
.B2(n_262),
.C(n_261),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_467),
.B(n_505),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_507),
.B(n_579),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_495),
.B(n_491),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_462),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_464),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_590),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_599),
.B(n_280),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_523),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_585),
.B(n_161),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_535),
.B(n_166),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_562),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_562),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_510),
.B(n_364),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_455),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_493),
.A2(n_234),
.B1(n_309),
.B2(n_307),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_535),
.B(n_462),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_535),
.B(n_166),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_505),
.Y(n_643)
);

AO22x2_ASAP7_75t_L g644 ( 
.A1(n_560),
.A2(n_366),
.B1(n_329),
.B2(n_328),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_582),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_505),
.B(n_302),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_563),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_582),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_551),
.B(n_234),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_551),
.B(n_170),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_563),
.B(n_313),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_582),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_565),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_491),
.B(n_318),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_462),
.B(n_480),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_462),
.B(n_318),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_506),
.A2(n_174),
.B1(n_309),
.B2(n_307),
.Y(n_657)
);

INVx8_ASAP7_75t_L g658 ( 
.A(n_543),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_565),
.B(n_323),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_595),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_472),
.B(n_247),
.C(n_246),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_489),
.A2(n_260),
.B1(n_328),
.B2(n_327),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_580),
.B(n_170),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_523),
.A2(n_173),
.B1(n_187),
.B2(n_185),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_597),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_551),
.B(n_173),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_501),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_501),
.B(n_174),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_323),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_516),
.B(n_517),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_516),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_517),
.B(n_182),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_552),
.B(n_182),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_521),
.B(n_184),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_486),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_513),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_526),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_486),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_486),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_526),
.B(n_184),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_519),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_520),
.B(n_185),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_530),
.B(n_537),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

OR2x6_ASAP7_75t_L g686 ( 
.A(n_523),
.B(n_324),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_564),
.B(n_187),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_579),
.B(n_279),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_L g689 ( 
.A(n_474),
.B(n_279),
.C(n_284),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_498),
.B(n_284),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_547),
.B(n_287),
.Y(n_691)
);

NAND2x1p5_ASAP7_75t_L g692 ( 
.A(n_559),
.B(n_324),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_574),
.B(n_287),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_514),
.B(n_288),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_537),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_477),
.B(n_288),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_522),
.B(n_290),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_525),
.Y(n_698)
);

INVxp67_ASAP7_75t_SL g699 ( 
.A(n_486),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_538),
.B(n_290),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_577),
.B(n_555),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_515),
.B(n_300),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_465),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_538),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_567),
.A2(n_329),
.B(n_327),
.C(n_3),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_539),
.B(n_300),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_556),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_523),
.B(n_474),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_532),
.A2(n_221),
.B(n_275),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_556),
.B(n_219),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_511),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_475),
.A2(n_568),
.B1(n_572),
.B2(n_550),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_571),
.B(n_214),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_490),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_571),
.B(n_222),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_559),
.B(n_211),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_573),
.B(n_241),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_573),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_586),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_534),
.A2(n_0),
.B(n_2),
.C(n_7),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_542),
.B(n_209),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_506),
.B(n_195),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_545),
.B(n_546),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_560),
.B(n_531),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_558),
.B(n_243),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_553),
.B(n_8),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_502),
.B(n_199),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_561),
.B(n_249),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_543),
.Y(n_731)
);

OAI21xp33_ASAP7_75t_L g732 ( 
.A1(n_569),
.A2(n_250),
.B(n_266),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_570),
.B(n_203),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_483),
.B(n_489),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_476),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_586),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_465),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_578),
.B(n_258),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_528),
.A2(n_251),
.B1(n_205),
.B2(n_204),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_594),
.B(n_295),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_502),
.B(n_12),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_581),
.Y(n_742)
);

AOI221xp5_ASAP7_75t_L g743 ( 
.A1(n_524),
.A2(n_295),
.B1(n_208),
.B2(n_19),
.C(n_23),
.Y(n_743)
);

BUFx5_ASAP7_75t_L g744 ( 
.A(n_482),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_503),
.B(n_14),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_483),
.B(n_14),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_587),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_584),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_528),
.A2(n_295),
.B1(n_19),
.B2(n_25),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_471),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_503),
.B(n_533),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_490),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_575),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_575),
.B(n_16),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_533),
.B(n_16),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_473),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_559),
.B(n_295),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_478),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_559),
.B(n_295),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_588),
.B(n_25),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_583),
.B(n_26),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_488),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_591),
.B(n_589),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_504),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_583),
.B(n_27),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_543),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_559),
.B(n_29),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_587),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_512),
.B(n_31),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_627),
.Y(n_770)
);

O2A1O1Ixp5_ASAP7_75t_L g771 ( 
.A1(n_602),
.A2(n_601),
.B(n_600),
.C(n_536),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_667),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_605),
.B(n_601),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_658),
.B(n_492),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_R g775 ( 
.A(n_620),
.B(n_492),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_627),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_626),
.B(n_601),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_701),
.A2(n_497),
.B1(n_482),
.B2(n_492),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_735),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_589),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_664),
.B(n_497),
.C(n_509),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_638),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_627),
.B(n_592),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_R g784 ( 
.A(n_713),
.B(n_716),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_671),
.Y(n_785)
);

AND3x1_ASAP7_75t_L g786 ( 
.A(n_612),
.B(n_600),
.C(n_536),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_741),
.A2(n_482),
.B1(n_598),
.B2(n_596),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_615),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_752),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_741),
.A2(n_482),
.B1(n_598),
.B2(n_596),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_603),
.B(n_600),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_656),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_660),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_607),
.B(n_592),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_665),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_710),
.B(n_714),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_714),
.B(n_592),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_658),
.Y(n_798)
);

BUFx12f_ASAP7_75t_L g799 ( 
.A(n_740),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_658),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_676),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_680),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_675),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_602),
.B(n_465),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_725),
.B(n_470),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_625),
.B(n_592),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_682),
.Y(n_807)
);

AND2x6_ASAP7_75t_L g808 ( 
.A(n_745),
.B(n_499),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_653),
.Y(n_809)
);

CKINVDCx11_ASAP7_75t_R g810 ( 
.A(n_740),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_651),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_698),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_647),
.B(n_470),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_725),
.B(n_470),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_659),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_704),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_677),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_742),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_675),
.Y(n_819)
);

AND3x1_ASAP7_75t_SL g820 ( 
.A(n_623),
.B(n_36),
.C(n_37),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_748),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_675),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_678),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_626),
.B(n_496),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_664),
.A2(n_482),
.B1(n_496),
.B2(n_529),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_637),
.B(n_482),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_619),
.A2(n_496),
.B1(n_529),
.B2(n_536),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_745),
.A2(n_500),
.B1(n_549),
.B2(n_548),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_750),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_686),
.B(n_500),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_756),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_728),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_751),
.B(n_529),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_606),
.B(n_499),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_606),
.B(n_494),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_622),
.B(n_494),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_614),
.A2(n_458),
.B1(n_549),
.B2(n_548),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_622),
.B(n_487),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_669),
.B(n_487),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_624),
.A2(n_481),
.B(n_544),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_758),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_726),
.B(n_481),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_762),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_686),
.B(n_656),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_644),
.A2(n_755),
.B1(n_631),
.B2(n_765),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_SL g846 ( 
.A1(n_624),
.A2(n_540),
.B(n_459),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_617),
.A2(n_609),
.B(n_754),
.C(n_630),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_764),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_678),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_643),
.B(n_544),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_643),
.B(n_540),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_656),
.Y(n_852)
);

AND2x4_ASAP7_75t_SL g853 ( 
.A(n_734),
.B(n_461),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_670),
.B(n_461),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_628),
.B(n_459),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_688),
.B(n_458),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_695),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_670),
.B(n_557),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_684),
.B(n_557),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_644),
.A2(n_509),
.B1(n_42),
.B2(n_43),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_644),
.A2(n_631),
.B1(n_761),
.B2(n_724),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_654),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_684),
.B(n_38),
.Y(n_863)
);

NOR2x1p5_ASAP7_75t_L g864 ( 
.A(n_632),
.B(n_38),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_654),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_753),
.B(n_49),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_678),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_679),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_705),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_679),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_679),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_731),
.B(n_766),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_768),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_634),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_604),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_629),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_708),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_709),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_720),
.B(n_69),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_729),
.A2(n_86),
.B1(n_96),
.B2(n_98),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_746),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_721),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_646),
.B(n_101),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_763),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_663),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_760),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_736),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_760),
.Y(n_888)
);

INVx6_ASAP7_75t_L g889 ( 
.A(n_769),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_747),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_646),
.B(n_109),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_641),
.B(n_110),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_618),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_691),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_689),
.B(n_124),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_668),
.A2(n_133),
.B(n_143),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_633),
.A2(n_154),
.B1(n_155),
.B2(n_642),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_635),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_702),
.B(n_611),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_703),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_668),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_650),
.B(n_666),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_636),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_743),
.A2(n_749),
.B(n_730),
.C(n_738),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_723),
.A2(n_730),
.B(n_738),
.C(n_727),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_661),
.B(n_655),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_SL g908 ( 
.A1(n_687),
.A2(n_723),
.B1(n_727),
.B2(n_610),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_672),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_SL g910 ( 
.A(n_608),
.B(n_639),
.C(n_722),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_645),
.Y(n_911)
);

NOR2x2_ASAP7_75t_L g912 ( 
.A(n_693),
.B(n_683),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_616),
.B(n_673),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_650),
.B(n_666),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_672),
.A2(n_700),
.B1(n_707),
.B2(n_681),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_648),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_692),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_674),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_652),
.B(n_640),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_674),
.A2(n_700),
.B1(n_707),
.B2(n_681),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_657),
.B(n_697),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_692),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_690),
.A2(n_694),
.B1(n_732),
.B2(n_696),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_739),
.A2(n_733),
.B1(n_737),
.B2(n_649),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_649),
.A2(n_613),
.B(n_706),
.C(n_717),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_712),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_767),
.Y(n_927)
);

AND2x4_ASAP7_75t_SL g928 ( 
.A(n_662),
.B(n_744),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_757),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_744),
.B(n_711),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_712),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_744),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_715),
.B(n_717),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_715),
.B(n_719),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_719),
.B(n_699),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_744),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_718),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_759),
.A2(n_605),
.B(n_602),
.C(n_664),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_744),
.B(n_603),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_603),
.B(n_602),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_735),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_627),
.B(n_641),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_SL g943 ( 
.A1(n_612),
.A2(n_664),
.B1(n_710),
.B2(n_631),
.Y(n_943)
);

BUFx4f_ASAP7_75t_L g944 ( 
.A(n_658),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_638),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_605),
.A2(n_701),
.B1(n_710),
.B2(n_714),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_627),
.Y(n_947)
);

AO22x1_ASAP7_75t_L g948 ( 
.A1(n_713),
.A2(n_457),
.B1(n_511),
.B2(n_315),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_627),
.B(n_621),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_782),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_875),
.B(n_940),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_847),
.A2(n_938),
.B(n_905),
.C(n_906),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_774),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_798),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_792),
.B(n_775),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_788),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_940),
.B(n_946),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_811),
.A2(n_815),
.B(n_921),
.C(n_910),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_862),
.B(n_902),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_909),
.A2(n_918),
.B(n_933),
.C(n_925),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_784),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_774),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_803),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_774),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_796),
.B(n_948),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_SL g966 ( 
.A1(n_773),
.A2(n_913),
.B(n_920),
.C(n_915),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_876),
.B(n_884),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_865),
.B(n_839),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_792),
.B(n_908),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_809),
.A2(n_808),
.B1(n_889),
.B2(n_943),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_886),
.A2(n_924),
.B1(n_923),
.B2(n_934),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_891),
.A2(n_933),
.B(n_804),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_944),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_944),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_800),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_901),
.B(n_792),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_926),
.B(n_931),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_810),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_792),
.B(n_786),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_799),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_885),
.A2(n_824),
.B(n_794),
.C(n_813),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_900),
.A2(n_888),
.B(n_781),
.C(n_896),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_832),
.B(n_779),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_805),
.A2(n_814),
.B1(n_804),
.B2(n_945),
.Y(n_984)
);

OAI22x1_ASAP7_75t_L g985 ( 
.A1(n_864),
.A2(n_852),
.B1(n_927),
.B2(n_881),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_883),
.A2(n_814),
.B(n_805),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_785),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_855),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_793),
.B(n_795),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_780),
.B(n_770),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_801),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_802),
.B(n_807),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_824),
.A2(n_941),
.B(n_789),
.C(n_863),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_896),
.A2(n_897),
.B(n_863),
.C(n_893),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_812),
.B(n_816),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_818),
.B(n_821),
.Y(n_996)
);

OAI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_860),
.A2(n_833),
.B(n_939),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_771),
.A2(n_833),
.B(n_840),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_844),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_844),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_844),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_873),
.A2(n_791),
.B(n_841),
.C(n_848),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_770),
.B(n_777),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_907),
.A2(n_935),
.B(n_949),
.C(n_873),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_808),
.B(n_826),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_834),
.A2(n_835),
.B(n_935),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_777),
.B(n_830),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_889),
.B(n_829),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_770),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_872),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_907),
.A2(n_838),
.B(n_836),
.C(n_939),
.Y(n_1011)
);

NOR2xp67_ASAP7_75t_L g1012 ( 
.A(n_901),
.B(n_776),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_SL g1013 ( 
.A1(n_932),
.A2(n_836),
.B(n_838),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_817),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_901),
.B(n_819),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_901),
.B(n_872),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_831),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_803),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_898),
.B(n_843),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_882),
.Y(n_1020)
);

AO22x1_ASAP7_75t_L g1021 ( 
.A1(n_808),
.A2(n_947),
.B1(n_868),
.B2(n_917),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_808),
.B(n_853),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_861),
.B(n_845),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_834),
.A2(n_835),
.B(n_930),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_791),
.A2(n_895),
.B(n_856),
.C(n_892),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_830),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_830),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_842),
.B(n_904),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_887),
.Y(n_1029)
);

AND3x1_ASAP7_75t_SL g1030 ( 
.A(n_912),
.B(n_820),
.C(n_898),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_904),
.B(n_787),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_858),
.A2(n_859),
.B(n_840),
.Y(n_1032)
);

OA22x2_ASAP7_75t_L g1033 ( 
.A1(n_825),
.A2(n_778),
.B1(n_911),
.B2(n_916),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_858),
.A2(n_859),
.B(n_854),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_857),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_874),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_890),
.A2(n_877),
.B1(n_878),
.B2(n_869),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_854),
.A2(n_850),
.B(n_851),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_797),
.A2(n_846),
.B(n_851),
.C(n_850),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_SL g1040 ( 
.A1(n_790),
.A2(n_894),
.B1(n_880),
.B2(n_942),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_874),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_819),
.B(n_867),
.Y(n_1042)
);

OAI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_827),
.A2(n_828),
.B(n_942),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_937),
.A2(n_879),
.B(n_866),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_837),
.A2(n_937),
.B(n_866),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_874),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_822),
.A2(n_867),
.B1(n_871),
.B2(n_823),
.Y(n_1047)
);

AND2x6_ASAP7_75t_L g1048 ( 
.A(n_922),
.B(n_871),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_806),
.B(n_783),
.C(n_822),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_823),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_928),
.A2(n_879),
.B(n_936),
.C(n_929),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_899),
.B(n_849),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_899),
.A2(n_919),
.B1(n_929),
.B2(n_870),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_919),
.A2(n_870),
.B(n_871),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_929),
.A2(n_605),
.B1(n_457),
.B2(n_946),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_903),
.A2(n_914),
.B(n_891),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_946),
.A2(n_938),
.B(n_847),
.C(n_605),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_772),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_840),
.A2(n_879),
.B(n_771),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_SL g1060 ( 
.A1(n_906),
.A2(n_847),
.B(n_914),
.C(n_903),
.Y(n_1060)
);

AO32x2_ASAP7_75t_L g1061 ( 
.A1(n_873),
.A2(n_714),
.A3(n_664),
.B1(n_753),
.B2(n_876),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_847),
.A2(n_605),
.B(n_875),
.C(n_602),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_946),
.A2(n_602),
.B1(n_847),
.B2(n_875),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_811),
.B(n_815),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_811),
.B(n_815),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_903),
.A2(n_914),
.B(n_891),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_844),
.B(n_798),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_875),
.B(n_315),
.Y(n_1068)
);

AO21x2_ASAP7_75t_L g1069 ( 
.A1(n_906),
.A2(n_914),
.B(n_903),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_784),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_875),
.B(n_593),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_774),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_903),
.A2(n_914),
.B(n_891),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_875),
.B(n_593),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_847),
.A2(n_605),
.B(n_875),
.C(n_602),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_798),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_782),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_946),
.A2(n_602),
.B1(n_847),
.B2(n_875),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_784),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_875),
.B(n_593),
.Y(n_1080)
);

INVx11_ASAP7_75t_L g1081 ( 
.A(n_799),
.Y(n_1081)
);

AND2x6_ASAP7_75t_L g1082 ( 
.A(n_932),
.B(n_627),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_903),
.A2(n_914),
.B(n_891),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_772),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_875),
.B(n_593),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_774),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_903),
.A2(n_914),
.B(n_891),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_950),
.Y(n_1088)
);

BUFx4_ASAP7_75t_SL g1089 ( 
.A(n_961),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_1079),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_1070),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_1055),
.B(n_957),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1071),
.B(n_1074),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1063),
.B(n_1078),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1080),
.B(n_1085),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_SL g1097 ( 
.A(n_954),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_953),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1057),
.A2(n_1075),
.B1(n_1062),
.B2(n_994),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_991),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_972),
.A2(n_986),
.B(n_984),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_965),
.B(n_971),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_977),
.B(n_960),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1017),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1082),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_998),
.A2(n_1034),
.B(n_1044),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_975),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_952),
.A2(n_982),
.B(n_1004),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_1081),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1056),
.A2(n_1073),
.B(n_1066),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_951),
.B(n_1064),
.Y(n_1111)
);

BUFx8_ASAP7_75t_L g1112 ( 
.A(n_973),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1077),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1065),
.B(n_1068),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_988),
.B(n_970),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1008),
.B(n_967),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1083),
.A2(n_1087),
.B(n_1038),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1006),
.A2(n_1045),
.B(n_1039),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_953),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_L g1120 ( 
.A(n_1054),
.B(n_999),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1011),
.A2(n_1051),
.B(n_1043),
.Y(n_1121)
);

AO22x2_ASAP7_75t_L g1122 ( 
.A1(n_1023),
.A2(n_969),
.B1(n_1061),
.B2(n_979),
.Y(n_1122)
);

AND2x2_ASAP7_75t_SL g1123 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1013),
.A2(n_1060),
.B(n_1002),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_968),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1033),
.A2(n_1025),
.B(n_993),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_997),
.A2(n_958),
.B(n_966),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_999),
.B(n_1050),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1040),
.A2(n_1069),
.B(n_1028),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_997),
.B(n_981),
.C(n_1019),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1005),
.A2(n_1047),
.B(n_1053),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_1076),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_973),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1010),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1031),
.A2(n_1058),
.A3(n_1014),
.B(n_1084),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_973),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1069),
.A2(n_995),
.B(n_989),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1046),
.A2(n_976),
.B(n_1016),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_953),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_992),
.A2(n_996),
.B(n_959),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1020),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_976),
.B(n_1086),
.Y(n_1142)
);

INVx5_ASAP7_75t_L g1143 ( 
.A(n_974),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_999),
.B(n_1000),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1029),
.B(n_1035),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1022),
.A2(n_990),
.B(n_963),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1015),
.A2(n_1012),
.B(n_1052),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_987),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_L g1149 ( 
.A(n_1003),
.B(n_955),
.C(n_983),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_962),
.B(n_1086),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_962),
.B(n_1086),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1026),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1021),
.A2(n_1015),
.B(n_1042),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1041),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1012),
.A2(n_1037),
.B(n_1042),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_974),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1036),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_962),
.B(n_964),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1027),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1048),
.B(n_1082),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1061),
.A2(n_985),
.A3(n_1030),
.B(n_1049),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1018),
.A2(n_1067),
.B(n_1061),
.Y(n_1162)
);

INVx5_ASAP7_75t_L g1163 ( 
.A(n_974),
.Y(n_1163)
);

INVx3_ASAP7_75t_SL g1164 ( 
.A(n_978),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_1067),
.A2(n_1082),
.B(n_1018),
.C(n_1009),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1018),
.A2(n_1009),
.B(n_964),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_964),
.B(n_1072),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1048),
.B(n_1072),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1009),
.A2(n_1048),
.B(n_980),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1063),
.A2(n_1078),
.B(n_1057),
.C(n_605),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1082),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_956),
.Y(n_1175)
);

INVx3_ASAP7_75t_SL g1176 ( 
.A(n_961),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1082),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_950),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_1057),
.A2(n_1078),
.B(n_1063),
.C(n_994),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_994),
.A2(n_1044),
.A3(n_972),
.B(n_1006),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_R g1184 ( 
.A(n_961),
.B(n_620),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_968),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1010),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1059),
.A2(n_998),
.B(n_1044),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1189)
);

INVxp67_ASAP7_75t_SL g1190 ( 
.A(n_968),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_956),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_994),
.A2(n_1044),
.A3(n_972),
.B(n_1006),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1063),
.A2(n_946),
.B1(n_1078),
.B2(n_605),
.Y(n_1197)
);

AOI211x1_ASAP7_75t_L g1198 ( 
.A1(n_1063),
.A2(n_1078),
.B(n_910),
.C(n_714),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_999),
.B(n_1007),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_SL g1200 ( 
.A1(n_952),
.A2(n_1078),
.B(n_1063),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_957),
.B(n_1063),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_961),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_957),
.A2(n_1057),
.B1(n_946),
.B2(n_1063),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_950),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_994),
.A2(n_1044),
.A3(n_972),
.B(n_1006),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_951),
.B(n_615),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_953),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_SL g1210 ( 
.A1(n_957),
.A2(n_1057),
.B(n_1011),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_957),
.B(n_1063),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_957),
.B(n_1063),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1213)
);

O2A1O1Ixp5_ASAP7_75t_SL g1214 ( 
.A1(n_969),
.A2(n_1078),
.B(n_1063),
.C(n_971),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_972),
.A2(n_986),
.B(n_994),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_968),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_961),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_965),
.A2(n_970),
.B1(n_946),
.B2(n_710),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_957),
.B(n_1063),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_950),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1059),
.A2(n_998),
.B(n_1044),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_999),
.B(n_1007),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1032),
.A2(n_1024),
.B(n_1059),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_957),
.B(n_1063),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1174),
.A2(n_1192),
.B(n_1179),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_1197),
.B(n_1171),
.C(n_1102),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1109),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1089),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1088),
.Y(n_1230)
);

AOI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1200),
.A2(n_1195),
.B1(n_1201),
.B2(n_1202),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1129),
.A2(n_1137),
.A3(n_1124),
.B(n_1099),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1100),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1095),
.A2(n_1173),
.B(n_1170),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1213),
.A2(n_1215),
.B(n_1101),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1199),
.B(n_1223),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1106),
.A2(n_1180),
.B(n_1177),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1183),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1185),
.A2(n_1196),
.B(n_1224),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1189),
.A2(n_1194),
.B(n_1217),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1104),
.Y(n_1242)
);

AO21x2_ASAP7_75t_L g1243 ( 
.A1(n_1127),
.A2(n_1197),
.B(n_1162),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1113),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1117),
.A2(n_1110),
.B(n_1118),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1181),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1091),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1112),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1132),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1126),
.A2(n_1182),
.B(n_1222),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1206),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1108),
.A2(n_1094),
.B(n_1205),
.C(n_1127),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1188),
.A2(n_1222),
.B(n_1108),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1094),
.A2(n_1103),
.B(n_1140),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1221),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1105),
.B(n_1172),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1112),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1188),
.A2(n_1131),
.B(n_1099),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1198),
.A2(n_1115),
.B1(n_1164),
.B2(n_1114),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1214),
.A2(n_1205),
.B(n_1210),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1141),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1198),
.A2(n_1225),
.B1(n_1203),
.B2(n_1220),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1155),
.A2(n_1225),
.B(n_1211),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1203),
.A2(n_1212),
.B(n_1220),
.C(n_1211),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1183),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1218),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1172),
.B(n_1178),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1107),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1212),
.A2(n_1103),
.B(n_1130),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1090),
.Y(n_1270)
);

BUFx12f_ASAP7_75t_L g1271 ( 
.A(n_1204),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1145),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1145),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1218),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1219),
.A2(n_1092),
.B1(n_1130),
.B2(n_1122),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1140),
.A2(n_1153),
.B(n_1186),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1208),
.A2(n_1125),
.B(n_1190),
.C(n_1216),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1147),
.A2(n_1146),
.B(n_1138),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1148),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1176),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1121),
.A2(n_1160),
.B(n_1165),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1199),
.B(n_1223),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1121),
.A2(n_1160),
.B(n_1183),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1193),
.A2(n_1207),
.B(n_1122),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1175),
.A2(n_1191),
.B(n_1149),
.C(n_1152),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1175),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_SL g1287 ( 
.A1(n_1169),
.A2(n_1166),
.B(n_1168),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1187),
.B(n_1154),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1120),
.A2(n_1168),
.B(n_1142),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1157),
.B(n_1134),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1159),
.B(n_1161),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_SL g1292 ( 
.A1(n_1133),
.A2(n_1136),
.B(n_1156),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1098),
.B(n_1209),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1098),
.B(n_1209),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1161),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1151),
.A2(n_1158),
.B(n_1128),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1144),
.B(n_1128),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1161),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1207),
.A2(n_1144),
.B(n_1123),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1133),
.A2(n_1143),
.B(n_1163),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1119),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1143),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1167),
.A2(n_1150),
.B(n_1139),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1143),
.A2(n_1163),
.B(n_1209),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_SL g1305 ( 
.A(n_1184),
.B(n_1097),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1167),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_R g1307 ( 
.A(n_1109),
.B(n_961),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1095),
.A2(n_1173),
.B(n_1170),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1088),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1095),
.A2(n_1173),
.B(n_1170),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1112),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1088),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1088),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1112),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1112),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1095),
.A2(n_1173),
.B(n_1170),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1135),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1197),
.A2(n_1171),
.B(n_946),
.C(n_1075),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1102),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1102),
.A2(n_1023),
.B1(n_861),
.B2(n_845),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1112),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1093),
.B(n_1096),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1135),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1088),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1111),
.B(n_1116),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1171),
.A2(n_1094),
.B(n_1101),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1171),
.A2(n_1094),
.B(n_1101),
.Y(n_1330)
);

NAND2xp33_ASAP7_75t_L g1331 ( 
.A(n_1197),
.B(n_1094),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1088),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_SL g1333 ( 
.A1(n_1171),
.A2(n_1197),
.B(n_1200),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1095),
.A2(n_1173),
.B(n_1170),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_1094),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1088),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1095),
.A2(n_1173),
.B(n_1170),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1199),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1174),
.A2(n_1192),
.B(n_1179),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1197),
.A2(n_1171),
.B(n_946),
.C(n_1075),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1171),
.A2(n_1094),
.B(n_1101),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1174),
.A2(n_1192),
.B(n_1179),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1284),
.A2(n_1258),
.B(n_1238),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1315),
.B(n_1286),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1290),
.B(n_1328),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1288),
.B(n_1230),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1252),
.A2(n_1227),
.B(n_1269),
.C(n_1321),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1331),
.A2(n_1330),
.B(n_1329),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1252),
.A2(n_1321),
.B1(n_1340),
.B2(n_1320),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1341),
.A2(n_1331),
.B(n_1335),
.C(n_1264),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1340),
.A2(n_1333),
.B(n_1264),
.C(n_1322),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1234),
.B(n_1242),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1257),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1249),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1244),
.B(n_1246),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1307),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1262),
.A2(n_1322),
.B(n_1335),
.C(n_1266),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1238),
.A2(n_1245),
.B(n_1283),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1251),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1233),
.A2(n_1313),
.B(n_1325),
.C(n_1277),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1260),
.A2(n_1275),
.B(n_1277),
.C(n_1323),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1259),
.B(n_1254),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1253),
.A2(n_1250),
.B(n_1337),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1255),
.B(n_1309),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1237),
.B(n_1282),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1254),
.B(n_1272),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1312),
.B(n_1314),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_SL g1368 ( 
.A1(n_1239),
.A2(n_1265),
.B(n_1294),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1274),
.B(n_1268),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1260),
.A2(n_1275),
.B(n_1323),
.C(n_1285),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1237),
.B(n_1282),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1249),
.A2(n_1231),
.B1(n_1302),
.B2(n_1247),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1327),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1235),
.A2(n_1241),
.B(n_1318),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1332),
.B(n_1336),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1273),
.B(n_1261),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1279),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1308),
.A2(n_1334),
.B(n_1310),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1291),
.B(n_1243),
.Y(n_1379)
);

OAI31xp33_ASAP7_75t_L g1380 ( 
.A1(n_1295),
.A2(n_1298),
.A3(n_1305),
.B(n_1267),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1243),
.B(n_1293),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1276),
.B(n_1301),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1236),
.A2(n_1226),
.B(n_1339),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1300),
.A2(n_1297),
.B(n_1299),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1263),
.A2(n_1281),
.B(n_1278),
.Y(n_1385)
);

AOI221xp5_ASAP7_75t_L g1386 ( 
.A1(n_1248),
.A2(n_1324),
.B1(n_1317),
.B2(n_1257),
.C(n_1311),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1302),
.A2(n_1316),
.B1(n_1311),
.B2(n_1280),
.Y(n_1387)
);

BUFx4f_ASAP7_75t_SL g1388 ( 
.A(n_1228),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1316),
.A2(n_1280),
.B1(n_1268),
.B2(n_1267),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1299),
.B(n_1232),
.Y(n_1390)
);

AOI21x1_ASAP7_75t_SL g1391 ( 
.A1(n_1226),
.A2(n_1342),
.B(n_1339),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_SL g1392 ( 
.A1(n_1226),
.A2(n_1342),
.B(n_1339),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1338),
.B(n_1232),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1232),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_SL g1395 ( 
.A1(n_1342),
.A2(n_1236),
.B(n_1232),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1338),
.B(n_1256),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1306),
.A2(n_1236),
.B1(n_1229),
.B2(n_1270),
.Y(n_1397)
);

AOI221x1_ASAP7_75t_SL g1398 ( 
.A1(n_1270),
.A2(n_1271),
.B1(n_1229),
.B2(n_1228),
.C(n_1307),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1306),
.B(n_1304),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1271),
.A2(n_1292),
.B1(n_1240),
.B2(n_1326),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_L g1401 ( 
.A(n_1303),
.B(n_1319),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1240),
.A2(n_1319),
.B1(n_1287),
.B2(n_1296),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1296),
.B(n_1289),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1240),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1284),
.A2(n_1258),
.B(n_1238),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1227),
.A2(n_1197),
.B1(n_1252),
.B2(n_1094),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1307),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1233),
.B(n_1313),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1230),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1307),
.Y(n_1410)
);

NOR2xp67_ASAP7_75t_L g1411 ( 
.A(n_1322),
.B(n_1266),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1331),
.A2(n_1094),
.B(n_1171),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1227),
.A2(n_1197),
.B1(n_1252),
.B2(n_1094),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1252),
.A2(n_965),
.B(n_1171),
.C(n_1197),
.Y(n_1414)
);

NOR2x1_ASAP7_75t_SL g1415 ( 
.A(n_1254),
.B(n_1102),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1233),
.B(n_1313),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1233),
.B(n_1313),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1230),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1233),
.B(n_1313),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1366),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1349),
.A2(n_1406),
.B1(n_1413),
.B2(n_1412),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1348),
.B(n_1412),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1404),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1394),
.B(n_1385),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1383),
.A2(n_1348),
.B(n_1361),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1350),
.B(n_1415),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_SL g1428 ( 
.A1(n_1347),
.A2(n_1414),
.B(n_1351),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1383),
.A2(n_1403),
.B(n_1382),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1390),
.B(n_1343),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1384),
.B(n_1401),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1343),
.B(n_1405),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1374),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1350),
.A2(n_1370),
.B(n_1362),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1378),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1378),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1362),
.A2(n_1393),
.B(n_1381),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1359),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1373),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1409),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1360),
.B(n_1351),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1363),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1418),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1367),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1391),
.A2(n_1392),
.B(n_1395),
.Y(n_1447)
);

NOR2x1_ASAP7_75t_SL g1448 ( 
.A(n_1397),
.B(n_1372),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1402),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1352),
.B(n_1355),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1364),
.B(n_1375),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1360),
.B(n_1357),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1379),
.B(n_1346),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1376),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1408),
.A2(n_1419),
.B1(n_1416),
.B2(n_1417),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1400),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1391),
.A2(n_1392),
.B(n_1368),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1344),
.B(n_1345),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1365),
.B(n_1371),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_SL g1460 ( 
.A(n_1399),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1437),
.Y(n_1461)
);

AOI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1427),
.A2(n_1411),
.B(n_1389),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1437),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1430),
.B(n_1459),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1430),
.B(n_1396),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1421),
.A2(n_1428),
.B1(n_1443),
.B2(n_1452),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1420),
.B(n_1380),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1450),
.B(n_1451),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1420),
.B(n_1369),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1450),
.B(n_1451),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1453),
.B(n_1354),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1424),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1424),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1420),
.B(n_1454),
.Y(n_1474)
);

BUFx2_ASAP7_75t_SL g1475 ( 
.A(n_1424),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1456),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1454),
.B(n_1386),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1422),
.B(n_1353),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1476),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1461),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1461),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1476),
.Y(n_1484)
);

AOI31xp33_ASAP7_75t_L g1485 ( 
.A1(n_1466),
.A2(n_1443),
.A3(n_1421),
.B(n_1452),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1466),
.A2(n_1434),
.B1(n_1449),
.B2(n_1423),
.Y(n_1486)
);

AOI33xp33_ASAP7_75t_L g1487 ( 
.A1(n_1477),
.A2(n_1449),
.A3(n_1458),
.B1(n_1442),
.B2(n_1445),
.B3(n_1441),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1461),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1476),
.A2(n_1388),
.B1(n_1443),
.B2(n_1456),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1476),
.A2(n_1448),
.B1(n_1434),
.B2(n_1423),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1478),
.A2(n_1434),
.B1(n_1449),
.B2(n_1423),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1479),
.A2(n_1428),
.B1(n_1455),
.B2(n_1434),
.C(n_1452),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1468),
.B(n_1455),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1467),
.A2(n_1434),
.B(n_1435),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1478),
.A2(n_1422),
.B1(n_1427),
.B2(n_1455),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1462),
.A2(n_1457),
.B(n_1447),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1478),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1467),
.A2(n_1434),
.B(n_1433),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1478),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_L g1500 ( 
.A(n_1480),
.Y(n_1500)
);

NAND4xp25_ASAP7_75t_L g1501 ( 
.A(n_1477),
.B(n_1444),
.C(n_1398),
.D(n_1427),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1468),
.B(n_1453),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1468),
.Y(n_1503)
);

NAND4xp25_ASAP7_75t_L g1504 ( 
.A(n_1477),
.B(n_1444),
.C(n_1439),
.D(n_1386),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_1471),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1469),
.B(n_1429),
.C(n_1440),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1463),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1463),
.Y(n_1508)
);

AOI211xp5_ASAP7_75t_L g1509 ( 
.A1(n_1472),
.A2(n_1448),
.B(n_1387),
.C(n_1432),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1469),
.B(n_1429),
.C(n_1440),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1465),
.A2(n_1425),
.B1(n_1438),
.B2(n_1460),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1470),
.B(n_1446),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1464),
.B(n_1470),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1502),
.B(n_1472),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1492),
.B(n_1474),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1513),
.B(n_1472),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1482),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1488),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1494),
.A2(n_1425),
.B(n_1433),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1499),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1503),
.B(n_1473),
.Y(n_1521)
);

OR2x6_ASAP7_75t_L g1522 ( 
.A(n_1506),
.B(n_1431),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1482),
.Y(n_1523)
);

NAND2x1_ASAP7_75t_L g1524 ( 
.A(n_1497),
.B(n_1473),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1483),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1483),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1507),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1510),
.B(n_1431),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1496),
.A2(n_1426),
.B(n_1444),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1484),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1513),
.B(n_1464),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1499),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1493),
.B(n_1474),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1508),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1511),
.A2(n_1426),
.B(n_1436),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1523),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1515),
.B(n_1485),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1519),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1523),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1535),
.B(n_1504),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1526),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1531),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1526),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1519),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1516),
.B(n_1497),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1527),
.B(n_1481),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1509),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1515),
.B(n_1512),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1537),
.A2(n_1486),
.B1(n_1490),
.B2(n_1491),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1531),
.B(n_1487),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1521),
.B(n_1481),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1534),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1536),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_L g1556 ( 
.A(n_1520),
.B(n_1484),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1536),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1518),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1518),
.B(n_1494),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1517),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1514),
.B(n_1501),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1517),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1514),
.B(n_1494),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1514),
.B(n_1498),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1527),
.B(n_1500),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1534),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1517),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1498),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1530),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1525),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1539),
.B(n_1498),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1550),
.B(n_1525),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1565),
.B(n_1527),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1558),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_L g1575 ( 
.A(n_1556),
.B(n_1489),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1565),
.B(n_1527),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1549),
.B(n_1527),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1549),
.B(n_1527),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1561),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1558),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1553),
.B(n_1532),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1551),
.A2(n_1522),
.B1(n_1529),
.B2(n_1495),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1560),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_SL g1584 ( 
.A(n_1551),
.B(n_1524),
.C(n_1533),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1550),
.B(n_1525),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1560),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1562),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1567),
.Y(n_1589)
);

INVx3_ASAP7_75t_SL g1590 ( 
.A(n_1566),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1546),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1556),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1567),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1570),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1570),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1548),
.B(n_1532),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1547),
.B(n_1532),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1546),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1542),
.B(n_1528),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1538),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1538),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1591),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1590),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1583),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1590),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1596),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1599),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1583),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1593),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1586),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1586),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1597),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1599),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1597),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1571),
.A2(n_1537),
.B1(n_1552),
.B2(n_1522),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1584),
.A2(n_1537),
.B1(n_1529),
.B2(n_1522),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1604),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1603),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1603),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1582),
.A2(n_1529),
.B1(n_1522),
.B2(n_1475),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1598),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1598),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1611),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1610),
.A2(n_1575),
.B(n_1602),
.C(n_1568),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1615),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1611),
.Y(n_1633)
);

AND2x2_ASAP7_75t_SL g1634 ( 
.A(n_1621),
.B(n_1575),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1612),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1615),
.Y(n_1636)
);

AOI332xp33_ASAP7_75t_L g1637 ( 
.A1(n_1629),
.A2(n_1580),
.A3(n_1574),
.B1(n_1557),
.B2(n_1555),
.B3(n_1543),
.C1(n_1541),
.C2(n_1545),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1620),
.A2(n_1569),
.B1(n_1602),
.B2(n_1559),
.C(n_1563),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1628),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1611),
.A2(n_1537),
.B1(n_1529),
.B2(n_1522),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1594),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1607),
.B(n_1593),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1628),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1620),
.A2(n_1529),
.B1(n_1522),
.B2(n_1537),
.Y(n_1644)
);

OAI32xp33_ASAP7_75t_L g1645 ( 
.A1(n_1621),
.A2(n_1585),
.A3(n_1572),
.B1(n_1564),
.B2(n_1578),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1572),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1612),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1646),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1646),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1642),
.B(n_1605),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1633),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1647),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1633),
.B(n_1605),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1630),
.Y(n_1657)
);

AOI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1634),
.A2(n_1625),
.B1(n_1622),
.B2(n_1606),
.C1(n_1623),
.C2(n_1614),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1636),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1635),
.B(n_1614),
.Y(n_1660)
);

OA22x2_ASAP7_75t_L g1661 ( 
.A1(n_1649),
.A2(n_1641),
.B1(n_1648),
.B2(n_1618),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_SL g1662 ( 
.A(n_1658),
.B(n_1637),
.C(n_1631),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1652),
.A2(n_1634),
.B(n_1645),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1650),
.B(n_1638),
.C(n_1639),
.Y(n_1664)
);

NOR3xp33_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1643),
.C(n_1623),
.Y(n_1665)
);

AOI221x1_ASAP7_75t_L g1666 ( 
.A1(n_1657),
.A2(n_1612),
.B1(n_1618),
.B2(n_1629),
.C(n_1617),
.Y(n_1666)
);

NOR4xp25_ASAP7_75t_L g1667 ( 
.A(n_1656),
.B(n_1653),
.C(n_1651),
.D(n_1659),
.Y(n_1667)
);

AOI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1651),
.A2(n_1624),
.B(n_1605),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1652),
.A2(n_1622),
.B(n_1625),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1655),
.A2(n_1644),
.B1(n_1640),
.B2(n_1612),
.C(n_1618),
.Y(n_1670)
);

AOI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1662),
.A2(n_1622),
.B1(n_1625),
.B2(n_1655),
.C(n_1640),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1663),
.A2(n_1619),
.B1(n_1613),
.B2(n_1608),
.C(n_1627),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1661),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1668),
.B(n_1624),
.Y(n_1674)
);

NAND5xp2_ASAP7_75t_L g1675 ( 
.A(n_1669),
.B(n_1660),
.C(n_1624),
.D(n_1578),
.E(n_1616),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_1667),
.B(n_1664),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1675),
.B(n_1674),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1673),
.B(n_1665),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_SL g1679 ( 
.A(n_1672),
.B(n_1608),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1674),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1672),
.B(n_1666),
.C(n_1670),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1678),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1677),
.B(n_1676),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1680),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1681),
.A2(n_1616),
.B(n_1613),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1679),
.A2(n_1619),
.B(n_1617),
.Y(n_1686)
);

NAND5xp2_ASAP7_75t_L g1687 ( 
.A(n_1683),
.B(n_1627),
.C(n_1573),
.D(n_1600),
.E(n_1581),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1684),
.B(n_1618),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1682),
.B(n_1585),
.Y(n_1689)
);

AND3x4_ASAP7_75t_L g1690 ( 
.A(n_1688),
.B(n_1685),
.C(n_1686),
.Y(n_1690)
);

AOI322xp5_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1606),
.A3(n_1687),
.B1(n_1569),
.B2(n_1591),
.C1(n_1601),
.C2(n_1592),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1689),
.C(n_1606),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1691),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1692),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1693),
.A2(n_1589),
.B1(n_1595),
.B2(n_1588),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1694),
.Y(n_1696)
);

XNOR2xp5_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1356),
.Y(n_1697)
);

NAND4xp25_ASAP7_75t_L g1698 ( 
.A(n_1696),
.B(n_1626),
.C(n_1353),
.D(n_1601),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1698),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1697),
.B1(n_1592),
.B2(n_1540),
.Y(n_1700)
);

OA22x2_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1410),
.B1(n_1407),
.B2(n_1587),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1576),
.B1(n_1573),
.B2(n_1626),
.Y(n_1702)
);

AOI211xp5_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1557),
.B(n_1541),
.C(n_1543),
.Y(n_1703)
);


endmodule