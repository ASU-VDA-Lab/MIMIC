module fake_jpeg_15041_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_21),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_48),
.B1(n_19),
.B2(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_52),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_23),
.CON(n_59),
.SN(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_63),
.B1(n_3),
.B2(n_4),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_27),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_77),
.B1(n_64),
.B2(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_95),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_94),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_59),
.A3(n_52),
.B1(n_51),
.B2(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_51),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_53),
.B1(n_49),
.B2(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_64),
.B1(n_80),
.B2(n_82),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_77),
.B1(n_86),
.B2(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_43),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_67),
.B(n_86),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_114),
.B(n_97),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_105),
.B(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_69),
.B1(n_71),
.B2(n_87),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_71),
.B1(n_87),
.B2(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_113),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_80),
.B1(n_92),
.B2(n_84),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_53),
.B1(n_43),
.B2(n_56),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_70),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_70),
.B(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_137),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_95),
.C(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_136),
.C(n_144),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_99),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_107),
.C(n_93),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_155),
.B(n_120),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_122),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_72),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_73),
.C(n_81),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_153),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_114),
.C(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_81),
.Y(n_173)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_92),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_118),
.A2(n_84),
.B1(n_30),
.B2(n_57),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_66),
.B1(n_57),
.B2(n_30),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_163),
.B(n_169),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_155),
.A2(n_131),
.B1(n_115),
.B2(n_126),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_143),
.B1(n_142),
.B2(n_146),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_147),
.A2(n_120),
.B(n_117),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_132),
.B1(n_130),
.B2(n_115),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_173),
.B1(n_177),
.B2(n_149),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_125),
.B(n_83),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_72),
.B1(n_66),
.B2(n_122),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_145),
.B1(n_134),
.B2(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_81),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_23),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_190),
.B1(n_193),
.B2(n_159),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_169),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_135),
.C(n_144),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_186),
.C(n_189),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_137),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_145),
.B1(n_153),
.B2(n_7),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_158),
.C(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_23),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_185),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_157),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_202),
.Y(n_216)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_179),
.B1(n_187),
.B2(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_162),
.C(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_208),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_180),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_217),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_183),
.B1(n_180),
.B2(n_166),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_213),
.A2(n_196),
.B1(n_206),
.B2(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_171),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_207),
.B1(n_195),
.B2(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_200),
.B1(n_201),
.B2(n_205),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_SL g232 ( 
.A(n_222),
.B(n_214),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_233),
.B(n_224),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_226),
.B(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_171),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_234),
.A2(n_211),
.B1(n_171),
.B2(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_16),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_241)
);

AOI321xp33_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_216),
.A3(n_177),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_8),
.B(n_11),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_229),
.Y(n_240)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_241),
.A3(n_243),
.B1(n_235),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_16),
.Y(n_248)
);


endmodule