module fake_jpeg_18845_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2x1_ASAP7_75t_R g45 ( 
.A(n_33),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_26),
.Y(n_54)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_23),
.B1(n_16),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_51),
.B1(n_24),
.B2(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_25),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_38),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_58),
.B1(n_72),
.B2(n_46),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_34),
.B1(n_48),
.B2(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_66),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_36),
.C(n_38),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_58),
.C(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_71),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_35),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_28),
.B(n_19),
.C(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_21),
.Y(n_89)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_29),
.B1(n_19),
.B2(n_28),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_18),
.B(n_20),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_1),
.B(n_2),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_20),
.B(n_31),
.C(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_11),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_92),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_52),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_89),
.B1(n_39),
.B2(n_4),
.Y(n_108)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_65),
.B(n_72),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_64),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_60),
.C(n_61),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_101),
.C(n_103),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_78),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_90),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_75),
.C(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_110),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_30),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_88),
.B(n_89),
.C(n_84),
.D(n_91),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_63),
.C(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_82),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_39),
.C(n_30),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_82),
.B1(n_81),
.B2(n_93),
.C(n_80),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_99),
.B(n_108),
.C(n_8),
.D(n_10),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_130),
.B1(n_4),
.B2(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_104),
.B(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_101),
.C(n_97),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_137),
.C(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_106),
.C(n_114),
.Y(n_137)
);

XOR2x1_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_141),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_134),
.C(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_125),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_149),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_122),
.B1(n_118),
.B2(n_119),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_151),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_124),
.B1(n_123),
.B2(n_116),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_131),
.C(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_158),
.C(n_143),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_151),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_137),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_145),
.C(n_141),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_158),
.C(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_145),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_7),
.B(n_10),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_167),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_161),
.B(n_12),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_167),
.B(n_14),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_14),
.C(n_6),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_170),
.C(n_39),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);


endmodule