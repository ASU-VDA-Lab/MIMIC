module fake_jpeg_24266_n_221 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_221);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_165;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_0),
.B(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_20),
.Y(n_66)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_28),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_28),
.B1(n_31),
.B2(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_33),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_27),
.B(n_26),
.C(n_25),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_22),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_72),
.Y(n_74)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_18),
.B1(n_21),
.B2(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_21),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_79),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_97),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_90),
.Y(n_122)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_38),
.B(n_37),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_51),
.B(n_49),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_95),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_32),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_37),
.C(n_35),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_95),
.C(n_77),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_46),
.B(n_23),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_2),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_63),
.B1(n_52),
.B2(n_68),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_127),
.B1(n_97),
.B2(n_100),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_26),
.B1(n_25),
.B2(n_16),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_68),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_125),
.Y(n_149)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_129),
.B1(n_112),
.B2(n_115),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_51),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_120),
.B(n_85),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_20),
.B1(n_19),
.B2(n_5),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_126),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_19),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_101),
.Y(n_134)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_138),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_140),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_146),
.B1(n_152),
.B2(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_145),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_77),
.B1(n_85),
.B2(n_86),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_73),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_113),
.B(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_93),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_86),
.B1(n_81),
.B2(n_87),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_104),
.C(n_125),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_141),
.C(n_149),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_122),
.C(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_169),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_127),
.B(n_109),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_161),
.B(n_162),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_79),
.B(n_123),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_147),
.B1(n_143),
.B2(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_153),
.B1(n_142),
.B2(n_133),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_173),
.C(n_180),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_146),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_182),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_151),
.C(n_134),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_137),
.C(n_132),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_158),
.B(n_165),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_179),
.B(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_153),
.B1(n_182),
.B2(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_162),
.B(n_133),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_191),
.A2(n_130),
.B(n_176),
.Y(n_195)
);

OAI22x1_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_162),
.B1(n_130),
.B2(n_154),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_192),
.A2(n_144),
.B1(n_168),
.B2(n_159),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_201),
.B1(n_191),
.B2(n_187),
.Y(n_204)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_200),
.B(n_186),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_193),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_172),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_203),
.C(n_189),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_173),
.B(n_140),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_159),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

AOI321xp33_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_208),
.A3(n_144),
.B1(n_15),
.B2(n_7),
.C(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_190),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_209),
.A3(n_203),
.B1(n_15),
.B2(n_10),
.C1(n_13),
.C2(n_103),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_200),
.B(n_202),
.C(n_184),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_4),
.B(n_6),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_213),
.B(n_4),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_211),
.A2(n_207),
.B(n_78),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_78),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_220),
.B(n_7),
.Y(n_221)
);


endmodule