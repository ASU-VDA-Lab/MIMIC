module fake_jpeg_294_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_31),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_44),
.B1(n_36),
.B2(n_41),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_49),
.B1(n_50),
.B2(n_37),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_37),
.C(n_40),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_45),
.C(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_36),
.B1(n_42),
.B2(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_54),
.B1(n_51),
.B2(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_59),
.B(n_47),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_48),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_54),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_50),
.B1(n_34),
.B2(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_57),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_51),
.B(n_55),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_67),
.A3(n_40),
.B1(n_43),
.B2(n_62),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_4),
.C(n_5),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_94),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_2),
.B(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_91),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_73),
.B1(n_82),
.B2(n_77),
.Y(n_99)
);

OR2x6_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_17),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_16),
.B(n_28),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.C(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_7),
.C(n_8),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_86),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_9),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_108),
.C(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_100),
.B(n_101),
.Y(n_112)
);

OA21x2_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_21),
.B(n_24),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_102),
.B1(n_100),
.B2(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_111),
.B1(n_105),
.B2(n_14),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_115),
.A3(n_113),
.B1(n_22),
.B2(n_18),
.C1(n_23),
.C2(n_29),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_14),
.C(n_11),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_13),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_13),
.Y(n_121)
);


endmodule