module fake_netlist_6_987_n_1792 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1792);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1792;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_25),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_89),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_56),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_100),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_0),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_92),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_78),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_69),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_113),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_82),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_29),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_123),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_26),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_66),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_23),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_80),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_138),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_71),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_66),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_23),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_5),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_7),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_96),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_29),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_116),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_61),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_81),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_46),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_154),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_5),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_90),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_95),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_97),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_36),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_102),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_62),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_64),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_115),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_48),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_150),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_3),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_61),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_11),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_104),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_137),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_47),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_105),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_73),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_117),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_0),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_37),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_147),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_128),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_47),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_65),
.Y(n_274)
);

BUFx8_ASAP7_75t_SL g275 ( 
.A(n_140),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_20),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_35),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_38),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_59),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_129),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_70),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_107),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_16),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_124),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_86),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_35),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_153),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_126),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_88),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_136),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_31),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_108),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_83),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_36),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_21),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_42),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_119),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_133),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_64),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_130),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_169),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_40),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_34),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_175),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_37),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_170),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_65),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_146),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_10),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_48),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_155),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_152),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_21),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_79),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_25),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_30),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_14),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_174),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_164),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_4),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_67),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_53),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_120),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_158),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_98),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_22),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_33),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_30),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_27),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_20),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_141),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_94),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_26),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_54),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_17),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_22),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_50),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_109),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_77),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_24),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_93),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_196),
.B(n_1),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_186),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_275),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_225),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_225),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_266),
.B(n_1),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_225),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_289),
.B(n_6),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_236),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_225),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_R g361 ( 
.A(n_266),
.B(n_6),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_225),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_179),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_182),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_197),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_225),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_202),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_227),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_350),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_190),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_201),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_242),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_176),
.B(n_8),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_209),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_201),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_191),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_246),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_246),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_246),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_251),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_266),
.B(n_9),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_246),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_251),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_176),
.B(n_10),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_199),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_204),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_246),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_205),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_246),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_177),
.B(n_183),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_210),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_252),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_252),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_298),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_177),
.B(n_183),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_213),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_299),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_187),
.B(n_11),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_264),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_299),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_189),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_215),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_300),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_224),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_266),
.B(n_12),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_300),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_333),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_216),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_228),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_236),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_234),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_237),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_209),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_247),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_249),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_219),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_219),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_201),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_258),
.Y(n_423)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_178),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_198),
.B(n_12),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_220),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_220),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_181),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_229),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_221),
.B(n_14),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_201),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_281),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_229),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_282),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_356),
.B(n_198),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_381),
.A2(n_323),
.B1(n_255),
.B2(n_212),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_391),
.B(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_226),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_370),
.B(n_287),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g448 ( 
.A1(n_376),
.A2(n_188),
.B(n_187),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_358),
.B(n_184),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_401),
.B(n_184),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_288),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_360),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_360),
.B(n_290),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_362),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_362),
.B(n_291),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_376),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_384),
.A2(n_268),
.B1(n_280),
.B2(n_344),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_366),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_422),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_259),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_422),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_359),
.B(n_224),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_431),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_378),
.B(n_293),
.Y(n_475)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_379),
.A2(n_383),
.B(n_380),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_409),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_388),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_407),
.B(n_226),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_403),
.A2(n_349),
.B1(n_346),
.B2(n_344),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_363),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_359),
.B(n_231),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_231),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_416),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_407),
.B(n_294),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_417),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_393),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_416),
.B(n_296),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_382),
.A2(n_261),
.B(n_256),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_353),
.B(n_184),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_374),
.B(n_297),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_238),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_420),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_393),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_420),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_427),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_425),
.B(n_256),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_375),
.B(n_238),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_385),
.B(n_400),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_429),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_394),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_429),
.B(n_421),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_361),
.A2(n_248),
.B1(n_345),
.B2(n_342),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_364),
.Y(n_513)
);

AND3x1_ASAP7_75t_L g514 ( 
.A(n_450),
.B(n_351),
.C(n_257),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_277),
.B1(n_250),
.B2(n_324),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_459),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_459),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_470),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_469),
.B(n_486),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_435),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_470),
.B(n_369),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_439),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_474),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_449),
.Y(n_526)
);

BUFx4f_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_450),
.A2(n_415),
.B1(n_418),
.B2(n_432),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_469),
.B(n_395),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_442),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_371),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_377),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_480),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_442),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_486),
.B(n_488),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_508),
.A2(n_314),
.B1(n_250),
.B2(n_257),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_386),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_489),
.Y(n_543)
);

BUFx6f_ASAP7_75t_SL g544 ( 
.A(n_505),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_467),
.B(n_512),
.C(n_498),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_444),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_489),
.B(n_387),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_449),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_389),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_449),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_447),
.B(n_392),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_484),
.B(n_430),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_R g558 ( 
.A(n_480),
.B(n_397),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_452),
.B(n_404),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_488),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_498),
.B(n_410),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_454),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_499),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_440),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_505),
.A2(n_306),
.B1(n_260),
.B2(n_346),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_452),
.B(n_412),
.Y(n_570)
);

BUFx16f_ASAP7_75t_R g571 ( 
.A(n_440),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_474),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_499),
.B(n_395),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_482),
.B(n_201),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_495),
.B(n_414),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_462),
.B(n_506),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_457),
.Y(n_578)
);

BUFx4f_ASAP7_75t_L g579 ( 
.A(n_448),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_495),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_463),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_505),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_463),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_465),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_485),
.B(n_419),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_465),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_466),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_456),
.B(n_423),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_506),
.A2(n_430),
.B1(n_434),
.B2(n_262),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_462),
.B(n_352),
.Y(n_592)
);

NOR2x1p5_ASAP7_75t_L g593 ( 
.A(n_511),
.B(n_180),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_477),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_458),
.B(n_269),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_478),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_479),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_460),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_461),
.A2(n_254),
.B1(n_194),
.B2(n_339),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_481),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_438),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_458),
.B(n_283),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_438),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_484),
.B(n_426),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_475),
.B(n_328),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_483),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_461),
.B(n_365),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_483),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_475),
.B(n_367),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_487),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_487),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_476),
.Y(n_618)
);

HB1xp67_ASAP7_75t_SL g619 ( 
.A(n_438),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_460),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_460),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_510),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_446),
.B(n_433),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_446),
.A2(n_331),
.B1(n_277),
.B2(n_279),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_476),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_482),
.B(n_207),
.C(n_203),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_497),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_510),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_510),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_446),
.B(n_408),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_446),
.B(n_305),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_476),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_492),
.B(n_368),
.Y(n_633)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_448),
.A2(n_192),
.B(n_188),
.Y(n_634)
);

AND3x2_ASAP7_75t_L g635 ( 
.A(n_493),
.B(n_292),
.C(n_261),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_493),
.B(n_307),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_448),
.A2(n_279),
.B1(n_343),
.B2(n_331),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_500),
.B(n_201),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_496),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_476),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_500),
.B(n_408),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_476),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_496),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_503),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_490),
.B(n_311),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_460),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_496),
.B(n_306),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_510),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_503),
.B(n_313),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_504),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_504),
.B(n_373),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_460),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_464),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_490),
.B(n_319),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_464),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_507),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_510),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_490),
.B(n_320),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_509),
.B(n_322),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_580),
.B(n_327),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_513),
.B(n_502),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_645),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_526),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_532),
.B(n_502),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_645),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_580),
.B(n_502),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_651),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_609),
.A2(n_437),
.B(n_436),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_564),
.B(n_502),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_607),
.B(n_230),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_651),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_517),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_655),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_607),
.B(n_230),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_545),
.B(n_211),
.C(n_208),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_618),
.A2(n_509),
.B(n_312),
.C(n_315),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_517),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_655),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_521),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_521),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_514),
.B(n_301),
.C(n_267),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_490),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_658),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_526),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_525),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_535),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_519),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_607),
.Y(n_691)
);

INVx8_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_582),
.B(n_230),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_530),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_632),
.A2(n_312),
.B1(n_315),
.B2(n_321),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_572),
.B(n_184),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_575),
.B(n_510),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_530),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_595),
.B(n_218),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_572),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_597),
.B(n_192),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_598),
.B(n_295),
.C(n_244),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_608),
.B(n_222),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_597),
.B(n_193),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_615),
.A2(n_332),
.B1(n_348),
.B2(n_347),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_582),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_577),
.B(n_232),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_611),
.B(n_235),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_582),
.B(n_527),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_619),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_625),
.A2(n_321),
.B(n_324),
.C(n_329),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_543),
.B(n_193),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_541),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_525),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_551),
.B(n_195),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_541),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_632),
.A2(n_329),
.B1(n_343),
.B2(n_200),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_641),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_556),
.B(n_195),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_640),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_559),
.B(n_200),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_560),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_577),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_641),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_527),
.A2(n_436),
.B(n_473),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_560),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_SL g727 ( 
.A(n_627),
.B(n_239),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_527),
.B(n_230),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_549),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_640),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_570),
.B(n_253),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_549),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_633),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_625),
.A2(n_241),
.B1(n_214),
.B2(n_217),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_520),
.B(n_310),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_573),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_563),
.B(n_230),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_563),
.B(n_230),
.Y(n_738)
);

NOR3xp33_ASAP7_75t_SL g739 ( 
.A(n_604),
.B(n_271),
.C(n_272),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_520),
.B(n_310),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_630),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_533),
.B(n_542),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_562),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_515),
.B(n_273),
.C(n_274),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_537),
.B(n_206),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_642),
.A2(n_233),
.B1(n_214),
.B2(n_217),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_566),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_630),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_537),
.B(n_548),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_562),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_579),
.B(n_316),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_578),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_548),
.B(n_206),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_522),
.B(n_223),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_524),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_610),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_578),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_579),
.B(n_642),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_553),
.B(n_223),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_524),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_579),
.B(n_316),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_637),
.B(n_334),
.Y(n_762)
);

CKINVDCx16_ASAP7_75t_R g763 ( 
.A(n_558),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_529),
.B(n_233),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_592),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_529),
.B(n_240),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_531),
.B(n_240),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_544),
.A2(n_340),
.B1(n_341),
.B2(n_241),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_531),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_536),
.B(n_243),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_536),
.B(n_243),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_539),
.B(n_245),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_539),
.B(n_546),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_581),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_546),
.B(n_245),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_555),
.B(n_263),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_573),
.B(n_310),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_555),
.B(n_263),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_623),
.B(n_276),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_623),
.B(n_265),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_639),
.A2(n_265),
.B(n_270),
.C(n_303),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_639),
.B(n_270),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_565),
.B(n_303),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_583),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_523),
.B(n_278),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_565),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_643),
.B(n_308),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_523),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_576),
.B(n_308),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_583),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_540),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_643),
.B(n_330),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_576),
.Y(n_794)
);

BUFx5_ASAP7_75t_L g795 ( 
.A(n_638),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_591),
.B(n_547),
.Y(n_796)
);

INVxp33_ASAP7_75t_L g797 ( 
.A(n_633),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_584),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_584),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_586),
.B(n_330),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_586),
.B(n_445),
.Y(n_801)
);

BUFx8_ASAP7_75t_L g802 ( 
.A(n_544),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_652),
.B(n_310),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_594),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_587),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_594),
.B(n_464),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_627),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_587),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_613),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_585),
.B(n_631),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_588),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_593),
.B(n_284),
.Y(n_812)
);

NAND2x1_ASAP7_75t_L g813 ( 
.A(n_516),
.B(n_445),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_557),
.A2(n_285),
.B1(n_286),
.B2(n_302),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_636),
.B(n_304),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_557),
.B(n_309),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_622),
.B(n_464),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_534),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_L g819 ( 
.A1(n_538),
.A2(n_317),
.B1(n_318),
.B2(n_325),
.C(n_326),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_557),
.B(n_335),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_534),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_596),
.B(n_464),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_557),
.B(n_336),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_650),
.B(n_338),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_588),
.B(n_445),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_589),
.B(n_600),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_540),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_596),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_589),
.B(n_445),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_600),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_691),
.A2(n_646),
.B(n_660),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_809),
.B(n_571),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_691),
.A2(n_656),
.B(n_647),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_742),
.B(n_602),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_720),
.B(n_730),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_723),
.B(n_610),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_674),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_690),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_810),
.B(n_602),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_700),
.Y(n_840)
);

AOI21xp33_ASAP7_75t_L g841 ( 
.A1(n_699),
.A2(n_610),
.B(n_626),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_697),
.A2(n_561),
.B(n_550),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_728),
.A2(n_648),
.B(n_634),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_720),
.B(n_622),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_688),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_821),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_796),
.A2(n_569),
.B(n_624),
.C(n_614),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_810),
.B(n_749),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_751),
.A2(n_761),
.B(n_737),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_728),
.A2(n_738),
.B(n_737),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_803),
.B(n_610),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_731),
.B(n_606),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_738),
.A2(n_648),
.B(n_634),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_731),
.B(n_606),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_679),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_796),
.A2(n_614),
.B(n_617),
.C(n_616),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_699),
.B(n_599),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_761),
.A2(n_561),
.B(n_550),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_720),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_758),
.A2(n_648),
.B(n_659),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_758),
.A2(n_620),
.B(n_550),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_714),
.B(n_661),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_789),
.B(n_703),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_730),
.B(n_605),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_692),
.B(n_648),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_778),
.B(n_568),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_671),
.A2(n_554),
.B(n_657),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_783),
.A2(n_574),
.B(n_612),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_703),
.B(n_612),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_L g870 ( 
.A(n_730),
.B(n_616),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_708),
.B(n_617),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_708),
.B(n_516),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_783),
.A2(n_628),
.B(n_629),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_672),
.A2(n_659),
.B(n_629),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_730),
.B(n_628),
.Y(n_875)
);

AOI22x1_ASAP7_75t_L g876 ( 
.A1(n_664),
.A2(n_644),
.B1(n_649),
.B2(n_653),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_788),
.A2(n_644),
.B(n_649),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_663),
.A2(n_568),
.B1(n_516),
.B2(n_653),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_788),
.A2(n_518),
.B(n_552),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_766),
.B(n_337),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_666),
.B(n_715),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_736),
.B(n_518),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_684),
.B(n_518),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_709),
.A2(n_725),
.B(n_668),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_696),
.B(n_398),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_719),
.A2(n_574),
.B1(n_567),
.B2(n_653),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_709),
.A2(n_657),
.B(n_654),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_721),
.B(n_552),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_667),
.B(n_552),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_792),
.A2(n_657),
.B(n_654),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_792),
.A2(n_657),
.B(n_654),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_745),
.A2(n_621),
.B1(n_567),
.B2(n_601),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_793),
.A2(n_621),
.B(n_567),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_792),
.A2(n_657),
.B(n_654),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_792),
.A2(n_654),
.B(n_647),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_763),
.B(n_398),
.C(n_399),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_678),
.A2(n_501),
.B(n_494),
.C(n_405),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_669),
.B(n_673),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_827),
.A2(n_826),
.B(n_774),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_706),
.B(n_722),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_675),
.B(n_601),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_827),
.A2(n_647),
.B(n_550),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_827),
.A2(n_647),
.B(n_550),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_734),
.A2(n_399),
.B(n_402),
.C(n_405),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_793),
.A2(n_621),
.B(n_601),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_717),
.A2(n_473),
.B(n_436),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_717),
.A2(n_676),
.B(n_693),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_827),
.A2(n_647),
.B(n_554),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_681),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_711),
.A2(n_501),
.B(n_494),
.C(n_402),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_680),
.B(n_554),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_682),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_676),
.A2(n_822),
.B(n_806),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_693),
.A2(n_620),
.B(n_603),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_685),
.B(n_554),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_686),
.B(n_554),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_734),
.A2(n_638),
.B1(n_494),
.B2(n_501),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_677),
.B(n_85),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_801),
.A2(n_620),
.B(n_603),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_735),
.B(n_635),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_701),
.A2(n_437),
.B(n_468),
.C(n_473),
.Y(n_922)
);

NOR2x1_ASAP7_75t_R g923 ( 
.A(n_807),
.B(n_464),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_825),
.A2(n_620),
.B(n_603),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_829),
.A2(n_620),
.B(n_603),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_755),
.B(n_603),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_706),
.A2(n_455),
.B(n_472),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_687),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_704),
.A2(n_455),
.B(n_472),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_687),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_746),
.A2(n_468),
.B1(n_437),
.B2(n_455),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_762),
.A2(n_455),
.B(n_472),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_760),
.B(n_770),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_689),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_787),
.B(n_638),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_806),
.A2(n_472),
.B(n_471),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_722),
.B(n_472),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_689),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_687),
.B(n_472),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_822),
.A2(n_472),
.B(n_471),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_794),
.B(n_638),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_687),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_741),
.A2(n_638),
.B1(n_471),
.B2(n_464),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_798),
.B(n_638),
.Y(n_944)
);

CKINVDCx8_ASAP7_75t_R g945 ( 
.A(n_692),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_726),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_799),
.B(n_468),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_805),
.B(n_471),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_781),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_713),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_718),
.B(n_471),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_740),
.B(n_18),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_748),
.A2(n_471),
.B1(n_173),
.B2(n_172),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_813),
.A2(n_471),
.B(n_171),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_662),
.A2(n_166),
.B(n_165),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_746),
.A2(n_160),
.B(n_156),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_695),
.A2(n_19),
.B(n_24),
.C(n_27),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_713),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_716),
.A2(n_148),
.B(n_144),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_716),
.A2(n_135),
.B(n_134),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_808),
.B(n_811),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_665),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_830),
.B(n_19),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_729),
.A2(n_131),
.B(n_127),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_732),
.A2(n_750),
.B(n_804),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_786),
.B(n_28),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_695),
.B(n_111),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_782),
.A2(n_712),
.B(n_698),
.C(n_694),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_732),
.A2(n_106),
.B(n_84),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_710),
.B(n_28),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_707),
.B(n_31),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_743),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_665),
.Y(n_973)
);

AOI21xp33_ASAP7_75t_L g974 ( 
.A1(n_815),
.A2(n_824),
.B(n_780),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_SL g975 ( 
.A(n_818),
.B(n_32),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_724),
.B(n_34),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_743),
.A2(n_39),
.B(n_40),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_780),
.B(n_39),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_750),
.B(n_41),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_812),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_670),
.A2(n_41),
.B(n_43),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_759),
.B(n_43),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_752),
.A2(n_828),
.B(n_804),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_752),
.B(n_44),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_757),
.B(n_44),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_757),
.B(n_828),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_765),
.A2(n_46),
.B(n_49),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_765),
.A2(n_775),
.B(n_791),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_775),
.A2(n_49),
.B(n_50),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_L g990 ( 
.A(n_795),
.B(n_51),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_785),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_785),
.B(n_51),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_764),
.A2(n_771),
.B(n_767),
.C(n_800),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_791),
.B(n_52),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_817),
.Y(n_995)
);

AND2x2_ASAP7_75t_SL g996 ( 
.A(n_815),
.B(n_52),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_753),
.B(n_53),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_768),
.B(n_55),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_754),
.A2(n_55),
.B(n_57),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_772),
.A2(n_57),
.B(n_58),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_773),
.B(n_58),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_816),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_776),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_777),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_779),
.B(n_60),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_784),
.A2(n_63),
.B(n_790),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_817),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_818),
.B(n_63),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_795),
.B(n_739),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_824),
.A2(n_702),
.B(n_692),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_945),
.Y(n_1011)
);

OAI21xp33_ASAP7_75t_SL g1012 ( 
.A1(n_956),
.A2(n_823),
.B(n_820),
.Y(n_1012)
);

NAND2xp33_ASAP7_75t_SL g1013 ( 
.A(n_851),
.B(n_756),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_844),
.Y(n_1014)
);

O2A1O1Ixp5_ASAP7_75t_L g1015 ( 
.A1(n_974),
.A2(n_727),
.B(n_683),
.C(n_814),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_846),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_996),
.A2(n_756),
.B1(n_769),
.B2(n_744),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_845),
.B(n_802),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_841),
.A2(n_705),
.B(n_819),
.C(n_733),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_928),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_928),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_917),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_848),
.B(n_817),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_840),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_849),
.A2(n_795),
.B(n_817),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_L g1026 ( 
.A(n_962),
.B(n_747),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_863),
.B(n_797),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_838),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_839),
.B(n_834),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_978),
.A2(n_795),
.B(n_817),
.C(n_850),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_852),
.B(n_795),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_854),
.B(n_795),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_844),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_863),
.B(n_881),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_832),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_966),
.A2(n_957),
.B(n_963),
.C(n_970),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1004),
.B(n_885),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_832),
.B(n_996),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_866),
.B(n_857),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_928),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_831),
.A2(n_884),
.B(n_833),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_837),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_880),
.B(n_1002),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_899),
.A2(n_870),
.B(n_853),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_966),
.A2(n_967),
.B1(n_952),
.B2(n_1003),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_869),
.B(n_871),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_898),
.B(n_933),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_961),
.B(n_847),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_1010),
.B(n_862),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_843),
.A2(n_872),
.B(n_842),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_836),
.B(n_980),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1002),
.B(n_896),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_855),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_835),
.A2(n_867),
.B(n_907),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_835),
.A2(n_888),
.B(n_860),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_836),
.A2(n_921),
.B1(n_878),
.B2(n_970),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_847),
.B(n_972),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_982),
.B(n_917),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_856),
.A2(n_965),
.B(n_988),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_972),
.B(n_856),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_968),
.A2(n_993),
.B(n_981),
.C(n_976),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_882),
.B(n_946),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_946),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_882),
.B(n_997),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_971),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_928),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_991),
.B(n_938),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_930),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_R g1069 ( 
.A(n_962),
.B(n_930),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_973),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_883),
.A2(n_864),
.B(n_875),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_957),
.A2(n_904),
.B1(n_918),
.B2(n_953),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1008),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_949),
.A2(n_990),
.B(n_1006),
.C(n_998),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1001),
.B(n_1005),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_SL g1076 ( 
.A1(n_1009),
.A2(n_979),
.B(n_994),
.C(n_904),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_865),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_975),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_942),
.B(n_859),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_865),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_979),
.A2(n_994),
.B(n_985),
.C(n_992),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_909),
.B(n_912),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_883),
.A2(n_864),
.B(n_875),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_900),
.B(n_942),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_934),
.B(n_950),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_986),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_868),
.A2(n_887),
.B(n_1009),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_918),
.A2(n_865),
.B1(n_995),
.B2(n_886),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_919),
.A2(n_983),
.B(n_999),
.C(n_1000),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_995),
.A2(n_984),
.B1(n_916),
.B2(n_926),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_844),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_900),
.B(n_915),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_1007),
.A2(n_877),
.B(n_873),
.C(n_955),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_939),
.Y(n_1094)
);

INVxp33_ASAP7_75t_SL g1095 ( 
.A(n_923),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_911),
.B(n_901),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_977),
.B(n_989),
.C(n_987),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_951),
.A2(n_897),
.B(n_889),
.C(n_910),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_951),
.A2(n_937),
.B1(n_935),
.B2(n_941),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_844),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_844),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_939),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_944),
.B(n_948),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_947),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_937),
.B(n_892),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_858),
.A2(n_861),
.B(n_908),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_906),
.A2(n_943),
.B1(n_905),
.B2(n_879),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_890),
.A2(n_903),
.B(n_902),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_922),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_891),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_931),
.Y(n_1111)
);

OA22x2_ASAP7_75t_L g1112 ( 
.A1(n_893),
.A2(n_913),
.B1(n_876),
.B2(n_874),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_929),
.B(n_924),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_914),
.A2(n_925),
.B(n_920),
.C(n_932),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_927),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_959),
.A2(n_969),
.B(n_964),
.C(n_960),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_SL g1117 ( 
.A1(n_954),
.A2(n_894),
.B1(n_895),
.B2(n_936),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_L g1118 ( 
.A1(n_940),
.A2(n_974),
.B(n_978),
.C(n_841),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_837),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_849),
.A2(n_691),
.B(n_563),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_974),
.A2(n_978),
.B(n_841),
.C(n_513),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_849),
.A2(n_691),
.B(n_563),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_974),
.A2(n_841),
.B(n_796),
.C(n_545),
.Y(n_1123)
);

BUFx8_ASAP7_75t_L g1124 ( 
.A(n_845),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_849),
.A2(n_691),
.B(n_563),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_958),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_837),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_974),
.A2(n_841),
.B(n_796),
.C(n_545),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_849),
.A2(n_691),
.B(n_563),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_974),
.A2(n_810),
.B(n_513),
.C(n_532),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_845),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_848),
.B(n_834),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_848),
.B(n_834),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_974),
.A2(n_978),
.B(n_841),
.C(n_513),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_865),
.B(n_692),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_849),
.A2(n_691),
.B(n_563),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_928),
.Y(n_1137)
);

BUFx5_ASAP7_75t_L g1138 ( 
.A(n_844),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_974),
.B(n_863),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_958),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_928),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_974),
.A2(n_841),
.B(n_796),
.C(n_545),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_974),
.B(n_513),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_848),
.B(n_834),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_838),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_974),
.A2(n_978),
.B(n_841),
.C(n_513),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_958),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_996),
.A2(n_746),
.B1(n_734),
.B2(n_717),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_SL g1149 ( 
.A1(n_974),
.A2(n_508),
.B(n_981),
.C(n_841),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_958),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_974),
.A2(n_841),
.B(n_796),
.C(n_545),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_849),
.A2(n_691),
.B(n_563),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_SL g1153 ( 
.A(n_945),
.B(n_720),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_848),
.B(n_839),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1131),
.Y(n_1155)
);

BUFx8_ASAP7_75t_L g1156 ( 
.A(n_1028),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1044),
.A2(n_1050),
.B(n_1041),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1143),
.A2(n_1027),
.B1(n_1035),
.B2(n_1038),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1123),
.B(n_1142),
.C(n_1128),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1061),
.A2(n_1046),
.B(n_1029),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1042),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1120),
.A2(n_1125),
.B(n_1122),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1030),
.A2(n_1151),
.A3(n_1089),
.B(n_1090),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1053),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1130),
.A2(n_1121),
.B(n_1146),
.C(n_1134),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1139),
.A2(n_1019),
.B(n_1036),
.C(n_1039),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1129),
.A2(n_1152),
.B(n_1136),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1091),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1144),
.B(n_1154),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1144),
.A2(n_1047),
.B(n_1054),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1059),
.A2(n_1097),
.B(n_1114),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1037),
.B(n_1048),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1014),
.A2(n_1033),
.B(n_1049),
.Y(n_1175)
);

AOI221xp5_ASAP7_75t_L g1176 ( 
.A1(n_1148),
.A2(n_1017),
.B1(n_1012),
.B2(n_1065),
.C(n_1078),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1149),
.A2(n_1118),
.B(n_1055),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1014),
.A2(n_1033),
.B(n_1059),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1043),
.B(n_1073),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1014),
.A2(n_1033),
.B(n_1113),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1135),
.B(n_1024),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1015),
.A2(n_1148),
.B(n_1045),
.C(n_1056),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1074),
.A2(n_1081),
.B(n_1075),
.C(n_1058),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1022),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1017),
.A2(n_1051),
.B(n_1064),
.C(n_1052),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1124),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1014),
.A2(n_1033),
.B(n_1032),
.Y(n_1187)
);

BUFx10_ASAP7_75t_L g1188 ( 
.A(n_1016),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1057),
.A2(n_1023),
.B(n_1072),
.C(n_1093),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1063),
.B(n_1145),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1072),
.A2(n_1057),
.B1(n_1101),
.B2(n_1094),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1091),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1090),
.A2(n_1107),
.A3(n_1116),
.B(n_1088),
.Y(n_1193)
);

AOI221x1_ASAP7_75t_L g1194 ( 
.A1(n_1108),
.A2(n_1109),
.B1(n_1083),
.B2(n_1071),
.C(n_1013),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1031),
.A2(n_1096),
.B(n_1025),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1060),
.A2(n_1062),
.B1(n_1119),
.B2(n_1127),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1115),
.A2(n_1103),
.B(n_1092),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1086),
.A2(n_1111),
.B1(n_1091),
.B2(n_1100),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1085),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1124),
.Y(n_1200)
);

AND2x6_ASAP7_75t_L g1201 ( 
.A(n_1021),
.B(n_1141),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1076),
.A2(n_1112),
.B(n_1098),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1070),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1110),
.A2(n_1084),
.A3(n_1104),
.B(n_1067),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1105),
.A2(n_1099),
.B(n_1102),
.C(n_1153),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1077),
.A2(n_1080),
.B1(n_1018),
.B2(n_1095),
.C(n_1082),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1117),
.A2(n_1087),
.B(n_1110),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1150),
.B(n_1147),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1135),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1040),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1069),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1087),
.A2(n_1138),
.B(n_1140),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1126),
.A2(n_1026),
.B(n_1020),
.C(n_1137),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1040),
.A2(n_1068),
.A3(n_1138),
.B(n_1079),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1021),
.B(n_1066),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1011),
.B(n_1021),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1138),
.A2(n_1068),
.B(n_1066),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1138),
.A2(n_1066),
.B(n_1141),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1138),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1138),
.A2(n_691),
.B(n_1044),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1044),
.A2(n_1054),
.B(n_1050),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1034),
.B(n_1132),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1061),
.A2(n_856),
.A3(n_1030),
.B(n_1123),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1143),
.B(n_974),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1148),
.A2(n_956),
.B(n_1061),
.Y(n_1227)
);

CKINVDCx16_ASAP7_75t_R g1228 ( 
.A(n_1018),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1061),
.A2(n_1041),
.B(n_974),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1143),
.A2(n_1027),
.B1(n_974),
.B2(n_807),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_1143),
.A2(n_1134),
.B(n_1121),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1011),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1061),
.A2(n_1059),
.B(n_1054),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1148),
.A2(n_1143),
.B1(n_1132),
.B2(n_1133),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_1024),
.B(n_690),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1061),
.A2(n_1041),
.B(n_974),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_SL g1242 ( 
.A1(n_1057),
.A2(n_956),
.B(n_981),
.Y(n_1242)
);

AOI31xp67_ASAP7_75t_L g1243 ( 
.A1(n_1112),
.A2(n_1049),
.A3(n_1113),
.B(n_1139),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1143),
.B(n_974),
.C(n_1123),
.Y(n_1244)
);

AOI31xp67_ASAP7_75t_L g1245 ( 
.A1(n_1112),
.A2(n_1049),
.A3(n_1113),
.B(n_1139),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1143),
.A2(n_974),
.B(n_1134),
.C(n_1121),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1061),
.A2(n_1059),
.B(n_1054),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1249)
);

NOR4xp25_ASAP7_75t_L g1250 ( 
.A(n_1123),
.B(n_1142),
.C(n_1151),
.D(n_1128),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1061),
.A2(n_856),
.A3(n_1030),
.B(n_1123),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1143),
.B(n_974),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1043),
.B(n_866),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1143),
.A2(n_974),
.B(n_1134),
.C(n_1121),
.Y(n_1254)
);

OAI22x1_ASAP7_75t_L g1255 ( 
.A1(n_1143),
.A2(n_1038),
.B1(n_1056),
.B2(n_966),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1148),
.A2(n_1143),
.B1(n_1132),
.B2(n_1133),
.Y(n_1256)
);

AOI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1143),
.A2(n_1134),
.B(n_1121),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1043),
.B(n_866),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1143),
.A2(n_974),
.B(n_1134),
.C(n_1121),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1143),
.A2(n_1130),
.B(n_974),
.C(n_1128),
.Y(n_1260)
);

CKINVDCx8_ASAP7_75t_R g1261 ( 
.A(n_1016),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1128),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1021),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1143),
.A2(n_974),
.B(n_1134),
.C(n_1121),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1061),
.A2(n_1059),
.B(n_1054),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1091),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1143),
.B(n_974),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1091),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1022),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1128),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1128),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1149),
.A2(n_1143),
.B(n_1128),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1043),
.B(n_866),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1282)
);

AOI31xp67_ASAP7_75t_L g1283 ( 
.A1(n_1112),
.A2(n_1049),
.A3(n_1113),
.B(n_1139),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1044),
.A2(n_691),
.B(n_1050),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1041),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1143),
.A2(n_1027),
.B1(n_974),
.B2(n_807),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1034),
.B(n_1132),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1131),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1143),
.A2(n_974),
.B(n_532),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1016),
.Y(n_1292)
);

OAI22x1_ASAP7_75t_L g1293 ( 
.A1(n_1226),
.A2(n_1271),
.B1(n_1252),
.B2(n_1244),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1235),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1244),
.A2(n_1160),
.B1(n_1256),
.B2(n_1238),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1291),
.A2(n_1230),
.B1(n_1288),
.B2(n_1159),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1272),
.B(n_1211),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1163),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1166),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1224),
.B(n_1289),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1156),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1156),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1255),
.A2(n_1231),
.B1(n_1160),
.B2(n_1257),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1257),
.A2(n_1238),
.B1(n_1256),
.B2(n_1176),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1171),
.A2(n_1234),
.B1(n_1157),
.B2(n_1249),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1216),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1161),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1171),
.A2(n_1233),
.B1(n_1157),
.B2(n_1280),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1292),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1291),
.A2(n_1281),
.B1(n_1258),
.B2(n_1253),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1261),
.Y(n_1311)
);

BUFx8_ASAP7_75t_SL g1312 ( 
.A(n_1200),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1181),
.Y(n_1313)
);

INVx5_ASAP7_75t_L g1314 ( 
.A(n_1201),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1264),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1162),
.A2(n_1232),
.B1(n_1280),
.B2(n_1234),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1162),
.B(n_1232),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1233),
.A2(n_1249),
.B1(n_1266),
.B2(n_1227),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1266),
.A2(n_1265),
.B1(n_1254),
.B2(n_1259),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1188),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1174),
.B(n_1179),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1239),
.A2(n_1206),
.B1(n_1247),
.B2(n_1191),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1272),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1182),
.A2(n_1174),
.B1(n_1191),
.B2(n_1185),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1262),
.A2(n_1279),
.B1(n_1278),
.B2(n_1277),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1188),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1208),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1242),
.A2(n_1262),
.B1(n_1279),
.B2(n_1278),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1277),
.A2(n_1229),
.B1(n_1240),
.B2(n_1268),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1199),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1229),
.A2(n_1240),
.B1(n_1248),
.B2(n_1268),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1184),
.B(n_1250),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_R g1334 ( 
.A1(n_1186),
.A2(n_1203),
.B1(n_1275),
.B2(n_1290),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1196),
.Y(n_1335)
);

BUFx8_ASAP7_75t_L g1336 ( 
.A(n_1155),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1215),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1168),
.B(n_1172),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1215),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1209),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1228),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1264),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1205),
.A2(n_1183),
.B1(n_1198),
.B2(n_1197),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1260),
.B(n_1167),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1170),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1213),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1192),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1237),
.A2(n_1248),
.B1(n_1202),
.B2(n_1173),
.Y(n_1348)
);

CKINVDCx11_ASAP7_75t_R g1349 ( 
.A(n_1219),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1237),
.A2(n_1173),
.B1(n_1177),
.B2(n_1198),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1204),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1204),
.Y(n_1352)
);

NAND2xp33_ASAP7_75t_SL g1353 ( 
.A(n_1192),
.B(n_1270),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1178),
.A2(n_1194),
.B1(n_1177),
.B2(n_1220),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1201),
.Y(n_1355)
);

BUFx8_ASAP7_75t_L g1356 ( 
.A(n_1201),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1270),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1214),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1210),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1210),
.A2(n_1243),
.B1(n_1283),
.B2(n_1245),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1207),
.A2(n_1195),
.B1(n_1158),
.B2(n_1285),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1175),
.A2(n_1180),
.B1(n_1187),
.B2(n_1212),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1222),
.A2(n_1284),
.B1(n_1282),
.B2(n_1269),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1217),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1236),
.A2(n_1263),
.B1(n_1164),
.B2(n_1169),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1218),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1193),
.A2(n_1165),
.B1(n_1251),
.B2(n_1225),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1221),
.A2(n_1246),
.B(n_1286),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1189),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1223),
.A2(n_1287),
.B1(n_1273),
.B2(n_1276),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_1241),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1267),
.A2(n_1274),
.B1(n_1193),
.B2(n_1251),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1193),
.A2(n_996),
.B1(n_1148),
.B2(n_1143),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1171),
.A2(n_1143),
.B1(n_1162),
.B2(n_1157),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1291),
.A2(n_1143),
.B(n_528),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1264),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1190),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1190),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1226),
.A2(n_996),
.B1(n_1148),
.B2(n_1143),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1226),
.A2(n_1148),
.B1(n_975),
.B2(n_1252),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1156),
.Y(n_1381)
);

CKINVDCx11_ASAP7_75t_R g1382 ( 
.A(n_1261),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1156),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1261),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1226),
.A2(n_1252),
.B1(n_1271),
.B2(n_1143),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1226),
.A2(n_1252),
.B1(n_1271),
.B2(n_1143),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1226),
.A2(n_996),
.B1(n_1148),
.B2(n_1143),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1156),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1264),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1264),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1171),
.A2(n_1143),
.B1(n_1162),
.B2(n_1157),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1261),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1226),
.A2(n_996),
.B1(n_1148),
.B2(n_1143),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1235),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1226),
.A2(n_1252),
.B1(n_1271),
.B2(n_1143),
.Y(n_1395)
);

BUFx2_ASAP7_75t_R g1396 ( 
.A(n_1261),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1373),
.B(n_1328),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1365),
.A2(n_1361),
.B(n_1363),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1307),
.A2(n_1338),
.B(n_1361),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1333),
.B(n_1332),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1298),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1354),
.A2(n_1368),
.B(n_1352),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1378),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1344),
.A2(n_1362),
.B(n_1343),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1337),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1351),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1339),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1328),
.B(n_1335),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1366),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1377),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1295),
.B(n_1367),
.Y(n_1411)
);

OAI21xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1307),
.A2(n_1304),
.B(n_1317),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1363),
.A2(n_1370),
.B(n_1331),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1330),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1293),
.A2(n_1319),
.B(n_1324),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1367),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1364),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1374),
.B(n_1391),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1299),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1371),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1325),
.A2(n_1329),
.B(n_1331),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1318),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1314),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1370),
.A2(n_1372),
.B(n_1329),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1358),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1372),
.A2(n_1350),
.B(n_1325),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1360),
.B(n_1297),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1348),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1316),
.B(n_1305),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1308),
.B(n_1385),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1295),
.B(n_1303),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1354),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1346),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1303),
.B(n_1379),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1358),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1350),
.A2(n_1304),
.B(n_1375),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1321),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1327),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1379),
.A2(n_1387),
.B1(n_1393),
.B2(n_1395),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_L g1441 ( 
.A(n_1386),
.B(n_1395),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1297),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1387),
.A2(n_1393),
.B(n_1380),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1380),
.A2(n_1296),
.B(n_1322),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1296),
.A2(n_1310),
.B1(n_1334),
.B2(n_1300),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1364),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1369),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1369),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1314),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1356),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1349),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1353),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1356),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1323),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1306),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1349),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1313),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1357),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1355),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1345),
.A2(n_1320),
.B(n_1381),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1294),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1355),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1359),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1315),
.B(n_1376),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1315),
.B(n_1376),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1383),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1342),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1342),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1443),
.A2(n_1340),
.B(n_1302),
.C(n_1301),
.Y(n_1469)
);

OAI211xp5_ASAP7_75t_L g1470 ( 
.A1(n_1443),
.A2(n_1326),
.B(n_1311),
.C(n_1392),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1440),
.A2(n_1431),
.B1(n_1445),
.B2(n_1411),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1424),
.A2(n_1347),
.B(n_1390),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_SL g1473 ( 
.A(n_1440),
.B(n_1396),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1429),
.B(n_1390),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1433),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1419),
.Y(n_1476)
);

NAND2x1_ASAP7_75t_L g1477 ( 
.A(n_1460),
.B(n_1388),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1415),
.A2(n_1341),
.B(n_1326),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1400),
.B(n_1389),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1441),
.A2(n_1376),
.B1(n_1311),
.B2(n_1392),
.C(n_1382),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1429),
.B(n_1336),
.Y(n_1481)
);

AOI211xp5_ASAP7_75t_L g1482 ( 
.A1(n_1439),
.A2(n_1382),
.B(n_1384),
.C(n_1309),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1400),
.B(n_1384),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1439),
.A2(n_1430),
.B(n_1418),
.C(n_1444),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1467),
.Y(n_1485)
);

INVx5_ASAP7_75t_SL g1486 ( 
.A(n_1451),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_SL g1487 ( 
.A1(n_1430),
.A2(n_1394),
.B(n_1309),
.C(n_1336),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1418),
.B(n_1437),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1403),
.B(n_1312),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1399),
.B(n_1427),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1404),
.A2(n_1412),
.B(n_1445),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1450),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1408),
.B(n_1455),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1444),
.A2(n_1431),
.B(n_1412),
.C(n_1434),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1413),
.A2(n_1424),
.B(n_1402),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1434),
.A2(n_1444),
.B1(n_1397),
.B2(n_1432),
.C(n_1411),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1424),
.A2(n_1426),
.B(n_1413),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1405),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1410),
.B(n_1417),
.Y(n_1499)
);

NAND2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1460),
.B(n_1442),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1397),
.A2(n_1447),
.B1(n_1448),
.B2(n_1436),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1425),
.B(n_1435),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1460),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1417),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1422),
.A2(n_1398),
.B(n_1436),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1422),
.B(n_1401),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1417),
.B(n_1446),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_SL g1508 ( 
.A1(n_1462),
.A2(n_1452),
.B(n_1423),
.C(n_1449),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1425),
.B(n_1435),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1444),
.A2(n_1446),
.B1(n_1436),
.B2(n_1448),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_SL g1511 ( 
.A(n_1461),
.B(n_1462),
.C(n_1454),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1467),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1436),
.A2(n_1446),
.B1(n_1425),
.B2(n_1435),
.Y(n_1513)
);

AO32x2_ASAP7_75t_L g1514 ( 
.A1(n_1409),
.A2(n_1420),
.A3(n_1457),
.B1(n_1423),
.B2(n_1459),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1407),
.B(n_1464),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1460),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1447),
.A2(n_1448),
.B1(n_1461),
.B2(n_1453),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_SL g1519 ( 
.A1(n_1452),
.A2(n_1423),
.B(n_1449),
.C(n_1463),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_SL g1520 ( 
.A(n_1466),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1447),
.A2(n_1448),
.B1(n_1456),
.B2(n_1451),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1467),
.Y(n_1522)
);

OAI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1458),
.A2(n_1447),
.B1(n_1448),
.B2(n_1451),
.C(n_1456),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1451),
.B(n_1456),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1438),
.B(n_1414),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1468),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1468),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1514),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1476),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1517),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1497),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1522),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1503),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1495),
.B(n_1402),
.Y(n_1535)
);

NOR2xp67_ASAP7_75t_L g1536 ( 
.A(n_1501),
.B(n_1420),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1475),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1498),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1488),
.B(n_1416),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1505),
.B(n_1402),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1505),
.B(n_1472),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1477),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1526),
.Y(n_1543)
);

AND2x2_ASAP7_75t_SL g1544 ( 
.A(n_1496),
.B(n_1421),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1472),
.B(n_1402),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1514),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1514),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1490),
.B(n_1426),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1506),
.Y(n_1550)
);

NOR2x1_ASAP7_75t_L g1551 ( 
.A(n_1523),
.B(n_1501),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1490),
.B(n_1426),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1484),
.A2(n_1421),
.B(n_1413),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1474),
.B(n_1428),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1524),
.B(n_1421),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1548),
.B(n_1421),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1534),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1538),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1530),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1542),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1543),
.B(n_1484),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1548),
.B(n_1510),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1537),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1529),
.B(n_1493),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1548),
.B(n_1555),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1534),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1516),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1548),
.B(n_1513),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1531),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1553),
.A2(n_1491),
.B(n_1406),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1555),
.B(n_1502),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_SL g1572 ( 
.A1(n_1538),
.A2(n_1469),
.B(n_1523),
.C(n_1470),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1530),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1555),
.B(n_1491),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1544),
.A2(n_1471),
.B1(n_1496),
.B2(n_1494),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1494),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1551),
.A2(n_1473),
.B1(n_1470),
.B2(n_1478),
.C(n_1480),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1553),
.A2(n_1471),
.B1(n_1473),
.B2(n_1480),
.C(n_1478),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1544),
.A2(n_1519),
.B(n_1508),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1542),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1532),
.Y(n_1581)
);

NOR2xp67_ASAP7_75t_L g1582 ( 
.A(n_1531),
.B(n_1492),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1541),
.B(n_1509),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1483),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1479),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1551),
.B(n_1521),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1509),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1558),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1576),
.B(n_1564),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1565),
.B(n_1574),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1581),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1574),
.B(n_1545),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1577),
.A2(n_1551),
.B1(n_1482),
.B2(n_1518),
.C(n_1481),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1558),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1581),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1564),
.B(n_1561),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1561),
.B(n_1550),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1562),
.B(n_1549),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1564),
.B(n_1554),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1556),
.B(n_1540),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1546),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1584),
.B(n_1533),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1559),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1569),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1557),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1585),
.B(n_1567),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1560),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1559),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1550),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1573),
.Y(n_1614)
);

NOR4xp25_ASAP7_75t_SL g1615 ( 
.A(n_1586),
.B(n_1525),
.C(n_1504),
.D(n_1533),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1507),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1573),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1611),
.B(n_1579),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1608),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1605),
.B(n_1489),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1617),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1583),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1594),
.A2(n_1575),
.B1(n_1578),
.B2(n_1577),
.Y(n_1623)
);

AOI21xp33_ASAP7_75t_L g1624 ( 
.A1(n_1594),
.A2(n_1575),
.B(n_1586),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1599),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1607),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1598),
.B(n_1568),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1607),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1598),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1599),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1632)
);

INVxp67_ASAP7_75t_SL g1633 ( 
.A(n_1591),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1588),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1617),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1606),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1590),
.B(n_1600),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1588),
.B(n_1571),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1591),
.B(n_1563),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1616),
.A2(n_1578),
.B(n_1544),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1609),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1590),
.B(n_1583),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1600),
.B(n_1602),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1600),
.B(n_1583),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1563),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1612),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1612),
.Y(n_1653)
);

OAI31xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1615),
.A2(n_1572),
.A3(n_1515),
.B(n_1549),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1614),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1602),
.B(n_1587),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1614),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1595),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1624),
.B(n_1595),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1621),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1610),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1654),
.B(n_1624),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1625),
.Y(n_1664)
);

AND3x1_ASAP7_75t_L g1665 ( 
.A(n_1654),
.B(n_1615),
.C(n_1579),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1604),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1634),
.B(n_1610),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1642),
.B(n_1635),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1649),
.Y(n_1670)
);

NAND3xp33_ASAP7_75t_L g1671 ( 
.A(n_1642),
.B(n_1572),
.C(n_1544),
.Y(n_1671)
);

OAI31xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1630),
.A2(n_1499),
.A3(n_1604),
.B(n_1593),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1618),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1618),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1621),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1620),
.B(n_1487),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1627),
.B(n_1451),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1604),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1633),
.B(n_1613),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1604),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1638),
.B(n_1627),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1636),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1625),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1637),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1626),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1628),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_SL g1688 ( 
.A(n_1618),
.B(n_1451),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1618),
.A2(n_1570),
.B1(n_1549),
.B2(n_1552),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1638),
.B(n_1456),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1618),
.A2(n_1536),
.B1(n_1540),
.B2(n_1486),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1637),
.Y(n_1692)
);

NOR2xp67_ASAP7_75t_L g1693 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1661),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1695)
);

AND4x1_ASAP7_75t_L g1696 ( 
.A(n_1671),
.B(n_1511),
.C(n_1650),
.D(n_1641),
.Y(n_1696)
);

OAI322xp33_ASAP7_75t_L g1697 ( 
.A1(n_1663),
.A2(n_1632),
.A3(n_1629),
.B1(n_1641),
.B2(n_1650),
.C1(n_1644),
.C2(n_1603),
.Y(n_1697)
);

CKINVDCx14_ASAP7_75t_R g1698 ( 
.A(n_1676),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1661),
.Y(n_1699)
);

NAND2xp33_ASAP7_75t_SL g1700 ( 
.A(n_1659),
.B(n_1456),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1693),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_SL g1702 ( 
.A(n_1671),
.B(n_1492),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1665),
.A2(n_1570),
.B1(n_1536),
.B2(n_1552),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1670),
.B(n_1656),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1678),
.B(n_1681),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1678),
.B(n_1656),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1669),
.A2(n_1536),
.B(n_1456),
.C(n_1468),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1660),
.B(n_1632),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1690),
.A2(n_1570),
.B1(n_1552),
.B2(n_1540),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1665),
.A2(n_1640),
.B1(n_1644),
.B2(n_1646),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1672),
.A2(n_1580),
.B1(n_1611),
.B2(n_1603),
.C(n_1652),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1675),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1681),
.B(n_1622),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1675),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1686),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1687),
.A2(n_1570),
.B1(n_1552),
.B2(n_1535),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1686),
.B(n_1622),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1672),
.B(n_1646),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1698),
.B(n_1679),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1693),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1715),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1702),
.A2(n_1677),
.B1(n_1688),
.B2(n_1689),
.Y(n_1723)
);

XOR2xp5_ASAP7_75t_L g1724 ( 
.A(n_1698),
.B(n_1485),
.Y(n_1724)
);

OAI321xp33_ASAP7_75t_L g1725 ( 
.A1(n_1710),
.A2(n_1674),
.A3(n_1682),
.B1(n_1691),
.B2(n_1668),
.C(n_1662),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1701),
.B(n_1658),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1694),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1699),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1708),
.B(n_1682),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1696),
.A2(n_1688),
.B1(n_1674),
.B2(n_1662),
.C(n_1668),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1695),
.B(n_1658),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1712),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1711),
.A2(n_1673),
.B1(n_1667),
.B2(n_1666),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1705),
.Y(n_1734)
);

AND3x1_ASAP7_75t_L g1735 ( 
.A(n_1707),
.B(n_1673),
.C(n_1667),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_1666),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1719),
.A2(n_1673),
.B1(n_1648),
.B2(n_1603),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1700),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1714),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1697),
.B(n_1700),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1720),
.B(n_1704),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_SL g1742 ( 
.A(n_1740),
.B(n_1707),
.C(n_1703),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1722),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1720),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1740),
.A2(n_1716),
.B(n_1673),
.C(n_1709),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1724),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1722),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1734),
.B(n_1704),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1721),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1730),
.A2(n_1718),
.B1(n_1705),
.B2(n_1706),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1725),
.A2(n_1717),
.B1(n_1713),
.B2(n_1706),
.C(n_1692),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1735),
.A2(n_1713),
.B1(n_1580),
.B2(n_1685),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1744),
.B(n_1726),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1752),
.B(n_1738),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1743),
.B(n_1731),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1747),
.B(n_1736),
.Y(n_1756)
);

CKINVDCx16_ASAP7_75t_R g1757 ( 
.A(n_1741),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1752),
.B(n_1723),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1748),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1749),
.B(n_1729),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1750),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1758),
.A2(n_1742),
.B1(n_1733),
.B2(n_1737),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1755),
.Y(n_1763)
);

OAI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1754),
.A2(n_1746),
.B1(n_1728),
.B2(n_1727),
.Y(n_1764)
);

OAI211xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1753),
.A2(n_1745),
.B(n_1751),
.C(n_1739),
.Y(n_1765)
);

NAND4xp25_ASAP7_75t_L g1766 ( 
.A(n_1760),
.B(n_1756),
.C(n_1732),
.D(n_1757),
.Y(n_1766)
);

A2O1A1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1762),
.A2(n_1761),
.B(n_1759),
.C(n_1692),
.Y(n_1767)
);

AOI21xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1764),
.A2(n_1683),
.B(n_1680),
.Y(n_1768)
);

AOI22x1_ASAP7_75t_L g1769 ( 
.A1(n_1763),
.A2(n_1685),
.B1(n_1683),
.B2(n_1684),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1765),
.A2(n_1684),
.B1(n_1664),
.B2(n_1625),
.C(n_1631),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1766),
.A2(n_1684),
.B(n_1664),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1764),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1772),
.B(n_1664),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1767),
.A2(n_1768),
.B1(n_1770),
.B2(n_1771),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1769),
.A2(n_1657),
.B1(n_1655),
.B2(n_1653),
.Y(n_1775)
);

NAND4xp75_ASAP7_75t_L g1776 ( 
.A(n_1772),
.B(n_1582),
.C(n_1528),
.D(n_1481),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1771),
.B(n_1648),
.Y(n_1777)
);

AOI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1774),
.A2(n_1643),
.B(n_1631),
.Y(n_1778)
);

AOI32xp33_ASAP7_75t_L g1779 ( 
.A1(n_1777),
.A2(n_1580),
.A3(n_1619),
.B1(n_1450),
.B2(n_1453),
.Y(n_1779)
);

NOR3xp33_ASAP7_75t_L g1780 ( 
.A(n_1773),
.B(n_1453),
.C(n_1450),
.Y(n_1780)
);

XNOR2x1_ASAP7_75t_L g1781 ( 
.A(n_1780),
.B(n_1776),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1778),
.B1(n_1775),
.B2(n_1779),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1782),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1782),
.A2(n_1619),
.B1(n_1643),
.B2(n_1631),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1783),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_SL g1786 ( 
.A1(n_1784),
.A2(n_1520),
.B1(n_1527),
.B2(n_1485),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1785),
.A2(n_1645),
.B(n_1643),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1786),
.B1(n_1619),
.B2(n_1645),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1788),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1789),
.Y(n_1790)
);

OAI221xp5_ASAP7_75t_R g1791 ( 
.A1(n_1790),
.A2(n_1619),
.B1(n_1592),
.B2(n_1596),
.C(n_1466),
.Y(n_1791)
);

AOI211xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1527),
.B(n_1512),
.C(n_1485),
.Y(n_1792)
);


endmodule