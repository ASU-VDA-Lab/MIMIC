module real_aes_1475_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_769;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_0), .B(n_144), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_1), .A2(n_126), .B(n_177), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_2), .A2(n_451), .B1(n_456), .B2(n_801), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_3), .B(n_447), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_4), .A2(n_11), .B1(n_111), .B2(n_112), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_4), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_5), .B(n_134), .Y(n_190) );
INVx1_ASAP7_75t_L g131 ( .A(n_6), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_7), .B(n_134), .Y(n_154) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_8), .A2(n_104), .B1(n_444), .B2(n_449), .C1(n_809), .C2(n_814), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_8), .A2(n_106), .B1(n_430), .B2(n_431), .Y(n_105) );
INVxp67_ASAP7_75t_L g431 ( .A(n_8), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_8), .B(n_121), .Y(n_492) );
INVx1_ASAP7_75t_L g520 ( .A(n_9), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_10), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_11), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_12), .Y(n_535) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_13), .B(n_138), .Y(n_171) );
INVx2_ASAP7_75t_L g123 ( .A(n_14), .Y(n_123) );
AOI221x1_ASAP7_75t_L g213 ( .A1(n_15), .A2(n_28), .B1(n_126), .B2(n_144), .C(n_214), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_16), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_17), .B(n_144), .Y(n_167) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_18), .A2(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g501 ( .A(n_19), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_20), .B(n_157), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_21), .B(n_134), .Y(n_133) );
AO21x1_ASAP7_75t_L g185 ( .A1(n_22), .A2(n_144), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g439 ( .A(n_23), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_24), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g499 ( .A(n_25), .Y(n_499) );
INVx1_ASAP7_75t_SL g485 ( .A(n_26), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_27), .B(n_145), .Y(n_579) );
NAND2x1_ASAP7_75t_L g199 ( .A(n_29), .B(n_134), .Y(n_199) );
AOI33xp33_ASAP7_75t_L g547 ( .A1(n_30), .A2(n_55), .A3(n_475), .B1(n_482), .B2(n_548), .B3(n_549), .Y(n_547) );
NAND2x1_ASAP7_75t_L g153 ( .A(n_31), .B(n_138), .Y(n_153) );
INVx1_ASAP7_75t_L g529 ( .A(n_32), .Y(n_529) );
OR2x2_ASAP7_75t_L g122 ( .A(n_33), .B(n_89), .Y(n_122) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_33), .A2(n_89), .B(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_34), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_35), .B(n_138), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_36), .B(n_134), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_37), .B(n_138), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_38), .A2(n_126), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g127 ( .A(n_39), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g142 ( .A(n_39), .B(n_131), .Y(n_142) );
INVx1_ASAP7_75t_L g481 ( .A(n_39), .Y(n_481) );
OR2x6_ASAP7_75t_L g437 ( .A(n_40), .B(n_438), .Y(n_437) );
XNOR2xp5_ASAP7_75t_L g452 ( .A(n_41), .B(n_453), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_42), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_43), .B(n_144), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_44), .B(n_473), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_45), .A2(n_121), .B1(n_161), .B2(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_46), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_47), .B(n_145), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_48), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_49), .B(n_138), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_50), .B(n_165), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_51), .B(n_145), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_52), .A2(n_126), .B(n_152), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_53), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_54), .B(n_138), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_56), .B(n_145), .Y(n_559) );
INVx1_ASAP7_75t_L g130 ( .A(n_57), .Y(n_130) );
INVx1_ASAP7_75t_L g140 ( .A(n_57), .Y(n_140) );
AND2x2_ASAP7_75t_L g560 ( .A(n_58), .B(n_157), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_59), .A2(n_76), .B1(n_473), .B2(n_479), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_60), .B(n_473), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_61), .B(n_134), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_62), .B(n_161), .Y(n_537) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_63), .A2(n_479), .B(n_510), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_64), .A2(n_126), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g495 ( .A(n_65), .Y(n_495) );
AO21x1_ASAP7_75t_L g187 ( .A1(n_66), .A2(n_126), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_67), .B(n_144), .Y(n_175) );
INVx1_ASAP7_75t_L g558 ( .A(n_68), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_69), .B(n_144), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_70), .A2(n_479), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g236 ( .A(n_71), .B(n_158), .Y(n_236) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g136 ( .A(n_72), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_73), .A2(n_99), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_73), .Y(n_454) );
AND2x2_ASAP7_75t_L g159 ( .A(n_74), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_75), .B(n_473), .Y(n_550) );
AND2x2_ASAP7_75t_L g488 ( .A(n_77), .B(n_160), .Y(n_488) );
INVx1_ASAP7_75t_L g496 ( .A(n_78), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_79), .A2(n_479), .B(n_484), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_80), .A2(n_479), .B(n_542), .C(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g440 ( .A(n_81), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_82), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g173 ( .A(n_83), .B(n_160), .Y(n_173) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_84), .B(n_160), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_85), .A2(n_479), .B1(n_545), .B2(n_546), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_86), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_86), .Y(n_108) );
XNOR2xp5_ASAP7_75t_L g451 ( .A(n_87), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g186 ( .A(n_88), .B(n_121), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_90), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g203 ( .A(n_91), .B(n_160), .Y(n_203) );
INVx1_ASAP7_75t_L g511 ( .A(n_92), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_93), .B(n_134), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_94), .A2(n_126), .B(n_132), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_95), .B(n_138), .Y(n_215) );
AND2x2_ASAP7_75t_L g551 ( .A(n_96), .B(n_160), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_97), .B(n_134), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_98), .A2(n_527), .B(n_528), .C(n_530), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_99), .Y(n_455) );
BUFx2_ASAP7_75t_L g448 ( .A(n_100), .Y(n_448) );
BUFx2_ASAP7_75t_SL g820 ( .A(n_100), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_101), .A2(n_126), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_102), .B(n_145), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_432), .B(n_441), .Y(n_104) );
INVx1_ASAP7_75t_L g430 ( .A(n_106), .Y(n_430) );
XNOR2x1_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_113), .A2(n_457), .B1(n_461), .B2(n_464), .Y(n_456) );
INVx2_ASAP7_75t_L g806 ( .A(n_113), .Y(n_806) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_328), .Y(n_113) );
NAND3xp33_ASAP7_75t_SL g114 ( .A(n_115), .B(n_240), .C(n_295), .Y(n_114) );
AOI221xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_180), .B1(n_204), .B2(n_208), .C(n_218), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_163), .Y(n_116) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_117), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g239 ( .A(n_117), .Y(n_239) );
AND2x2_ASAP7_75t_L g284 ( .A(n_117), .B(n_221), .Y(n_284) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_148), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g272 ( .A(n_119), .Y(n_272) );
INVx1_ASAP7_75t_L g282 ( .A(n_119), .Y(n_282) );
AO21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_146), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_120), .B(n_147), .Y(n_146) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_120), .A2(n_124), .B(n_146), .Y(n_246) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_121), .A2(n_167), .B(n_168), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_121), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_121), .B(n_141), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_121), .A2(n_509), .B(n_513), .Y(n_508) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_122), .B(n_123), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_143), .Y(n_124) );
AND2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
BUFx3_ASAP7_75t_L g477 ( .A(n_127), .Y(n_477) );
AND2x6_ASAP7_75t_L g138 ( .A(n_128), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g483 ( .A(n_128), .Y(n_483) );
AND2x4_ASAP7_75t_L g479 ( .A(n_129), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x4_ASAP7_75t_L g134 ( .A(n_130), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g475 ( .A(n_130), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_131), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_137), .B(n_141), .Y(n_132) );
INVxp67_ASAP7_75t_L g502 ( .A(n_134), .Y(n_502) );
AND2x4_ASAP7_75t_L g145 ( .A(n_135), .B(n_139), .Y(n_145) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVxp67_ASAP7_75t_L g500 ( .A(n_138), .Y(n_500) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_141), .A2(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_141), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_141), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_141), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_141), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_141), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_141), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_141), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_141), .A2(n_486), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_141), .A2(n_486), .B(n_520), .C(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g545 ( .A(n_141), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_141), .A2(n_486), .B(n_558), .C(n_559), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_141), .A2(n_579), .B(n_580), .Y(n_578) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g144 ( .A(n_142), .B(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_142), .Y(n_530) );
INVx1_ASAP7_75t_L g497 ( .A(n_145), .Y(n_497) );
OR2x2_ASAP7_75t_L g261 ( .A(n_148), .B(n_164), .Y(n_261) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_148), .B(n_207), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_148), .B(n_172), .Y(n_305) );
INVx2_ASAP7_75t_L g314 ( .A(n_148), .Y(n_314) );
AND2x2_ASAP7_75t_L g335 ( .A(n_148), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g419 ( .A(n_148), .B(n_238), .Y(n_419) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g247 ( .A(n_149), .B(n_172), .Y(n_247) );
AND2x2_ASAP7_75t_L g380 ( .A(n_149), .B(n_207), .Y(n_380) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_149), .Y(n_406) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_156), .B(n_159), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
AO21x2_ASAP7_75t_L g470 ( .A1(n_156), .A2(n_471), .B(n_488), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_157), .A2(n_175), .B(n_176), .Y(n_174) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_157), .A2(n_213), .B(n_217), .Y(n_212) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_157), .A2(n_213), .B(n_217), .Y(n_224) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g202 ( .A(n_160), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_160), .A2(n_202), .B1(n_526), .B2(n_531), .Y(n_525) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_161), .B(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_162), .Y(n_165) );
AND2x4_ASAP7_75t_L g334 ( .A(n_163), .B(n_335), .Y(n_334) );
AOI321xp33_ASAP7_75t_L g348 ( .A1(n_163), .A2(n_277), .A3(n_278), .B1(n_310), .B2(n_349), .C(n_352), .Y(n_348) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_172), .Y(n_163) );
BUFx3_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx2_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_164), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g271 ( .A(n_164), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g304 ( .A(n_164), .Y(n_304) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_165), .A2(n_518), .B(n_522), .Y(n_517) );
INVx2_ASAP7_75t_SL g542 ( .A(n_165), .Y(n_542) );
INVx5_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
NOR2x1_ASAP7_75t_SL g256 ( .A(n_172), .B(n_246), .Y(n_256) );
BUFx2_ASAP7_75t_L g351 ( .A(n_172), .Y(n_351) );
OR2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVxp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_193), .Y(n_181) );
NOR2xp33_ASAP7_75t_SL g249 ( .A(n_182), .B(n_250), .Y(n_249) );
NOR4xp25_ASAP7_75t_L g352 ( .A(n_182), .B(n_346), .C(n_350), .D(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g390 ( .A(n_182), .Y(n_390) );
AND2x2_ASAP7_75t_L g424 ( .A(n_182), .B(n_364), .Y(n_424) );
BUFx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g279 ( .A(n_184), .Y(n_279) );
OAI21x1_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_187), .B(n_191), .Y(n_184) );
INVx1_ASAP7_75t_L g192 ( .A(n_186), .Y(n_192) );
AOI33xp33_ASAP7_75t_L g420 ( .A1(n_193), .A2(n_222), .A3(n_253), .B1(n_269), .B2(n_375), .B3(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g210 ( .A(n_194), .B(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g220 ( .A(n_194), .B(n_221), .Y(n_220) );
BUFx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g227 ( .A(n_195), .Y(n_227) );
INVxp67_ASAP7_75t_L g308 ( .A(n_195), .Y(n_308) );
AND2x2_ASAP7_75t_L g364 ( .A(n_195), .B(n_229), .Y(n_364) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_202), .B(n_203), .Y(n_195) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_196), .A2(n_202), .B(n_203), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_201), .Y(n_196) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_202), .A2(n_230), .B(n_236), .Y(n_229) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_202), .A2(n_230), .B(n_236), .Y(n_265) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_202), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x2_ASAP7_75t_L g591 ( .A1(n_202), .A2(n_554), .B(n_560), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_204), .A2(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AND2x2_ASAP7_75t_L g373 ( .A(n_205), .B(n_247), .Y(n_373) );
AND3x2_ASAP7_75t_L g375 ( .A(n_205), .B(n_259), .C(n_314), .Y(n_375) );
INVx3_ASAP7_75t_SL g327 ( .A(n_206), .Y(n_327) );
INVx4_ASAP7_75t_L g221 ( .A(n_207), .Y(n_221) );
AND2x2_ASAP7_75t_L g259 ( .A(n_207), .B(n_246), .Y(n_259) );
INVxp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
BUFx2_ASAP7_75t_L g253 ( .A(n_211), .Y(n_253) );
AND2x4_ASAP7_75t_L g278 ( .A(n_211), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g341 ( .A(n_211), .B(n_229), .Y(n_341) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g311 ( .A(n_212), .Y(n_311) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_212), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_R g218 ( .A1(n_219), .A2(n_222), .B(n_226), .C(n_237), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_221), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_221), .B(n_238), .Y(n_399) );
INVx1_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g381 ( .A(n_223), .B(n_371), .Y(n_381) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_L g228 ( .A(n_224), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g250 ( .A(n_224), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g266 ( .A(n_224), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g299 ( .A(n_224), .B(n_279), .Y(n_299) );
AND2x4_ASAP7_75t_L g264 ( .A(n_225), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g288 ( .A(n_225), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g326 ( .A(n_225), .B(n_251), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_L g254 ( .A(n_227), .B(n_251), .Y(n_254) );
AND2x2_ASAP7_75t_L g269 ( .A(n_227), .B(n_229), .Y(n_269) );
BUFx2_ASAP7_75t_L g325 ( .A(n_227), .Y(n_325) );
AND2x2_ASAP7_75t_L g339 ( .A(n_227), .B(n_250), .Y(n_339) );
INVx2_ASAP7_75t_L g251 ( .A(n_229), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_231), .B(n_235), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g287 ( .A1(n_237), .A2(n_288), .B1(n_290), .B2(n_294), .Y(n_287) );
INVx2_ASAP7_75t_SL g318 ( .A(n_237), .Y(n_318) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g293 ( .A(n_238), .B(n_246), .Y(n_293) );
INVx1_ASAP7_75t_L g400 ( .A(n_239), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_273), .C(n_287), .Y(n_240) );
OAI221xp5_ASAP7_75t_SL g241 ( .A1(n_242), .A2(n_248), .B1(n_252), .B2(n_255), .C(n_257), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
INVxp67_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_245), .Y(n_429) );
INVx1_ASAP7_75t_L g392 ( .A(n_247), .Y(n_392) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_247), .B(n_271), .Y(n_402) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_251), .B(n_279), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OR2x2_ASAP7_75t_L g285 ( .A(n_253), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g363 ( .A(n_253), .Y(n_363) );
AND2x2_ASAP7_75t_L g298 ( .A(n_254), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g344 ( .A(n_256), .B(n_304), .Y(n_344) );
AND2x2_ASAP7_75t_L g421 ( .A(n_256), .B(n_419), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B1(n_269), .B2(n_270), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g280 ( .A(n_261), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx2_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
AND2x4_ASAP7_75t_L g310 ( .A(n_264), .B(n_311), .Y(n_310) );
OAI21xp33_ASAP7_75t_SL g340 ( .A1(n_264), .A2(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g367 ( .A(n_264), .B(n_325), .Y(n_367) );
INVx2_ASAP7_75t_L g289 ( .A(n_265), .Y(n_289) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_265), .Y(n_322) );
INVx1_ASAP7_75t_SL g346 ( .A(n_266), .Y(n_346) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g277 ( .A(n_268), .Y(n_277) );
AND2x4_ASAP7_75t_SL g371 ( .A(n_268), .B(n_289), .Y(n_371) );
AND2x2_ASAP7_75t_L g368 ( .A(n_271), .B(n_314), .Y(n_368) );
AND2x2_ASAP7_75t_L g394 ( .A(n_271), .B(n_380), .Y(n_394) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_272), .Y(n_316) );
INVx1_ASAP7_75t_L g336 ( .A(n_272), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_280), .B1(n_283), .B2(n_285), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_278), .B(n_289), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_278), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g417 ( .A(n_278), .Y(n_417) );
INVx2_ASAP7_75t_SL g342 ( .A(n_280), .Y(n_342) );
AND2x2_ASAP7_75t_L g354 ( .A(n_282), .B(n_314), .Y(n_354) );
INVx2_ASAP7_75t_L g360 ( .A(n_282), .Y(n_360) );
INVxp33_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_288), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g410 ( .A(n_288), .Y(n_410) );
INVx1_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_291), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g349 ( .A(n_293), .B(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_293), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_317), .C(n_320), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B1(n_302), .B2(n_306), .C(n_309), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g415 ( .A(n_300), .Y(n_415) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g384 ( .A(n_301), .B(n_350), .Y(n_384) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g315 ( .A(n_304), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g386 ( .A(n_306), .Y(n_386) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g383 ( .A(n_307), .Y(n_383) );
INVx1_ASAP7_75t_L g389 ( .A(n_308), .Y(n_389) );
OR2x2_ASAP7_75t_L g412 ( .A(n_308), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_SL g321 ( .A(n_311), .Y(n_321) );
AND2x2_ASAP7_75t_L g391 ( .A(n_311), .B(n_371), .Y(n_391) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_311), .B(n_324), .Y(n_423) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g428 ( .A(n_314), .Y(n_428) );
INVx1_ASAP7_75t_L g378 ( .A(n_316), .Y(n_378) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_323), .C(n_327), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_321), .B(n_371), .Y(n_395) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_324), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g332 ( .A(n_326), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g413 ( .A(n_326), .Y(n_413) );
NAND4xp75_ASAP7_75t_L g328 ( .A(n_329), .B(n_385), .C(n_401), .D(n_422), .Y(n_328) );
NOR3x1_ASAP7_75t_L g329 ( .A(n_330), .B(n_347), .C(n_369), .Y(n_329) );
NAND4xp75_ASAP7_75t_L g330 ( .A(n_331), .B(n_337), .C(n_340), .D(n_343), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g382 ( .A(n_333), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g407 ( .A(n_334), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_SL g396 ( .A(n_339), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_355), .Y(n_347) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_351), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .B(n_365), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI322xp33_ASAP7_75t_L g387 ( .A1(n_359), .A2(n_388), .A3(n_392), .B1(n_393), .B2(n_395), .C1(n_396), .C2(n_397), .Y(n_387) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_360), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_363), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_364), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B(n_374), .C(n_376), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_382), .B2(n_384), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_391), .Y(n_388) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_394), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g404 ( .A(n_399), .B(n_405), .Y(n_404) );
O2A1O1Ixp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_408), .C(n_411), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B1(n_416), .B2(n_418), .C(n_420), .Y(n_411) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_432), .A2(n_446), .B(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g443 ( .A(n_434), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
AND2x6_ASAP7_75t_SL g460 ( .A(n_435), .B(n_437), .Y(n_460) );
OR2x6_ASAP7_75t_SL g463 ( .A(n_435), .B(n_436), .Y(n_463) );
OR2x2_ASAP7_75t_L g802 ( .A(n_435), .B(n_437), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g810 ( .A(n_443), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx2_ASAP7_75t_L g813 ( .A(n_446), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g812 ( .A(n_448), .B(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_450), .B(n_803), .Y(n_449) );
INVx1_ASAP7_75t_L g804 ( .A(n_451), .Y(n_804) );
CKINVDCx6p67_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
INVx4_ASAP7_75t_SL g807 ( .A(n_458), .Y(n_807) );
INVx3_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
CKINVDCx11_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
OAI22x1_ASAP7_75t_L g805 ( .A1(n_463), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_464), .Y(n_808) );
OR3x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_666), .C(n_737), .Y(n_464) );
NAND3x1_ASAP7_75t_SL g465 ( .A(n_466), .B(n_593), .C(n_615), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_583), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_514), .B1(n_561), .B2(n_565), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_468), .A2(n_769), .B1(n_770), .B2(n_772), .Y(n_768) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_489), .Y(n_468) );
AND2x2_ASAP7_75t_L g584 ( .A(n_469), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_469), .B(n_631), .Y(n_650) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g568 ( .A(n_470), .Y(n_568) );
AND2x2_ASAP7_75t_L g618 ( .A(n_470), .B(n_491), .Y(n_618) );
INVx1_ASAP7_75t_L g657 ( .A(n_470), .Y(n_657) );
OR2x2_ASAP7_75t_L g694 ( .A(n_470), .B(n_506), .Y(n_694) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_470), .Y(n_706) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_470), .Y(n_730) );
AND2x2_ASAP7_75t_L g787 ( .A(n_470), .B(n_614), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_478), .Y(n_471) );
INVx1_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_477), .Y(n_473) );
INVx1_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
OR2x6_ASAP7_75t_L g486 ( .A(n_475), .B(n_483), .Y(n_486) );
INVxp33_ASAP7_75t_L g548 ( .A(n_475), .Y(n_548) );
INVx1_ASAP7_75t_L g575 ( .A(n_477), .Y(n_575) );
INVxp67_ASAP7_75t_L g536 ( .A(n_479), .Y(n_536) );
NOR2x1p5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g549 ( .A(n_482), .Y(n_549) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_486), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
INVxp67_ASAP7_75t_L g527 ( .A(n_486), .Y(n_527) );
INVx2_ASAP7_75t_L g581 ( .A(n_486), .Y(n_581) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_504), .Y(n_489) );
INVx1_ASAP7_75t_L g662 ( .A(n_490), .Y(n_662) );
AND2x2_ASAP7_75t_L g688 ( .A(n_490), .B(n_506), .Y(n_688) );
NAND2x1_ASAP7_75t_L g704 ( .A(n_490), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g585 ( .A(n_491), .B(n_571), .Y(n_585) );
INVx3_ASAP7_75t_L g614 ( .A(n_491), .Y(n_614) );
NOR2x1_ASAP7_75t_SL g733 ( .A(n_491), .B(n_506), .Y(n_733) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .B(n_503), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_497), .B(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_501), .B2(n_502), .Y(n_498) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_504), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g612 ( .A(n_505), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx4_ASAP7_75t_L g582 ( .A(n_506), .Y(n_582) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_506), .Y(n_627) );
AND2x2_ASAP7_75t_L g699 ( .A(n_506), .B(n_571), .Y(n_699) );
AND2x4_ASAP7_75t_L g716 ( .A(n_506), .B(n_660), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_506), .B(n_658), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_506), .B(n_567), .Y(n_792) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_514), .A2(n_609), .B1(n_680), .B2(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_539), .Y(n_514) );
INVx2_ASAP7_75t_L g682 ( .A(n_515), .Y(n_682) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_523), .Y(n_515) );
BUFx3_ASAP7_75t_L g672 ( .A(n_516), .Y(n_672) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_517), .B(n_541), .Y(n_564) );
INVx2_ASAP7_75t_L g588 ( .A(n_517), .Y(n_588) );
INVx1_ASAP7_75t_L g600 ( .A(n_517), .Y(n_600) );
AND2x4_ASAP7_75t_L g607 ( .A(n_517), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g624 ( .A(n_517), .B(n_524), .Y(n_624) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_517), .Y(n_638) );
INVxp67_ASAP7_75t_L g646 ( .A(n_517), .Y(n_646) );
AND2x2_ASAP7_75t_L g675 ( .A(n_523), .B(n_591), .Y(n_675) );
AND2x2_ASAP7_75t_L g691 ( .A(n_523), .B(n_592), .Y(n_691) );
NOR2xp67_ASAP7_75t_L g778 ( .A(n_523), .B(n_591), .Y(n_778) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g587 ( .A(n_524), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g598 ( .A(n_524), .Y(n_598) );
INVx1_ASAP7_75t_L g611 ( .A(n_524), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_524), .B(n_553), .Y(n_648) );
OR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_536), .B1(n_537), .B2(n_538), .Y(n_532) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g771 ( .A(n_539), .Y(n_771) );
AND2x4_ASAP7_75t_L g539 ( .A(n_540), .B(n_552), .Y(n_539) );
AND2x2_ASAP7_75t_L g645 ( .A(n_540), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
AND2x2_ASAP7_75t_L g776 ( .A(n_540), .B(n_591), .Y(n_776) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_541), .B(n_553), .Y(n_636) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_551), .Y(n_541) );
AO21x2_ASAP7_75t_L g592 ( .A1(n_542), .A2(n_543), .B(n_551), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_550), .Y(n_543) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g562 ( .A(n_552), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g751 ( .A(n_552), .B(n_672), .Y(n_751) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_553), .Y(n_665) );
AND2x2_ASAP7_75t_L g692 ( .A(n_553), .B(n_638), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g606 ( .A(n_562), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g622 ( .A(n_562), .Y(n_622) );
AND2x2_ASAP7_75t_L g710 ( .A(n_562), .B(n_587), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_562), .B(n_730), .Y(n_735) );
AND2x2_ASAP7_75t_L g745 ( .A(n_562), .B(n_624), .Y(n_745) );
OR2x2_ASAP7_75t_L g782 ( .A(n_562), .B(n_682), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_563), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g742 ( .A(n_563), .B(n_598), .Y(n_742) );
AND2x2_ASAP7_75t_L g758 ( .A(n_563), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g752 ( .A(n_564), .B(n_648), .Y(n_752) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g634 ( .A(n_566), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_566), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g732 ( .A(n_566), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_566), .B(n_613), .Y(n_757) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_567), .Y(n_604) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_568), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_569), .A2(n_602), .B1(n_620), .B2(n_623), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_569), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g736 ( .A(n_569), .Y(n_736) );
AND2x4_ASAP7_75t_SL g569 ( .A(n_570), .B(n_582), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g613 ( .A(n_571), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
INVx1_ASAP7_75t_L g660 ( .A(n_571), .Y(n_660) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .C(n_576), .Y(n_573) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_582), .Y(n_602) );
AND2x4_ASAP7_75t_L g659 ( .A(n_582), .B(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_L g720 ( .A(n_582), .B(n_689), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
AND2x2_ASAP7_75t_L g684 ( .A(n_584), .B(n_627), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g764 ( .A1(n_584), .A2(n_765), .B(n_766), .Y(n_764) );
INVx2_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_586), .A2(n_696), .B1(n_700), .B2(n_703), .Y(n_695) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_587), .Y(n_653) );
AND2x2_ASAP7_75t_L g663 ( .A(n_587), .B(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g702 ( .A(n_587), .Y(n_702) );
NAND2x1_ASAP7_75t_SL g727 ( .A(n_587), .B(n_596), .Y(n_727) );
AND2x2_ASAP7_75t_L g623 ( .A(n_589), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_591), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g596 ( .A(n_592), .Y(n_596) );
INVx2_ASAP7_75t_L g608 ( .A(n_592), .Y(n_608) );
AOI21xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_601), .B(n_605), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_596), .B(n_790), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_597), .A2(n_686), .B1(n_690), .B2(n_693), .Y(n_685) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
BUFx2_ASAP7_75t_L g790 ( .A(n_598), .Y(n_790) );
INVx1_ASAP7_75t_SL g797 ( .A(n_598), .Y(n_797) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_599), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OA21x2_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B(n_612), .Y(n_605) );
AND2x2_ASAP7_75t_L g609 ( .A(n_607), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g651 ( .A(n_607), .B(n_647), .Y(n_651) );
AND2x2_ASAP7_75t_L g766 ( .A(n_607), .B(n_664), .Y(n_766) );
AND2x2_ASAP7_75t_L g769 ( .A(n_607), .B(n_675), .Y(n_769) );
AND2x4_ASAP7_75t_L g777 ( .A(n_607), .B(n_778), .Y(n_777) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_609), .A2(n_732), .B(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g759 ( .A(n_611), .Y(n_759) );
AND2x2_ASAP7_75t_L g775 ( .A(n_611), .B(n_776), .Y(n_775) );
INVx4_ASAP7_75t_L g689 ( .A(n_613), .Y(n_689) );
INVx1_ASAP7_75t_L g658 ( .A(n_614), .Y(n_658) );
AND2x2_ASAP7_75t_L g680 ( .A(n_614), .B(n_633), .Y(n_680) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_639), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B(n_625), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g626 ( .A(n_618), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_SL g779 ( .A(n_618), .B(n_631), .Y(n_779) );
AND2x2_ASAP7_75t_L g800 ( .A(n_618), .B(n_716), .Y(n_800) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g726 ( .A(n_623), .Y(n_726) );
OAI21xp5_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_628), .B(n_635), .Y(n_625) );
OR2x6_ASAP7_75t_L g678 ( .A(n_627), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OR2x2_ASAP7_75t_L g701 ( .A(n_636), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g798 ( .A(n_636), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_637), .B(n_771), .Y(n_770) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_652), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_649), .B2(n_651), .Y(n_640) );
OR2x2_ASAP7_75t_L g712 ( .A(n_642), .B(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_644), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g718 ( .A(n_647), .Y(n_718) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_661), .B2(n_663), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
AND2x4_ASAP7_75t_SL g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g722 ( .A(n_662), .B(n_716), .Y(n_722) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_667), .B(n_707), .Y(n_666) );
NOR2xp67_ASAP7_75t_L g667 ( .A(n_668), .B(n_681), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_670), .B(n_676), .Y(n_668) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp33_ASAP7_75t_SL g746 ( .A1(n_678), .A2(n_747), .B1(n_749), .B2(n_752), .Y(n_746) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_679), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g729 ( .A(n_680), .B(n_730), .Y(n_729) );
OAI211xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B(n_685), .C(n_695), .Y(n_681) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVxp33_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g698 ( .A(n_689), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_690), .A2(n_710), .B1(n_711), .B2(n_714), .C(n_717), .Y(n_709) );
AND2x4_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g750 ( .A(n_691), .Y(n_750) );
INVx2_ASAP7_75t_SL g748 ( .A(n_694), .Y(n_748) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NAND2x1_ASAP7_75t_L g747 ( .A(n_698), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g744 ( .A(n_704), .Y(n_744) );
INVx1_ASAP7_75t_L g773 ( .A(n_705), .Y(n_773) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_723), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_721), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g762 ( .A(n_713), .Y(n_762) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g783 ( .A(n_716), .B(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g788 ( .A(n_716), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVxp33_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g741 ( .A(n_720), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g723 ( .A1(n_724), .A2(n_728), .B(n_731), .Y(n_723) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g784 ( .A(n_730), .Y(n_784) );
AND2x2_ASAP7_75t_L g772 ( .A(n_733), .B(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_R g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_753), .C(n_780), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_746), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_740), .B(n_743), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_767), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_755), .B(n_764), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_756), .A2(n_758), .B1(n_760), .B2(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_763), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_768), .B(n_774), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_777), .B(n_779), .Y(n_774) );
INVx1_ASAP7_75t_L g793 ( .A(n_777), .Y(n_793) );
AOI211xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_783), .B(n_785), .C(n_794), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_789), .B1(n_791), .B2(n_793), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_799), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
INVxp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVxp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
CKINVDCx11_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
CKINVDCx8_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
endmodule