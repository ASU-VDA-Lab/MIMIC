module fake_jpeg_19351_n_201 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_31),
.B1(n_34),
.B2(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_16),
.B1(n_23),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_50),
.B1(n_55),
.B2(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_29),
.B(n_18),
.C(n_27),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_25),
.B(n_21),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_39),
.B1(n_36),
.B2(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_60),
.B1(n_66),
.B2(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_39),
.B1(n_36),
.B2(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_75),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_36),
.B1(n_33),
.B2(n_31),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_70)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_80),
.B(n_7),
.Y(n_112)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_87),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_38),
.B1(n_30),
.B2(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_84),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_12),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_62),
.B1(n_73),
.B2(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_4),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_6),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_80),
.B(n_83),
.C(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_131),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_81),
.B(n_71),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_122),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_75),
.B1(n_61),
.B2(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_120),
.B1(n_123),
.B2(n_93),
.Y(n_137)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_88),
.C(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_12),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_126),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_10),
.C(n_11),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_127),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_10),
.C(n_11),
.Y(n_127)
);

AOI22x1_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_11),
.B1(n_112),
.B2(n_111),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_104),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_110),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_96),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_117),
.B(n_123),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_91),
.B1(n_94),
.B2(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_89),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_93),
.B1(n_98),
.B2(n_96),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_149),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_109),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_154),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_116),
.B(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_138),
.B1(n_136),
.B2(n_121),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_141),
.B(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_148),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_129),
.A3(n_121),
.B1(n_114),
.B2(n_127),
.C1(n_119),
.C2(n_109),
.Y(n_161)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_139),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_171),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_162),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_144),
.C(n_168),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_137),
.B1(n_135),
.B2(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_171),
.A2(n_159),
.B1(n_154),
.B2(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_163),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_160),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_164),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_180),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_153),
.B1(n_163),
.B2(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_164),
.B1(n_173),
.B2(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_178),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_187),
.C(n_175),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_190),
.B(n_188),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_167),
.B(n_182),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_174),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_191),
.A2(n_184),
.B(n_176),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_186),
.C(n_156),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_190),
.B1(n_152),
.B2(n_181),
.C(n_146),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_197),
.Y(n_201)
);


endmodule