module fake_jpeg_23417_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_19),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_2),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_16),
.B1(n_14),
.B2(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_29),
.B1(n_14),
.B2(n_24),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_12),
.B1(n_10),
.B2(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_19),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.C(n_26),
.Y(n_42)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_11),
.B1(n_30),
.B2(n_7),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_26),
.C(n_25),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_39),
.C(n_36),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_44),
.B(n_45),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_45)
);

AO21x2_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_11),
.B(n_39),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_33),
.B(n_13),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_50),
.C(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_40),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_36),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_43),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_53),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B(n_30),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_49),
.B1(n_6),
.B2(n_7),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_5),
.Y(n_61)
);


endmodule