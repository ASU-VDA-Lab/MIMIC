module fake_jpeg_13599_n_432 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_432);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_432;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_56),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_62),
.Y(n_136)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_58),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_61),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_35),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_64),
.B(n_73),
.Y(n_129)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_88),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_75),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_15),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_80),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_86),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_19),
.B(n_6),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_92),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_7),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_15),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_101),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_98),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_31),
.B(n_14),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_106),
.Y(n_127)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_9),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_109),
.Y(n_177)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_34),
.B(n_10),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_25),
.B(n_10),
.C(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_36),
.B(n_0),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_45),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_36),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_0),
.Y(n_145)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_73),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_37),
.B1(n_41),
.B2(n_30),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_119),
.A2(n_122),
.B1(n_181),
.B2(n_164),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_60),
.A2(n_37),
.B1(n_41),
.B2(n_30),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_33),
.B1(n_49),
.B2(n_40),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_123),
.A2(n_147),
.B1(n_152),
.B2(n_157),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_124),
.B(n_134),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_132),
.B(n_129),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_64),
.A2(n_51),
.B1(n_20),
.B2(n_32),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_133),
.B(n_165),
.C(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_45),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_33),
.B1(n_49),
.B2(n_40),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_141),
.A2(n_154),
.B1(n_163),
.B2(n_151),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_44),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_142),
.B(n_153),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_145),
.B(n_161),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_44),
.B1(n_38),
.B2(n_83),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_105),
.A2(n_38),
.B1(n_54),
.B2(n_28),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_67),
.A2(n_54),
.B1(n_20),
.B2(n_32),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_82),
.A2(n_51),
.B1(n_1),
.B2(n_3),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_58),
.A2(n_0),
.B1(n_4),
.B2(n_65),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_85),
.A2(n_4),
.B1(n_86),
.B2(n_70),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_104),
.A2(n_84),
.B1(n_100),
.B2(n_80),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_176),
.B1(n_178),
.B2(n_128),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_72),
.B(n_59),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_174),
.B(n_179),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g176 ( 
.A1(n_71),
.A2(n_68),
.B1(n_61),
.B2(n_89),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_72),
.B(n_97),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_116),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_61),
.A2(n_87),
.B1(n_77),
.B2(n_56),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_182),
.Y(n_280)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_184),
.Y(n_279)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_187),
.Y(n_281)
);

OR2x2_ASAP7_75t_SL g188 ( 
.A(n_133),
.B(n_129),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_188),
.B(n_193),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_154),
.B1(n_122),
.B2(n_165),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_189),
.A2(n_196),
.B1(n_205),
.B2(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_194),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_121),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_192),
.B(n_199),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_139),
.A2(n_150),
.B1(n_178),
.B2(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_136),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_127),
.B(n_114),
.C(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_195),
.B(n_206),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_130),
.A2(n_123),
.B1(n_133),
.B2(n_138),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_118),
.Y(n_197)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_203),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_156),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_200),
.B(n_210),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_135),
.Y(n_204)
);

BUFx24_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_119),
.B1(n_138),
.B2(n_146),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_213),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_117),
.B(n_126),
.Y(n_210)
);

INVx6_ASAP7_75t_SL g211 ( 
.A(n_150),
.Y(n_211)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_144),
.B(n_167),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_137),
.B(n_130),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_217),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_115),
.B(n_171),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_207),
.C(n_233),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_128),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_221),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_139),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_162),
.B(n_160),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_223),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_224),
.A2(n_235),
.B1(n_237),
.B2(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_160),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_115),
.B(n_158),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_236),
.Y(n_243)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_232),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_168),
.A2(n_120),
.B(n_158),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_220),
.B(n_224),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_142),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_227),
.B(n_212),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_129),
.A2(n_177),
.B(n_127),
.C(n_142),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_177),
.A2(n_134),
.B1(n_142),
.B2(n_154),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_127),
.B(n_114),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_240),
.Y(n_257)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_135),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_244),
.A2(n_281),
.B1(n_241),
.B2(n_255),
.Y(n_302)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_188),
.Y(n_246)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_246),
.A2(n_231),
.B(n_240),
.C(n_206),
.D(n_204),
.Y(n_291)
);

OAI21x1_ASAP7_75t_R g248 ( 
.A1(n_211),
.A2(n_189),
.B(n_184),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_248),
.A2(n_281),
.B(n_273),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_250),
.A2(n_186),
.B(n_201),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_234),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_268),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_278),
.B1(n_250),
.B2(n_261),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_207),
.B(n_219),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_265),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_198),
.B(n_218),
.C(n_203),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_235),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_282),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_185),
.B(n_239),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_225),
.B(n_218),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_221),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_285),
.B(n_292),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_229),
.A3(n_217),
.B1(n_223),
.B2(n_209),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_303),
.B(n_263),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_257),
.B(n_197),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_298),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_294),
.A2(n_307),
.B(n_279),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_202),
.B1(n_244),
.B2(n_248),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_302),
.B1(n_318),
.B2(n_252),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_249),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_301),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_245),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_300),
.A2(n_316),
.B1(n_280),
.B2(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_249),
.B(n_241),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_241),
.B(n_243),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_304),
.B(n_305),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_253),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_314),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_273),
.A2(n_277),
.B(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_243),
.B(n_259),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_271),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_258),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_264),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_317),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_248),
.A2(n_280),
.B1(n_276),
.B2(n_246),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_319),
.A2(n_294),
.B1(n_299),
.B2(n_316),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_330),
.B1(n_341),
.B2(n_300),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_266),
.A3(n_260),
.B1(n_269),
.B2(n_272),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_292),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_287),
.A2(n_260),
.B1(n_275),
.B2(n_274),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_SL g347 ( 
.A1(n_337),
.A2(n_343),
.B(n_302),
.C(n_307),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_304),
.A2(n_264),
.B(n_258),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_339),
.A2(n_340),
.B(n_342),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_303),
.A2(n_251),
.B(n_283),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_287),
.A2(n_275),
.B1(n_272),
.B2(n_247),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_286),
.A2(n_251),
.B(n_283),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_346),
.A2(n_356),
.B1(n_361),
.B2(n_363),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_347),
.A2(n_352),
.B(n_291),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_333),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_349),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_298),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_293),
.Y(n_350)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_297),
.C(n_301),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_358),
.Y(n_376)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_314),
.B(n_317),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_318),
.B1(n_290),
.B2(n_285),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_354),
.A2(n_364),
.B1(n_339),
.B2(n_342),
.Y(n_373)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_344),
.Y(n_355)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_297),
.C(n_296),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_309),
.C(n_289),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_344),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_360),
.Y(n_370)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_329),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_324),
.B(n_305),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_288),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_365),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_373),
.A2(n_375),
.B1(n_378),
.B2(n_371),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_362),
.B(n_329),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_382),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_364),
.A2(n_334),
.B1(n_331),
.B2(n_341),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_346),
.A2(n_334),
.B1(n_343),
.B2(n_331),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_377),
.A2(n_354),
.B1(n_347),
.B2(n_330),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_336),
.B1(n_323),
.B2(n_291),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_345),
.B(n_340),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_351),
.B(n_337),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_384),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_385),
.A2(n_347),
.B1(n_368),
.B2(n_361),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_345),
.B(n_365),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_392),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_367),
.B(n_357),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_372),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_373),
.A2(n_375),
.B(n_347),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_SL g399 ( 
.A(n_389),
.B(n_391),
.C(n_394),
.Y(n_399)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_348),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_359),
.Y(n_392)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_393),
.A2(n_377),
.B1(n_347),
.B2(n_370),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_338),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_379),
.C(n_358),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_379),
.C(n_376),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_371),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_400),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_370),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_401),
.A2(n_405),
.B1(n_387),
.B2(n_384),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_403),
.B1(n_385),
.B2(n_383),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_404),
.B(n_395),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_408),
.Y(n_414)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_407),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_389),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_383),
.C(n_393),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_411),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_386),
.C(n_382),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_412),
.A2(n_413),
.B1(n_397),
.B2(n_398),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_400),
.A2(n_388),
.B1(n_390),
.B2(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_408),
.Y(n_424)
);

NOR2x1_ASAP7_75t_R g418 ( 
.A(n_411),
.B(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_419),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_399),
.B(n_401),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_410),
.Y(n_421)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_421),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_414),
.B(n_407),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_423),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_413),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_424),
.A2(n_416),
.B(n_355),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_427),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_425),
.C(n_420),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_429),
.B(n_335),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_335),
.Y(n_432)
);


endmodule