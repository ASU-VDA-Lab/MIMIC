module fake_jpeg_20855_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_1),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_51),
.B(n_3),
.C(n_41),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_35),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_3),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_43),
.B1(n_34),
.B2(n_38),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_34),
.B1(n_42),
.B2(n_47),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_14),
.C(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_61),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_36),
.B1(n_4),
.B2(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_32),
.B1(n_7),
.B2(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_13),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_31),
.B1(n_10),
.B2(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_67),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_80),
.B1(n_81),
.B2(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_17),
.Y(n_79)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_60),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_88),
.Y(n_94)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_18),
.C(n_19),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_91),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_100),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.C(n_98),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_84),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_86),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_87),
.B1(n_77),
.B2(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_24),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_25),
.Y(n_108)
);


endmodule