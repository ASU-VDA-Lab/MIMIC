module fake_jpeg_11741_n_78 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_5),
.B(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_1),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_28),
.B(n_32),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_30),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_4),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_12),
.C(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_7),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_11),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_19),
.C(n_20),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_17),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_21),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.C(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_67),
.C(n_62),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_73),
.B(n_58),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_70),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_60),
.B(n_22),
.Y(n_78)
);


endmodule