module fake_jpeg_19530_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_44),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_46),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_27),
.B1(n_17),
.B2(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_27),
.B1(n_20),
.B2(n_31),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_65),
.B(n_67),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_75),
.Y(n_114)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_73),
.B1(n_76),
.B2(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_29),
.B(n_21),
.C(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_43),
.B1(n_17),
.B2(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_54),
.B(n_26),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_32),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_94),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_98),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_37),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_84),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_32),
.B1(n_23),
.B2(n_33),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_103),
.B1(n_109),
.B2(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_24),
.B1(n_25),
.B2(n_3),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_25),
.B1(n_24),
.B2(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_24),
.B1(n_25),
.B2(n_4),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_1),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_5),
.Y(n_125)
);

OAI22x1_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_133),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_70),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_143),
.B(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_135),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_80),
.C(n_85),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_137),
.C(n_149),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_68),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_85),
.B1(n_74),
.B2(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_142),
.B1(n_11),
.B2(n_12),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_106),
.B1(n_114),
.B2(n_118),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_83),
.B(n_66),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_84),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_146),
.B1(n_115),
.B2(n_122),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_102),
.A2(n_74),
.B1(n_66),
.B2(n_9),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_6),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_150),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_9),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_10),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_100),
.B(n_124),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_153),
.B(n_167),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_100),
.B(n_115),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_109),
.B(n_112),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_161),
.B(n_166),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_168),
.B1(n_131),
.B2(n_146),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_117),
.B(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_171),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_117),
.C(n_119),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_108),
.B(n_12),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_108),
.B(n_12),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_145),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_149),
.CI(n_141),
.CON(n_171),
.SN(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_138),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_176),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_125),
.C(n_147),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_183),
.B(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_126),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_130),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_189),
.B1(n_158),
.B2(n_154),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_161),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_11),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_155),
.B(n_153),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_13),
.C(n_171),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_164),
.C(n_160),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_196),
.Y(n_209)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_170),
.A3(n_155),
.B1(n_171),
.B2(n_156),
.C1(n_163),
.C2(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_199),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_198),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_172),
.B1(n_166),
.B2(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_157),
.C(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_178),
.C(n_177),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_188),
.C(n_191),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_157),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_166),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_182),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_215),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_184),
.B(n_175),
.C(n_181),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_207),
.B1(n_201),
.B2(n_198),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_183),
.B(n_187),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_195),
.B(n_202),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g216 ( 
.A(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_204),
.C(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_209),
.C(n_206),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_200),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_225),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_219),
.B(n_203),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_222),
.C(n_227),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_190),
.B1(n_199),
.B2(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_223),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_SL g234 ( 
.A(n_228),
.B(n_164),
.C(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_234),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_239),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_230),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_237),
.Y(n_243)
);

AOI21x1_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_240),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_236),
.B(n_234),
.C(n_213),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_227),
.B(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_13),
.Y(n_247)
);


endmodule