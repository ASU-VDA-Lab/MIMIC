module fake_aes_6254_n_700 (n_20, n_12, n_56, n_47, n_52, n_67, n_50, n_7, n_1, n_60, n_16, n_22, n_3, n_19, n_10, n_34, n_40, n_68, n_25, n_30, n_36, n_9, n_13, n_53, n_26, n_11, n_64, n_72, n_69, n_39, n_43, n_73, n_62, n_38, n_23, n_0, n_33, n_4, n_59, n_24, n_35, n_6, n_32, n_8, n_15, n_57, n_61, n_51, n_44, n_71, n_66, n_70, n_46, n_45, n_42, n_21, n_2, n_37, n_48, n_27, n_63, n_18, n_17, n_54, n_28, n_41, n_58, n_65, n_55, n_49, n_5, n_29, n_14, n_31, n_700, n_678);
input n_20;
input n_12;
input n_56;
input n_47;
input n_52;
input n_67;
input n_50;
input n_7;
input n_1;
input n_60;
input n_16;
input n_22;
input n_3;
input n_19;
input n_10;
input n_34;
input n_40;
input n_68;
input n_25;
input n_30;
input n_36;
input n_9;
input n_13;
input n_53;
input n_26;
input n_11;
input n_64;
input n_72;
input n_69;
input n_39;
input n_43;
input n_73;
input n_62;
input n_38;
input n_23;
input n_0;
input n_33;
input n_4;
input n_59;
input n_24;
input n_35;
input n_6;
input n_32;
input n_8;
input n_15;
input n_57;
input n_61;
input n_51;
input n_44;
input n_71;
input n_66;
input n_70;
input n_46;
input n_45;
input n_42;
input n_21;
input n_2;
input n_37;
input n_48;
input n_27;
input n_63;
input n_18;
input n_17;
input n_54;
input n_28;
input n_41;
input n_58;
input n_65;
input n_55;
input n_49;
input n_5;
input n_29;
input n_14;
input n_31;
output n_700;
output n_678;
wire n_107;
wire n_646;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_169;
wire n_384;
wire n_370;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_357;
wire n_74;
wire n_308;
wire n_518;
wire n_44;
wire n_394;
wire n_189;
wire n_681;
wire n_352;
wire n_226;
wire n_447;
wire n_66;
wire n_379;
wire n_535;
wire n_689;
wire n_595;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_475;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_436;
wire n_438;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_223;
wire n_405;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_534;
wire n_569;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_303;
wire n_502;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_340;
wire n_301;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_246;
wire n_676;
wire n_191;
wire n_143;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_555;
wire n_553;
wire n_135;
wire n_481;
wire n_621;
wire n_397;
wire n_315;
wire n_53;
wire n_213;
wire n_196;
wire n_293;
wire n_127;
wire n_312;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_155;
wire n_162;
wire n_114;
wire n_50;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_9;
wire n_428;
wire n_478;
wire n_178;
wire n_652;
wire n_678;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_699;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_441;
wire n_628;
wire n_425;
wire n_314;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_172;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_228;
wire n_671;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_599;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_362;
wire n_617;
wire n_688;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_152;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_491;
wire n_388;
wire n_266;
wire n_80;
wire n_632;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_326;
wire n_532;
wire n_635;
wire n_544;
wire n_576;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_493;
wire n_274;
wire n_150;
wire n_235;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_100;
wire n_299;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_147;
wire n_185;
wire n_367;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_212;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_435;
wire n_583;
wire n_64;
wire n_69;
wire n_248;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_119;
wire n_667;
wire n_503;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_79;
wire n_129;
wire n_611;
wire n_521;
wire n_157;
wire n_103;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_325;
wire n_273;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_163;
wire n_348;
wire n_96;
wire n_685;
wire n_669;
wire n_72;
wire n_77;
wire n_90;
wire n_594;
wire n_214;
wire n_167;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_413;
wire n_65;
wire n_537;
wire n_560;
wire n_525;
wire n_5;
wire n_496;
wire n_393;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_290;
wire n_217;
wire n_201;
wire n_277;
wire n_259;
wire n_612;
wire n_244;
wire n_666;
wire n_297;
wire n_276;
wire n_225;
wire n_631;
wire n_350;
wire n_208;
wire n_616;
wire n_523;
wire n_528;
wire n_419;
wire n_252;
wire n_519;
wire n_168;
wire n_271;
wire n_693;
wire n_94;
wire n_194;
wire n_282;
wire n_58;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_116;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_597;
wire n_554;
wire n_698;
wire n_257;
wire n_26;
wire n_203;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_146;
wire n_337;
wire n_32;
wire n_637;
wire n_641;
wire n_531;
wire n_93;
wire n_539;
wire n_406;
wire n_372;
wire n_467;
wire n_41;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_647;
wire n_445;
wire n_500;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_75;
wire n_82;
wire n_183;
wire n_550;
wire n_132;
wire n_643;
wire n_582;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_510;
wire n_360;
wire n_363;
wire n_427;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_437;
wire n_620;
wire n_89;
wire n_480;
wire n_130;
wire n_341;
wire n_310;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_136;
wire n_260;
wire n_580;
wire n_610;
wire n_222;
wire n_657;
wire n_381;
wire n_34;
wire n_142;
wire n_385;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_606;
wire n_190;
wire n_62;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_376;
wire n_694;
wire n_240;
wire n_459;
wire n_88;
wire n_568;
wire n_46;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_672;
wire n_87;
wire n_466;
wire n_207;
wire n_197;
wire n_81;
wire n_541;
wire n_572;
wire n_298;
wire n_112;
wire n_630;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_36;
wire n_416;
wire n_432;
wire n_465;
wire n_414;
wire n_680;
wire n_369;
wire n_469;
wire n_361;
wire n_237;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_591;
wire n_391;
wire n_241;
wire n_209;
wire n_84;
wire n_20;
wire n_449;
wire n_12;
wire n_412;
wire n_56;
wire n_455;
wire n_67;
wire n_504;
wire n_618;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_383;
wire n_202;
wire n_319;
wire n_542;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_508;
wire n_486;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_400;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_173;
wire n_488;
wire n_556;
wire n_382;
wire n_138;
wire n_60;
wire n_462;
wire n_573;
wire n_536;
wire n_474;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_505;
wire n_358;
wire n_92;
wire n_313;
wire n_333;
wire n_627;
wire n_589;
wire n_175;
wire n_128;
wire n_306;
wire n_415;
wire n_31;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_234;
wire n_607;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_349;
INVx1_ASAP7_75t_L g74 ( .A(n_10), .Y(n_74) );
BUFx2_ASAP7_75t_L g75 ( .A(n_19), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_10), .Y(n_76) );
HB1xp67_ASAP7_75t_L g77 ( .A(n_13), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_50), .Y(n_79) );
INVxp33_ASAP7_75t_L g80 ( .A(n_64), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_68), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_38), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_12), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_22), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_11), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_45), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_70), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_72), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_61), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_42), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_9), .Y(n_92) );
INVxp67_ASAP7_75t_L g93 ( .A(n_16), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_67), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_54), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_15), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_36), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_35), .Y(n_98) );
INVx1_ASAP7_75t_SL g99 ( .A(n_21), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_3), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_26), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_28), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_58), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_53), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_71), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_57), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_49), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_13), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_66), .Y(n_113) );
INVxp33_ASAP7_75t_L g114 ( .A(n_34), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_17), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
OR2x2_ASAP7_75t_L g119 ( .A(n_47), .B(n_43), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_37), .Y(n_120) );
INVx4_ASAP7_75t_R g121 ( .A(n_44), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_63), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_75), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_82), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_75), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_82), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_122), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_107), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_76), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_107), .Y(n_137) );
NOR2xp33_ASAP7_75t_R g138 ( .A(n_113), .B(n_27), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_107), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_77), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_90), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_74), .B(n_0), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_112), .Y(n_147) );
OR2x2_ASAP7_75t_L g148 ( .A(n_74), .B(n_0), .Y(n_148) );
NOR2xp67_ASAP7_75t_L g149 ( .A(n_81), .B(n_1), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_99), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_92), .B(n_2), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_99), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_108), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_98), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_98), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_98), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_93), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_93), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_88), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_80), .B(n_2), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_91), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_97), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_91), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_100), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_97), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_83), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
NAND2x1p5_ASAP7_75t_L g169 ( .A(n_146), .B(n_119), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_153), .B(n_84), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_125), .B(n_102), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_123), .B(n_114), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
OR2x2_ASAP7_75t_L g177 ( .A(n_123), .B(n_100), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
NAND3xp33_ASAP7_75t_L g179 ( .A(n_162), .B(n_83), .C(n_85), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_133), .B(n_94), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_133), .B(n_106), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_156), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_136), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_140), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_164), .A2(n_115), .B1(n_96), .B2(n_85), .Y(n_191) );
INVx5_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_156), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_150), .B(n_106), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_140), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_124), .B(n_94), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_164), .B(n_116), .Y(n_199) );
BUFx10_ASAP7_75t_L g200 ( .A(n_127), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_126), .B(n_95), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_131), .Y(n_206) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_152), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_149), .B(n_116), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_132), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_126), .B(n_95), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_131), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_131), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_132), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_129), .B(n_103), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_129), .B(n_103), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_130), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
NOR2xp33_ASAP7_75t_SL g218 ( .A(n_160), .B(n_119), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_148), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_137), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_130), .B(n_104), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_151), .B(n_96), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_158), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_135), .B(n_104), .Y(n_226) );
NOR3xp33_ASAP7_75t_L g227 ( .A(n_151), .B(n_117), .C(n_105), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_135), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_149), .B(n_117), .Y(n_229) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_139), .A2(n_105), .B1(n_111), .B2(n_118), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_139), .B(n_111), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_219), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_223), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g234 ( .A1(n_218), .A2(n_166), .B1(n_145), .B2(n_128), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_219), .B(n_163), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_223), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_220), .Y(n_238) );
NOR2xp33_ASAP7_75t_R g239 ( .A(n_200), .B(n_147), .Y(n_239) );
NOR3xp33_ASAP7_75t_SL g240 ( .A(n_179), .B(n_163), .C(n_161), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_220), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_220), .B(n_161), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_203), .B(n_159), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
NOR3xp33_ASAP7_75t_SL g245 ( .A(n_196), .B(n_159), .C(n_144), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_203), .B(n_144), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_230), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_192), .B(n_143), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_203), .B(n_143), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_230), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_167), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_177), .B(n_134), .Y(n_252) );
NOR3xp33_ASAP7_75t_SL g253 ( .A(n_171), .B(n_87), .C(n_89), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_230), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_216), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_172), .B(n_138), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g258 ( .A(n_200), .B(n_3), .Y(n_258) );
BUFx4f_ASAP7_75t_L g259 ( .A(n_169), .Y(n_259) );
NOR2x1p5_ASAP7_75t_L g260 ( .A(n_177), .B(n_172), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_207), .B(n_101), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_167), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_216), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_200), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_167), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_224), .B(n_120), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_174), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_169), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_228), .A2(n_118), .B1(n_109), .B2(n_110), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_224), .B(n_118), .Y(n_271) );
BUFx4f_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_182), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_174), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_182), .B(n_109), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_208), .B(n_109), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_208), .B(n_4), .Y(n_277) );
NOR3xp33_ASAP7_75t_SL g278 ( .A(n_198), .B(n_121), .C(n_5), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_202), .B(n_141), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_183), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_182), .Y(n_282) );
INVx5_ASAP7_75t_L g283 ( .A(n_212), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_185), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_175), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_202), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_225), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_170), .B(n_137), .Y(n_288) );
AND2x6_ASAP7_75t_SL g289 ( .A(n_208), .B(n_229), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_185), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_202), .Y(n_291) );
XOR2xp5_ASAP7_75t_L g292 ( .A(n_191), .B(n_4), .Y(n_292) );
NAND2x1_ASAP7_75t_L g293 ( .A(n_212), .B(n_121), .Y(n_293) );
BUFx6f_ASAP7_75t_SL g294 ( .A(n_229), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_199), .B(n_137), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_199), .B(n_191), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_227), .A2(n_141), .B1(n_137), .B2(n_7), .Y(n_298) );
NAND2xp33_ASAP7_75t_SL g299 ( .A(n_210), .B(n_141), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_180), .B(n_137), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_242), .A2(n_192), .B(n_222), .Y(n_301) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_264), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_244), .B(n_229), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_263), .A2(n_192), .B(n_184), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_244), .B(n_186), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_243), .B(n_193), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_267), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_235), .A2(n_231), .B(n_226), .C(n_205), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_287), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_250), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_239), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_280), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_239), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_250), .A2(n_254), .B1(n_247), .B2(n_255), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_281), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_243), .B(n_214), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_295), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g326 ( .A1(n_259), .A2(n_192), .B1(n_215), .B2(n_193), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_251), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_269), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_259), .A2(n_192), .B1(n_212), .B2(n_206), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_243), .Y(n_330) );
BUFx12f_ASAP7_75t_L g331 ( .A(n_233), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_293), .A2(n_168), .B(n_176), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_237), .Y(n_333) );
INVx5_ASAP7_75t_L g334 ( .A(n_282), .Y(n_334) );
BUFx12f_ASAP7_75t_L g335 ( .A(n_289), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_275), .A2(n_194), .B(n_197), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_272), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_286), .B(n_5), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_272), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_252), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_251), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_297), .A2(n_206), .B1(n_197), .B2(n_194), .C(n_211), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_277), .A2(n_211), .B1(n_168), .B2(n_173), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_235), .A2(n_176), .B1(n_173), .B2(n_188), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_262), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_285), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_260), .B(n_6), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_249), .B(n_6), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_285), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_257), .B(n_7), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_246), .A2(n_141), .B1(n_175), .B2(n_181), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_SL g353 ( .A1(n_288), .A2(n_181), .B(n_187), .C(n_188), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_262), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_347), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
CKINVDCx16_ASAP7_75t_R g358 ( .A(n_316), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_307), .B(n_249), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_340), .B(n_277), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_306), .B(n_291), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_303), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_307), .B(n_277), .Y(n_363) );
AO22x2_ASAP7_75t_L g364 ( .A1(n_339), .A2(n_292), .B1(n_276), .B2(n_236), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_334), .B(n_283), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_310), .B(n_234), .Y(n_366) );
OAI22xp5_ASAP7_75t_SL g367 ( .A1(n_316), .A2(n_298), .B1(n_271), .B2(n_266), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_334), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_303), .B(n_232), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_304), .A2(n_253), .B1(n_240), .B2(n_276), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_308), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_308), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_314), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_311), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_314), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_330), .B(n_276), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_333), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_319), .Y(n_382) );
INVx6_ASAP7_75t_L g383 ( .A(n_334), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_330), .B(n_238), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_338), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_331), .Y(n_386) );
INVx4_ASAP7_75t_SL g387 ( .A(n_340), .Y(n_387) );
NAND2xp33_ASAP7_75t_SL g388 ( .A(n_340), .B(n_258), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_358), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_364), .A2(n_341), .B1(n_309), .B2(n_261), .C(n_351), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_364), .A2(n_339), .B1(n_311), .B2(n_317), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_364), .A2(n_335), .B1(n_348), .B2(n_331), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_364), .A2(n_335), .B1(n_348), .B2(n_339), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_355), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_367), .A2(n_339), .B1(n_294), .B2(n_312), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_376), .A2(n_332), .B(n_305), .Y(n_396) );
AOI21x1_ASAP7_75t_L g397 ( .A1(n_382), .A2(n_332), .B(n_349), .Y(n_397) );
INVx11_ASAP7_75t_L g398 ( .A(n_386), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_359), .B(n_319), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_367), .A2(n_294), .B1(n_312), .B2(n_258), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_323), .B1(n_320), .B2(n_321), .Y(n_401) );
BUFx12f_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_366), .A2(n_323), .B1(n_320), .B2(n_321), .Y(n_403) );
OAI33xp33_ASAP7_75t_L g404 ( .A1(n_382), .A2(n_322), .A3(n_324), .B1(n_345), .B2(n_300), .B3(n_352), .Y(n_404) );
AO21x2_ASAP7_75t_L g405 ( .A1(n_362), .A2(n_353), .B(n_301), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_360), .A2(n_350), .B(n_347), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_383), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g412 ( .A1(n_375), .A2(n_324), .B(n_336), .Y(n_412) );
BUFx6f_ASAP7_75t_SL g413 ( .A(n_369), .Y(n_413) );
AOI21xp33_ASAP7_75t_L g414 ( .A1(n_375), .A2(n_326), .B(n_338), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_378), .A2(n_340), .B1(n_302), .B2(n_328), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_368), .B(n_328), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_379), .A2(n_245), .B(n_278), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_413), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_393), .A2(n_378), .B1(n_359), .B2(n_360), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_407), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_407), .B(n_379), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_408), .B(n_387), .Y(n_423) );
OAI321xp33_ASAP7_75t_L g424 ( .A1(n_392), .A2(n_373), .A3(n_298), .B1(n_360), .B2(n_279), .C(n_270), .Y(n_424) );
OAI332xp33_ASAP7_75t_L g425 ( .A1(n_394), .A2(n_358), .A3(n_381), .B1(n_361), .B2(n_337), .B3(n_380), .C1(n_384), .C2(n_241), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
BUFx2_ASAP7_75t_SL g427 ( .A(n_413), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
INVx4_ASAP7_75t_L g429 ( .A(n_413), .Y(n_429) );
OAI222xp33_ASAP7_75t_L g430 ( .A1(n_391), .A2(n_360), .B1(n_373), .B2(n_369), .C1(n_377), .C2(n_357), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_400), .A2(n_270), .B(n_388), .C(n_363), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_411), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_390), .B(n_299), .C(n_141), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_398), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_397), .A2(n_371), .B(n_248), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_411), .B(n_387), .Y(n_436) );
AO21x2_ASAP7_75t_L g437 ( .A1(n_397), .A2(n_371), .B(n_248), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_395), .A2(n_360), .B1(n_363), .B2(n_338), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_402), .Y(n_440) );
NOR2xp33_ASAP7_75t_R g441 ( .A(n_389), .B(n_302), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_401), .A2(n_343), .B1(n_337), .B2(n_299), .C(n_344), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g444 ( .A1(n_403), .A2(n_340), .B1(n_329), .B2(n_342), .C(n_369), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_391), .A2(n_394), .B1(n_415), .B2(n_416), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_409), .A2(n_356), .B(n_372), .Y(n_446) );
OAI33xp33_ASAP7_75t_L g447 ( .A1(n_416), .A2(n_327), .A3(n_354), .B1(n_213), .B2(n_217), .B3(n_14), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_398), .A2(n_369), .B1(n_383), .B2(n_365), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_417), .A2(n_338), .B1(n_383), .B2(n_357), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_399), .A2(n_338), .B1(n_377), .B2(n_370), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_412), .B(n_357), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_449), .B(n_439), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_449), .B(n_417), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_429), .B(n_413), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_419), .A2(n_445), .B1(n_429), .B2(n_427), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_443), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_427), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_453), .B(n_405), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_439), .B(n_412), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_420), .B(n_405), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_428), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_428), .B(n_405), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_432), .B(n_417), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_453), .B(n_405), .Y(n_467) );
AOI221xp5_ASAP7_75t_SL g468 ( .A1(n_430), .A2(n_414), .B1(n_357), .B2(n_377), .C(n_370), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_418), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_438), .A2(n_417), .B1(n_404), .B2(n_414), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_443), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_448), .B(n_421), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_448), .B(n_385), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_422), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_421), .B(n_385), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
NAND3xp33_ASAP7_75t_SL g477 ( .A(n_434), .B(n_365), .C(n_279), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_425), .A2(n_410), .B1(n_315), .B2(n_325), .C(n_318), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_447), .A2(n_410), .B1(n_383), .B2(n_377), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_422), .B(n_8), .C(n_9), .D(n_11), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_418), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_440), .B(n_370), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_440), .B(n_370), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_426), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
AOI221xp5_ASAP7_75t_SL g487 ( .A1(n_450), .A2(n_175), .B1(n_354), .B2(n_327), .C(n_315), .Y(n_487) );
INVx4_ASAP7_75t_L g488 ( .A(n_429), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_437), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_437), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_423), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_423), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_423), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_418), .Y(n_495) );
OAI33xp33_ASAP7_75t_L g496 ( .A1(n_434), .A2(n_8), .A3(n_12), .B1(n_14), .B2(n_16), .B3(n_18), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_436), .B(n_396), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_436), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_426), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_452), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_446), .B(n_356), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_444), .A2(n_365), .B1(n_315), .B2(n_318), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_431), .B(n_387), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_459), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_454), .B(n_451), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_459), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_485), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_467), .B(n_396), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_458), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_458), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_455), .B(n_433), .Y(n_512) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_456), .B(n_488), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_454), .B(n_442), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_467), .B(n_18), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_472), .B(n_19), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_500), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_464), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_463), .B(n_20), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_464), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_466), .B(n_472), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_462), .B(n_20), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_463), .B(n_175), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_459), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_474), .B(n_424), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_465), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_462), .B(n_175), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_465), .B(n_387), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_471), .B(n_356), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_471), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_460), .Y(n_532) );
AOI31xp33_ASAP7_75t_L g533 ( .A1(n_460), .A2(n_441), .A3(n_387), .B(n_273), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_481), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_456), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_493), .B(n_372), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_475), .B(n_325), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_475), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_461), .B(n_23), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_498), .B(n_325), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_493), .B(n_372), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_499), .B(n_318), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_461), .B(n_24), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_499), .B(n_372), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_461), .B(n_25), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_461), .B(n_29), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_493), .B(n_494), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_497), .B(n_31), .Y(n_551) );
INVx3_ASAP7_75t_SL g552 ( .A(n_456), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_473), .B(n_372), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_473), .B(n_356), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_469), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_494), .B(n_490), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_494), .B(n_356), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_491), .B(n_32), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_480), .B(n_342), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_457), .B(n_342), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_560), .A2(n_480), .B1(n_496), .B2(n_478), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_521), .B(n_491), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_513), .B(n_488), .Y(n_564) );
AOI322xp5_ASAP7_75t_L g565 ( .A1(n_508), .A2(n_468), .A3(n_470), .B1(n_477), .B2(n_487), .C1(n_501), .C2(n_482), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_517), .B(n_495), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_516), .B(n_484), .C(n_483), .Y(n_567) );
O2A1O1Ixp5_ASAP7_75t_L g568 ( .A1(n_525), .A2(n_488), .B(n_504), .C(n_503), .Y(n_568) );
OAI221xp5_ASAP7_75t_L g569 ( .A1(n_522), .A2(n_468), .B1(n_483), .B2(n_488), .C(n_487), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_508), .B(n_495), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_533), .A2(n_482), .B(n_479), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_513), .A2(n_502), .B1(n_492), .B2(n_490), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_515), .A2(n_502), .B(n_489), .Y(n_573) );
AOI32xp33_ASAP7_75t_L g574 ( .A1(n_515), .A2(n_476), .A3(n_486), .B1(n_346), .B2(n_265), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_505), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_511), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_514), .A2(n_486), .B1(n_476), .B2(n_502), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_552), .A2(n_346), .B1(n_283), .B2(n_265), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_532), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_518), .Y(n_580) );
NOR2xp33_ASAP7_75t_R g581 ( .A(n_552), .B(n_33), .Y(n_581) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_519), .A2(n_178), .B(n_195), .C(n_209), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_519), .B(n_39), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_539), .B(n_40), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_518), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_521), .B(n_41), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_535), .A2(n_283), .B1(n_350), .B2(n_347), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_561), .A2(n_283), .B1(n_273), .B2(n_209), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_527), .B(n_48), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_527), .B(n_52), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_535), .A2(n_195), .B1(n_209), .B2(n_178), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_544), .B(n_56), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_507), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_529), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_520), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_556), .Y(n_597) );
NAND4xp25_ASAP7_75t_SL g598 ( .A(n_551), .B(n_59), .C(n_60), .D(n_62), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_529), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_556), .B(n_65), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
AOI21xp33_ASAP7_75t_SL g602 ( .A1(n_551), .A2(n_213), .B(n_217), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_540), .A2(n_221), .B(n_187), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_540), .A2(n_546), .B1(n_548), .B2(n_549), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_550), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_506), .B(n_178), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_509), .B(n_178), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_546), .B(n_178), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_597), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_566), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_588), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_596), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_604), .A2(n_559), .B1(n_537), .B2(n_549), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_594), .Y(n_615) );
AO21x1_ASAP7_75t_L g616 ( .A1(n_564), .A2(n_548), .B(n_531), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_601), .B(n_509), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_605), .B(n_563), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_576), .Y(n_619) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_565), .A2(n_557), .B(n_512), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_573), .A2(n_557), .B(n_512), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_580), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_575), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_606), .B(n_523), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_585), .Y(n_625) );
OAI33xp33_ASAP7_75t_L g626 ( .A1(n_579), .A2(n_545), .A3(n_541), .B1(n_553), .B2(n_554), .B3(n_547), .Y(n_626) );
NAND2xp33_ASAP7_75t_R g627 ( .A(n_581), .B(n_524), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_575), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_607), .Y(n_629) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_570), .A2(n_528), .B(n_543), .C(n_538), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_595), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_562), .B(n_507), .Y(n_632) );
AOI22x1_ASAP7_75t_L g633 ( .A1(n_571), .A2(n_528), .B1(n_526), .B2(n_538), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_599), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_567), .B(n_526), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_577), .B(n_543), .Y(n_636) );
XOR2x2_ASAP7_75t_L g637 ( .A(n_567), .B(n_530), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_586), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_598), .B(n_530), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_574), .B(n_534), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_569), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_608), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_590), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_632), .B(n_562), .Y(n_644) );
NAND3xp33_ASAP7_75t_SL g645 ( .A(n_616), .B(n_582), .C(n_568), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_632), .B(n_572), .Y(n_646) );
AOI21xp33_ASAP7_75t_L g647 ( .A1(n_641), .A2(n_568), .B(n_583), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_620), .A2(n_591), .B1(n_600), .B2(n_584), .C(n_602), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_617), .B(n_558), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g650 ( .A1(n_621), .A2(n_609), .B(n_589), .Y(n_650) );
OAI21xp33_ASAP7_75t_L g651 ( .A1(n_637), .A2(n_603), .B(n_578), .Y(n_651) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_643), .A2(n_593), .B(n_587), .C(n_592), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_628), .B(n_542), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_611), .B(n_542), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_612), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_635), .B(n_536), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_626), .A2(n_587), .B(n_536), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_637), .B(n_629), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_626), .A2(n_350), .B(n_209), .Y(n_659) );
NOR2xp67_ASAP7_75t_SL g660 ( .A(n_627), .B(n_209), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_633), .A2(n_195), .B1(n_190), .B2(n_189), .Y(n_661) );
OA22x2_ASAP7_75t_L g662 ( .A1(n_627), .A2(n_189), .B1(n_190), .B2(n_201), .Y(n_662) );
XOR2x2_ASAP7_75t_L g663 ( .A(n_614), .B(n_195), .Y(n_663) );
XNOR2xp5_ASAP7_75t_L g664 ( .A(n_631), .B(n_201), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_630), .A2(n_195), .B1(n_285), .B2(n_274), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_613), .Y(n_666) );
NAND2xp33_ASAP7_75t_R g667 ( .A(n_660), .B(n_638), .Y(n_667) );
NAND2xp33_ASAP7_75t_R g668 ( .A(n_644), .B(n_638), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_658), .B(n_634), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_664), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_654), .B(n_646), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_657), .B(n_636), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_662), .Y(n_673) );
AOI21xp33_ASAP7_75t_SL g674 ( .A1(n_651), .A2(n_640), .B(n_623), .Y(n_674) );
NOR2xp33_ASAP7_75t_R g675 ( .A(n_645), .B(n_639), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_653), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_647), .A2(n_610), .B1(n_625), .B2(n_619), .C(n_622), .Y(n_677) );
UNKNOWN g678 ( );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_656), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_650), .A2(n_618), .B1(n_615), .B2(n_624), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g681 ( .A(n_652), .B(n_615), .C(n_642), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_655), .B(n_268), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_649), .B(n_268), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_666), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_661), .B(n_665), .C(n_659), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_663), .A2(n_651), .B(n_660), .C(n_644), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_675), .B(n_674), .C(n_680), .Y(n_687) );
AND3x4_ASAP7_75t_L g688 ( .A(n_678), .B(n_681), .C(n_685), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_668), .A2(n_673), .B1(n_686), .B2(n_672), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_670), .Y(n_690) );
NOR4xp25_ASAP7_75t_L g691 ( .A(n_677), .B(n_671), .C(n_676), .D(n_684), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_690), .Y(n_692) );
OR3x1_ASAP7_75t_L g693 ( .A(n_687), .B(n_668), .C(n_667), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_689), .B(n_682), .C(n_683), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_692), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_693), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_696), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_695), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_697), .A2(n_696), .B1(n_694), .B2(n_688), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_691), .B1(n_698), .B2(n_669), .C(n_679), .Y(n_700) );
endmodule