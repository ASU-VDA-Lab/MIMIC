module fake_jpeg_29650_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_31;
wire n_25;
wire n_17;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx6p67_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_13),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_37),
.Y(n_43)
);

OA21x2_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_21),
.B(n_14),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_36),
.B(n_21),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_19),
.B1(n_24),
.B2(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_21),
.B1(n_15),
.B2(n_11),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_33),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_35),
.C(n_37),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_39),
.B(n_28),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_49),
.B(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_15),
.Y(n_55)
);

AOI321xp33_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_7),
.A3(n_13),
.B1(n_17),
.B2(n_46),
.C(n_52),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_48),
.B(n_50),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_57),
.B(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);


endmodule