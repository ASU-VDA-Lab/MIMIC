module fake_jpeg_12430_n_569 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_569);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_569;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g155 ( 
.A(n_59),
.Y(n_155)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_8),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_60),
.B(n_42),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_63),
.Y(n_114)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_6),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_96),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_74),
.Y(n_157)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx4f_ASAP7_75t_SL g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_22),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_87),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_111),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_6),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_34),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_5),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_34),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_110),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_22),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_43),
.B1(n_52),
.B2(n_47),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_117),
.A2(n_174),
.B1(n_44),
.B2(n_36),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_120),
.B(n_134),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_97),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_137),
.B(n_148),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_102),
.B1(n_55),
.B2(n_48),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_138),
.A2(n_152),
.B1(n_87),
.B2(n_95),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_74),
.B(n_32),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_147),
.B(n_178),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_59),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_42),
.B1(n_48),
.B2(n_52),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_156),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_161),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_79),
.B(n_35),
.Y(n_161)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_37),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_177),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_79),
.A2(n_17),
.B(n_28),
.Y(n_172)
);

OR2x4_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_14),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_70),
.A2(n_44),
.B1(n_47),
.B2(n_52),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_35),
.Y(n_178)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_183),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_17),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_195),
.Y(n_252)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_185),
.Y(n_265)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_110),
.B1(n_85),
.B2(n_99),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_192),
.B(n_223),
.Y(n_280)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

CKINVDCx12_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_37),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_53),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_199),
.A2(n_211),
.B1(n_214),
.B2(n_182),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_53),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_200),
.B(n_201),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_121),
.B(n_122),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_38),
.B1(n_30),
.B2(n_48),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_204),
.A2(n_210),
.B1(n_227),
.B2(n_228),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_123),
.A2(n_54),
.B1(n_108),
.B2(n_105),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_205),
.A2(n_128),
.B(n_136),
.Y(n_268)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_209),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_30),
.B1(n_38),
.B2(n_31),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_152),
.A2(n_107),
.B1(n_109),
.B2(n_94),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_40),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_213),
.B(n_215),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_138),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_39),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_39),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_217),
.B(n_220),
.Y(n_274)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_219),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_124),
.B(n_36),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_239),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_141),
.B(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_226),
.B(n_236),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_157),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_157),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

CKINVDCx6p67_ASAP7_75t_R g232 ( 
.A(n_167),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_243),
.Y(n_275)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_233),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_162),
.Y(n_234)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_116),
.Y(n_235)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_2),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_172),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_237),
.B(n_238),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_119),
.B(n_0),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_140),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g244 ( 
.A(n_155),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_244),
.Y(n_251)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_144),
.B(n_4),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_247),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_135),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_126),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_158),
.B(n_143),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_250),
.A2(n_257),
.B(n_271),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_158),
.B(n_143),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_184),
.B(n_135),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_260),
.B(n_195),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_142),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_261),
.B(n_283),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_196),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_262),
.B(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_180),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_285),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_279),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_155),
.B(n_169),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_198),
.A2(n_128),
.B(n_168),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_205),
.A2(n_116),
.B(n_163),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_206),
.B(n_115),
.C(n_150),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_201),
.B(n_139),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_289),
.A2(n_302),
.B1(n_202),
.B2(n_224),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_200),
.A2(n_116),
.B1(n_132),
.B2(n_130),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_SL g340 ( 
.A(n_292),
.B(n_294),
.C(n_232),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_233),
.A2(n_230),
.B1(n_234),
.B2(n_245),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_247),
.A2(n_115),
.B1(n_132),
.B2(n_130),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_298),
.A2(n_183),
.B1(n_191),
.B2(n_219),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_222),
.A2(n_126),
.B1(n_139),
.B2(n_12),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_189),
.B(n_4),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_188),
.Y(n_306)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_300),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_308),
.A2(n_241),
.B(n_190),
.C(n_273),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_275),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_312),
.Y(n_382)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_285),
.Y(n_314)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_320),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_207),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_318),
.B(n_323),
.Y(n_365)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_319),
.B(n_338),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_213),
.Y(n_320)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_267),
.Y(n_322)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_322),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_251),
.B(n_186),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_215),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_325),
.Y(n_371)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_328),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_252),
.B(n_242),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_303),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_329),
.B(n_330),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_249),
.Y(n_330)
);

XOR2x2_ASAP7_75t_L g331 ( 
.A(n_261),
.B(n_264),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_342),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_248),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_333),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_216),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_334),
.B(n_337),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_264),
.A2(n_230),
.B1(n_234),
.B2(n_240),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_259),
.B(n_187),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_288),
.B(n_279),
.Y(n_359)
);

INVx6_ASAP7_75t_SL g341 ( 
.A(n_267),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_341),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_250),
.B(n_218),
.Y(n_342)
);

INVx13_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_343),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_232),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_348),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_345),
.A2(n_347),
.B1(n_355),
.B2(n_256),
.Y(n_396)
);

CKINVDCx12_ASAP7_75t_R g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_346),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_253),
.B(n_232),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_264),
.A2(n_191),
.B1(n_203),
.B2(n_185),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_349),
.A2(n_353),
.B1(n_257),
.B2(n_268),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_208),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_350),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_282),
.B(n_241),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_354),
.C(n_293),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_289),
.A2(n_235),
.B1(n_221),
.B2(n_193),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_241),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_302),
.A2(n_209),
.B1(n_225),
.B2(n_212),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_276),
.B(n_0),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_270),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_367),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_352),
.A2(n_271),
.B(n_280),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_369),
.Y(n_408)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_329),
.A2(n_280),
.A3(n_281),
.B1(n_304),
.B2(n_296),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_317),
.B(n_322),
.Y(n_409)
);

FAx1_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_281),
.CI(n_273),
.CON(n_375),
.SN(n_375)
);

A2O1A1O1Ixp25_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_354),
.B(n_342),
.C(n_351),
.D(n_317),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_341),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_377),
.B(n_384),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_314),
.A2(n_290),
.B1(n_255),
.B2(n_291),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_378),
.A2(n_381),
.B1(n_390),
.B2(n_395),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_330),
.A2(n_356),
.B1(n_310),
.B2(n_320),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_348),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_266),
.C(n_296),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_388),
.C(n_392),
.Y(n_406)
);

AO22x1_ASAP7_75t_SL g386 ( 
.A1(n_347),
.A2(n_265),
.B1(n_266),
.B2(n_277),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_345),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_258),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_310),
.A2(n_290),
.B1(n_291),
.B2(n_265),
.Y(n_390)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_339),
.B(n_277),
.C(n_258),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_331),
.B(n_270),
.C(n_293),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_342),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_327),
.A2(n_256),
.B1(n_0),
.B2(n_12),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_396),
.A2(n_355),
.B1(n_309),
.B2(n_319),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_332),
.B(n_4),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_312),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_374),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_412),
.Y(n_433)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_399),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_387),
.Y(n_437)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_328),
.A3(n_337),
.B1(n_336),
.B2(n_308),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_418),
.Y(n_436)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_404),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_405),
.B(n_414),
.C(n_427),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_407),
.A2(n_381),
.B(n_392),
.Y(n_453)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_324),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_379),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_416),
.Y(n_434)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_359),
.A2(n_349),
.B1(n_317),
.B2(n_311),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_419),
.B1(n_362),
.B2(n_394),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_316),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_367),
.A2(n_353),
.B1(n_340),
.B2(n_313),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_326),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_422),
.Y(n_446)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_428),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_334),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_387),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_425),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_365),
.B(n_333),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_424),
.B(n_426),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_318),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_321),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_325),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_376),
.B(n_315),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_315),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_431),
.Y(n_449)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_432),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g484 ( 
.A(n_437),
.B(n_322),
.C(n_338),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_375),
.Y(n_438)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_402),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_439),
.B(n_455),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_442),
.A2(n_463),
.B1(n_389),
.B2(n_357),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_429),
.A2(n_419),
.B1(n_413),
.B2(n_400),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_443),
.A2(n_458),
.B(n_459),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_393),
.Y(n_450)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_423),
.B(n_420),
.Y(n_451)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_451),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_427),
.B(n_364),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_393),
.Y(n_454)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_454),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_397),
.Y(n_457)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_457),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_413),
.A2(n_364),
.B(n_391),
.Y(n_458)
);

FAx1_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_395),
.CI(n_379),
.CON(n_459),
.SN(n_459)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_363),
.B(n_358),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_SL g468 ( 
.A1(n_461),
.A2(n_448),
.B(n_449),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_385),
.C(n_405),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_406),
.C(n_401),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_408),
.A2(n_378),
.B1(n_358),
.B2(n_386),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_471),
.C(n_478),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_468),
.A2(n_438),
.B(n_461),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_407),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_408),
.C(n_368),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_438),
.Y(n_475)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_416),
.Y(n_476)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_476),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_460),
.A2(n_429),
.B1(n_410),
.B2(n_411),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_477),
.A2(n_481),
.B1(n_463),
.B2(n_449),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_411),
.C(n_399),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_447),
.A2(n_431),
.B1(n_403),
.B2(n_386),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_479),
.A2(n_480),
.B1(n_486),
.B2(n_460),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_435),
.A2(n_373),
.B1(n_357),
.B2(n_346),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_434),
.Y(n_483)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_488),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_309),
.C(n_343),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_487),
.C(n_440),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_447),
.A2(n_372),
.B1(n_343),
.B2(n_13),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_372),
.C(n_0),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_372),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_489),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_469),
.B(n_442),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_490),
.B(n_480),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_458),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_441),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_500),
.C(n_504),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_469),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_501),
.Y(n_514)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_495),
.B(n_503),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_497),
.A2(n_507),
.B1(n_487),
.B2(n_498),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_441),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_443),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_437),
.Y(n_502)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_508),
.C(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_433),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_505),
.B(n_436),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g508 ( 
.A(n_475),
.B(n_436),
.CI(n_446),
.CON(n_508),
.SN(n_508)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_510),
.B(n_523),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_496),
.B(n_456),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_511),
.B(n_522),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_485),
.C(n_484),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_512),
.B(n_519),
.Y(n_531)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

XNOR2x1_ASAP7_75t_L g530 ( 
.A(n_517),
.B(n_518),
.Y(n_530)
);

XNOR2x1_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_470),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_473),
.C(n_470),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_491),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_521),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_473),
.C(n_464),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_472),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_495),
.B(n_454),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_524),
.B(n_450),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_501),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_525),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_527),
.B(n_538),
.Y(n_542)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_529),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_512),
.C(n_519),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_510),
.C(n_490),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_514),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_517),
.B(n_507),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_540),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_513),
.A2(n_498),
.B(n_492),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_435),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g545 ( 
.A(n_539),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_513),
.A2(n_481),
.B1(n_477),
.B2(n_445),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_544),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_523),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_548),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_508),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_534),
.B(n_508),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_549),
.B(n_451),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_528),
.A2(n_464),
.B1(n_455),
.B2(n_445),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_550),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_536),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_555),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_542),
.A2(n_532),
.B(n_531),
.Y(n_553)
);

AOI21x1_ASAP7_75t_L g561 ( 
.A1(n_553),
.A2(n_554),
.B(n_547),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_546),
.A2(n_535),
.B(n_446),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_552),
.B(n_541),
.C(n_543),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_558),
.A2(n_560),
.B(n_556),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_544),
.C(n_547),
.Y(n_560)
);

AOI31xp67_ASAP7_75t_L g563 ( 
.A1(n_561),
.A2(n_530),
.A3(n_550),
.B(n_459),
.Y(n_563)
);

AOI322xp5_ASAP7_75t_L g564 ( 
.A1(n_562),
.A2(n_563),
.A3(n_559),
.B1(n_530),
.B2(n_459),
.C1(n_537),
.C2(n_518),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_564),
.A2(n_499),
.B(n_537),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_565),
.B(n_499),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_566),
.B(n_459),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_440),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_568),
.A2(n_13),
.B(n_553),
.Y(n_569)
);


endmodule