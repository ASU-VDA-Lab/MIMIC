module real_jpeg_5185_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_1),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_23),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_159),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_2),
.A2(n_89),
.B1(n_159),
.B2(n_336),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_2),
.A2(n_159),
.B1(n_358),
.B2(n_361),
.Y(n_357)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_22),
.B1(n_86),
.B2(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_4),
.A2(n_22),
.B1(n_126),
.B2(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_27),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_22),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_4),
.A2(n_324),
.B(n_326),
.C(n_330),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_4),
.B(n_348),
.C(n_350),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_4),
.B(n_142),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_4),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_4),
.B(n_74),
.Y(n_387)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_6),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_6),
.Y(n_375)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_6),
.Y(n_383)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_7),
.Y(n_178)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_9),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_10),
.Y(n_179)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_11),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_12),
.A2(n_43),
.B1(n_118),
.B2(n_121),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_12),
.A2(n_43),
.B1(n_192),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_12),
.A2(n_43),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_134),
.B1(n_138),
.B2(n_140),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_13),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_140),
.B1(n_187),
.B2(n_191),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_13),
.A2(n_140),
.B1(n_251),
.B2(n_255),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_13),
.A2(n_140),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_450),
.B(n_453),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_148),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_57),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_19),
.B(n_58),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_20),
.B(n_235),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_21),
.B(n_46),
.Y(n_156)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_21),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_22),
.A2(n_327),
.B(n_329),
.Y(n_326)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_24),
.Y(n_180)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_27),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_27),
.B(n_40),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_27),
.B(n_158),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_31),
.Y(n_182)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_33),
.Y(n_176)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_36),
.Y(n_167)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_39),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_39),
.B(n_157),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_46),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_46),
.B(n_158),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_52),
.B2(n_55),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_51),
.Y(n_184)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_141),
.C(n_144),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_59),
.B(n_446),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_92),
.C(n_130),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_60),
.A2(n_162),
.B1(n_170),
.B2(n_171),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_60),
.B(n_155),
.C(n_162),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_60),
.B(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_60),
.A2(n_92),
.B1(n_170),
.B2(n_438),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_83),
.B(n_84),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_61),
.A2(n_225),
.B(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_62),
.B(n_85),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_62),
.B(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_62),
.B(n_335),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_74),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_66),
.Y(n_230)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_66),
.Y(n_256)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_66),
.Y(n_338)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_73),
.Y(n_254)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_74),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_74),
.B(n_335),
.Y(n_352)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_78),
.Y(n_361)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_82),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_82),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_83),
.A2(n_250),
.B(n_257),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_83),
.B(n_84),
.Y(n_305)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_88),
.Y(n_227)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_88),
.Y(n_346)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_92),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_123),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_93),
.A2(n_142),
.B(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_116),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_109),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_103),
.B2(n_105),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_99),
.Y(n_328)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_102),
.Y(n_300)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_115),
.Y(n_325)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_117),
.B(n_142),
.Y(n_205)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_122),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_125),
.B(n_143),
.Y(n_274)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_130),
.A2(n_131),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_132),
.A2(n_145),
.B(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_141),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_141),
.A2(n_144),
.B1(n_262),
.B2(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_143),
.B(n_165),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_143),
.A2(n_298),
.B(n_427),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_144),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_146),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_146),
.B(n_156),
.Y(n_423)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_416),
.B(n_441),
.C(n_444),
.D(n_449),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_408),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_264),
.C(n_313),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_238),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_218),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_153),
.B(n_218),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_172),
.C(n_203),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_154),
.B(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_164),
.B(n_274),
.Y(n_397)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_170),
.B(n_423),
.C(n_426),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_172),
.A2(n_173),
.B1(n_203),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_174),
.B(n_185),
.Y(n_232)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_177),
.A3(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_194),
.B(n_196),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_217),
.B(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_197),
.A2(n_211),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_197),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_201),
.Y(n_217)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_204),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_274),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_205),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_209),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_210),
.B(n_373),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_214),
.Y(n_360)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_217),
.B(n_356),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_218),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_218),
.B(n_239),
.Y(n_412)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.CI(n_231),
.CON(n_218),
.SN(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_223),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_224),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_225),
.B(n_334),
.Y(n_363)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_234),
.C(n_236),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_238),
.A2(n_411),
.B(n_412),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_240),
.B(n_242),
.C(n_258),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_258),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_244),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_248),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_257),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_257),
.B(n_352),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_261),
.C(n_262),
.Y(n_283)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_309),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_265),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_284),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_266),
.B(n_284),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_275),
.C(n_283),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_275),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_272),
.C(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_275)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_282),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_276),
.A2(n_282),
.B1(n_323),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_282),
.A2(n_288),
.B(n_293),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_308),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_295),
.B2(n_296),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_287),
.B(n_295),
.C(n_308),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_304),
.B(n_307),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_304),
.Y(n_307)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_307),
.A2(n_420),
.B1(n_421),
.B2(n_428),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_307),
.Y(n_428)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_309),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_310),
.B(n_312),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_339),
.B(n_407),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_315),
.B(n_318),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.C(n_331),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_322),
.A2(n_331),
.B1(n_332),
.B2(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_401),
.B(n_406),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_391),
.B(n_400),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_367),
.B(n_390),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_353),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_353),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_351),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_344),
.A2(n_345),
.B1(n_351),
.B2(n_370),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_362),
.Y(n_353)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_363),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_364),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_365),
.C(n_393),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_376),
.B(n_389),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_371),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_385),
.B(n_388),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_384),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_387),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_394),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_397),
.C(n_398),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_405),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_402),
.B(n_405),
.Y(n_406)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_410),
.B(n_413),
.C(n_414),
.D(n_415),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_431),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_430),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_430),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_429),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_428),
.C(n_429),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_422),
.A2(n_423),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_434),
.C(n_439),
.Y(n_448)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_431),
.A2(n_442),
.B(n_443),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_440),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_440),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_439),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_448),
.Y(n_449)
);

BUFx4f_ASAP7_75t_SL g450 ( 
.A(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

INVx13_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);


endmodule