module real_aes_4778_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g326 ( .A(n_0), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_1), .A2(n_15), .B1(n_220), .B2(n_223), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_2), .A2(n_20), .B1(n_118), .B2(n_125), .Y(n_117) );
INVx2_ASAP7_75t_L g286 ( .A(n_3), .Y(n_286) );
INVx1_ASAP7_75t_SL g351 ( .A(n_4), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_5), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_6), .B(n_337), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_7), .A2(n_49), .B1(n_142), .B2(n_145), .Y(n_141) );
XOR2xp5_ASAP7_75t_L g635 ( .A(n_8), .B(n_81), .Y(n_635) );
INVx1_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVxp67_ASAP7_75t_L g153 ( .A(n_9), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_9), .B(n_56), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_10), .A2(n_44), .B1(n_332), .B2(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_11), .B(n_161), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g84 ( .A1(n_12), .A2(n_36), .B1(n_85), .B2(n_107), .Y(n_84) );
NAND2xp5_ASAP7_75t_SL g100 ( .A(n_13), .B(n_89), .Y(n_100) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_14), .A2(n_54), .B(n_236), .Y(n_235) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_14), .A2(n_54), .B(n_236), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_16), .B(n_221), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_17), .A2(n_63), .B1(n_277), .B2(n_279), .Y(n_276) );
INVx2_ASAP7_75t_L g268 ( .A(n_18), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_19), .A2(n_53), .B1(n_131), .B2(n_136), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_21), .A2(n_26), .B1(n_227), .B2(n_229), .Y(n_226) );
AOI21xp33_ASAP7_75t_L g164 ( .A1(n_22), .A2(n_165), .B(n_167), .Y(n_164) );
BUFx3_ASAP7_75t_L g195 ( .A(n_23), .Y(n_195) );
O2A1O1Ixp5_ASAP7_75t_L g260 ( .A1(n_24), .A2(n_224), .B(n_261), .C(n_265), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_25), .A2(n_50), .B1(n_262), .B2(n_282), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_27), .Y(n_374) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_29), .A2(n_64), .B1(n_340), .B2(n_343), .Y(n_339) );
INVx1_ASAP7_75t_L g254 ( .A(n_30), .Y(n_254) );
INVx1_ASAP7_75t_L g90 ( .A(n_31), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_31), .B(n_55), .Y(n_150) );
INVx1_ASAP7_75t_L g168 ( .A(n_32), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_33), .B(n_250), .Y(n_321) );
INVx2_ASAP7_75t_L g266 ( .A(n_34), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_35), .Y(n_375) );
INVx2_ASAP7_75t_L g296 ( .A(n_37), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_38), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g354 ( .A(n_39), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_40), .A2(n_59), .B1(n_155), .B2(n_158), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_41), .Y(n_188) );
INVx1_ASAP7_75t_L g369 ( .A(n_42), .Y(n_369) );
INVx1_ASAP7_75t_L g236 ( .A(n_43), .Y(n_236) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_45), .Y(n_206) );
AND2x4_ASAP7_75t_L g238 ( .A(n_45), .B(n_204), .Y(n_238) );
AND2x4_ASAP7_75t_L g258 ( .A(n_45), .B(n_204), .Y(n_258) );
INVx1_ASAP7_75t_L g358 ( .A(n_46), .Y(n_358) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_47), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_48), .A2(n_60), .B1(n_128), .B2(n_129), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_51), .B(n_302), .Y(n_301) );
OA22x2_ASAP7_75t_L g94 ( .A1(n_52), .A2(n_56), .B1(n_89), .B2(n_93), .Y(n_94) );
INVx1_ASAP7_75t_L g114 ( .A(n_52), .Y(n_114) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_55), .B(n_112), .Y(n_177) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_55), .Y(n_198) );
OAI21xp33_ASAP7_75t_L g115 ( .A1(n_56), .A2(n_62), .B(n_116), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_57), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_58), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_61), .B(n_230), .Y(n_356) );
INVx1_ASAP7_75t_L g92 ( .A(n_62), .Y(n_92) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_62), .B(n_75), .Y(n_175) );
INVx1_ASAP7_75t_L g182 ( .A(n_64), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_65), .Y(n_183) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_66), .Y(n_222) );
BUFx5_ASAP7_75t_L g228 ( .A(n_66), .Y(n_228) );
INVx1_ASAP7_75t_L g264 ( .A(n_66), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_67), .B(n_302), .Y(n_352) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_67), .Y(n_643) );
INVx2_ASAP7_75t_L g299 ( .A(n_68), .Y(n_299) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_69), .Y(n_187) );
INVx1_ASAP7_75t_L g306 ( .A(n_70), .Y(n_306) );
INVx2_ASAP7_75t_L g377 ( .A(n_71), .Y(n_377) );
INVx2_ASAP7_75t_SL g204 ( .A(n_72), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_73), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_74), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g98 ( .A(n_75), .B(n_99), .Y(n_98) );
AO32x2_ASAP7_75t_L g217 ( .A1(n_76), .A2(n_218), .A3(n_233), .B1(n_237), .B2(n_239), .Y(n_217) );
AO22x2_ASAP7_75t_L g382 ( .A1(n_76), .A2(n_218), .B1(n_383), .B2(n_385), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_190), .B1(n_207), .B2(n_623), .C(n_630), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_180), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_178), .B2(n_179), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_80), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_81), .Y(n_179) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_140), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_117), .C(n_127), .D(n_130), .Y(n_83) );
AND2x4_ASAP7_75t_L g85 ( .A(n_86), .B(n_95), .Y(n_85) );
AND2x4_ASAP7_75t_L g128 ( .A(n_86), .B(n_123), .Y(n_128) );
AND2x2_ASAP7_75t_L g157 ( .A(n_86), .B(n_134), .Y(n_157) );
AND2x2_ASAP7_75t_L g163 ( .A(n_86), .B(n_138), .Y(n_163) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_94), .Y(n_86) );
INVx1_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
NAND2xp33_ASAP7_75t_L g88 ( .A(n_89), .B(n_90), .Y(n_88) );
INVx2_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx3_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g105 ( .A(n_89), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g116 ( .A(n_89), .Y(n_116) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_90), .B(n_114), .Y(n_113) );
INVxp67_ASAP7_75t_L g199 ( .A(n_90), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g91 ( .A(n_92), .B(n_93), .Y(n_91) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_92), .A2(n_116), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g122 ( .A(n_94), .Y(n_122) );
AND2x2_ASAP7_75t_L g144 ( .A(n_94), .B(n_121), .Y(n_144) );
AND2x2_ASAP7_75t_L g151 ( .A(n_94), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g109 ( .A(n_95), .B(n_110), .Y(n_109) );
AND2x4_ASAP7_75t_L g126 ( .A(n_95), .B(n_120), .Y(n_126) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_101), .Y(n_96) );
AND2x4_ASAP7_75t_L g123 ( .A(n_97), .B(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g134 ( .A(n_97), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
AND2x2_ASAP7_75t_L g147 ( .A(n_97), .B(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_99), .B(n_104), .Y(n_103) );
INVxp67_ASAP7_75t_L g112 ( .A(n_99), .Y(n_112) );
NAND3xp33_ASAP7_75t_L g176 ( .A(n_100), .B(n_111), .C(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx6_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g129 ( .A(n_110), .B(n_123), .Y(n_129) );
AND2x4_ASAP7_75t_L g159 ( .A(n_110), .B(n_138), .Y(n_159) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_114), .Y(n_200) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
AND2x4_ASAP7_75t_L g133 ( .A(n_120), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g137 ( .A(n_120), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g143 ( .A(n_134), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g138 ( .A(n_135), .B(n_139), .Y(n_138) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g166 ( .A(n_138), .B(n_144), .Y(n_166) );
NAND4xp25_ASAP7_75t_L g140 ( .A(n_141), .B(n_154), .C(n_160), .D(n_164), .Y(n_140) );
BUFx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx4f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_176), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_179), .B(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B1(n_185), .B2(n_189), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_181), .Y(n_189) );
XNOR2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
XOR2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
CKINVDCx14_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
BUFx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g634 ( .A(n_194), .B(n_201), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .C(n_200), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_205), .Y(n_201) );
OR2x2_ASAP7_75t_L g637 ( .A(n_202), .B(n_206), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_202), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_202), .B(n_205), .Y(n_641) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_528), .Y(n_210) );
NAND4xp25_ASAP7_75t_L g211 ( .A(n_212), .B(n_424), .C(n_471), .D(n_503), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_408), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_378), .Y(n_213) );
OAI21xp33_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_287), .B(n_309), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_242), .Y(n_215) );
INVx1_ASAP7_75t_L g423 ( .A(n_216), .Y(n_423) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_216), .B(n_291), .Y(n_428) );
AND2x2_ASAP7_75t_L g507 ( .A(n_216), .B(n_401), .Y(n_507) );
OR2x2_ASAP7_75t_L g531 ( .A(n_216), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g549 ( .A(n_216), .B(n_431), .Y(n_549) );
AND2x2_ASAP7_75t_L g571 ( .A(n_216), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g587 ( .A(n_216), .Y(n_587) );
BUFx8_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g455 ( .A(n_217), .Y(n_455) );
AND2x2_ASAP7_75t_L g603 ( .A(n_217), .B(n_454), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_224), .B1(n_226), .B2(n_231), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_220), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g248 ( .A(n_221), .Y(n_248) );
INVx1_ASAP7_75t_L g282 ( .A(n_221), .Y(n_282) );
INVx2_ASAP7_75t_L g327 ( .A(n_221), .Y(n_327) );
INVx6_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g223 ( .A(n_222), .Y(n_223) );
INVx3_ASAP7_75t_L g230 ( .A(n_222), .Y(n_230) );
INVx2_ASAP7_75t_L g342 ( .A(n_222), .Y(n_342) );
INVx2_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_223), .Y(n_343) );
INVx1_ASAP7_75t_L g628 ( .A(n_223), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_224), .A2(n_316), .B(n_318), .Y(n_315) );
INVx4_ASAP7_75t_L g372 ( .A(n_224), .Y(n_372) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_225), .Y(n_232) );
INVx4_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
INVx3_ASAP7_75t_L g284 ( .A(n_225), .Y(n_284) );
INVx1_ASAP7_75t_L g345 ( .A(n_225), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_227), .A2(n_327), .B1(n_374), .B2(n_375), .Y(n_373) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g319 ( .A(n_228), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_228), .Y(n_323) );
INVx2_ASAP7_75t_L g332 ( .A(n_228), .Y(n_332) );
INVx2_ASAP7_75t_L g355 ( .A(n_228), .Y(n_355) );
INVx1_ASAP7_75t_L g350 ( .A(n_229), .Y(n_350) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx2_ASAP7_75t_L g279 ( .A(n_230), .Y(n_279) );
INVx1_ASAP7_75t_L g317 ( .A(n_230), .Y(n_317) );
INVx1_ASAP7_75t_L g333 ( .A(n_230), .Y(n_333) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g280 ( .A(n_232), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_232), .A2(n_299), .B(n_300), .C(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_232), .B(n_335), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_232), .A2(n_350), .B(n_351), .C(n_352), .Y(n_349) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_233), .A2(n_245), .A3(n_259), .B(n_267), .Y(n_244) );
INVx2_ASAP7_75t_L g385 ( .A(n_233), .Y(n_385) );
BUFx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_234), .B(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_234), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g313 ( .A(n_234), .Y(n_313) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
BUFx3_ASAP7_75t_L g396 ( .A(n_235), .Y(n_396) );
AND2x2_ASAP7_75t_L g624 ( .A(n_237), .B(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g271 ( .A(n_238), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
AND2x2_ASAP7_75t_L g383 ( .A(n_238), .B(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g360 ( .A(n_239), .Y(n_360) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_240), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_241), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_241), .B(n_304), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_241), .B(n_304), .Y(n_335) );
BUFx3_ASAP7_75t_L g337 ( .A(n_241), .Y(n_337) );
INVx1_ASAP7_75t_L g384 ( .A(n_241), .Y(n_384) );
AND2x2_ASAP7_75t_L g511 ( .A(n_242), .B(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g592 ( .A(n_242), .B(n_448), .Y(n_592) );
INVxp67_ASAP7_75t_SL g608 ( .A(n_242), .Y(n_608) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_269), .Y(n_242) );
INVx1_ASAP7_75t_L g468 ( .A(n_243), .Y(n_468) );
INVx2_ASAP7_75t_SL g565 ( .A(n_243), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_243), .B(n_455), .Y(n_578) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g308 ( .A(n_244), .Y(n_308) );
OR2x2_ASAP7_75t_L g388 ( .A(n_244), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g401 ( .A(n_244), .B(n_292), .Y(n_401) );
AND2x2_ASAP7_75t_L g431 ( .A(n_244), .B(n_386), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_244), .B(n_389), .Y(n_484) );
AOI221x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_249), .B1(n_253), .B2(n_255), .C(n_257), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
AND2x2_ASAP7_75t_L g253 ( .A(n_250), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_251), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_257), .B(n_283), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g368 ( .A(n_257), .B(n_283), .C(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_257), .B(n_372), .Y(n_371) );
INVx4_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_269), .Y(n_414) );
INVx2_ASAP7_75t_L g447 ( .A(n_269), .Y(n_447) );
AND2x2_ASAP7_75t_L g614 ( .A(n_269), .B(n_386), .Y(n_614) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g290 ( .A(n_270), .Y(n_290) );
INVx1_ASAP7_75t_L g389 ( .A(n_270), .Y(n_389) );
AOI21x1_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_275), .B(n_285), .Y(n_270) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_273), .B(n_304), .Y(n_348) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B1(n_281), .B2(n_283), .Y(n_275) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g300 ( .A(n_278), .Y(n_300) );
INVx1_ASAP7_75t_L g295 ( .A(n_282), .Y(n_295) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_284), .A2(n_295), .B(n_296), .C(n_297), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_284), .A2(n_354), .B(n_355), .C(n_356), .Y(n_353) );
INVx2_ASAP7_75t_L g536 ( .A(n_287), .Y(n_536) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
NAND2x1p5_ASAP7_75t_L g400 ( .A(n_288), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_288), .B(n_381), .Y(n_486) );
INVx4_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_SL g426 ( .A(n_289), .Y(n_426) );
AND2x2_ASAP7_75t_L g545 ( .A(n_289), .B(n_431), .Y(n_545) );
AND2x2_ASAP7_75t_L g558 ( .A(n_289), .B(n_291), .Y(n_558) );
INVx2_ASAP7_75t_L g561 ( .A(n_289), .Y(n_561) );
BUFx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g454 ( .A(n_290), .Y(n_454) );
INVx2_ASAP7_75t_L g532 ( .A(n_291), .Y(n_532) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_308), .Y(n_291) );
INVx2_ASAP7_75t_L g386 ( .A(n_292), .Y(n_386) );
INVx1_ASAP7_75t_L g449 ( .A(n_292), .Y(n_449) );
BUFx3_ASAP7_75t_L g467 ( .A(n_292), .Y(n_467) );
AND2x4_ASAP7_75t_L g512 ( .A(n_292), .B(n_455), .Y(n_512) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_298), .A3(n_303), .B(n_305), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_300), .B(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NOR2xp33_ASAP7_75t_SL g357 ( .A(n_307), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_346), .Y(n_309) );
AND2x2_ASAP7_75t_L g574 ( .A(n_310), .B(n_406), .Y(n_574) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_329), .Y(n_310) );
INVx2_ASAP7_75t_L g398 ( .A(n_311), .Y(n_398) );
INVx1_ASAP7_75t_L g421 ( .A(n_311), .Y(n_421) );
AND2x2_ASAP7_75t_L g437 ( .A(n_311), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g500 ( .A(n_311), .Y(n_500) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_311), .Y(n_611) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_320), .B(n_328), .Y(n_314) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_L g397 ( .A(n_329), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g417 ( .A(n_329), .Y(n_417) );
INVx2_ASAP7_75t_L g435 ( .A(n_329), .Y(n_435) );
INVx1_ASAP7_75t_L g459 ( .A(n_329), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_330), .B(n_338), .Y(n_329) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_330), .B(n_338), .Y(n_405) );
OA21x2_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B(n_336), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_335), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
INVx1_ASAP7_75t_L g485 ( .A(n_346), .Y(n_485) );
AND2x2_ASAP7_75t_L g534 ( .A(n_346), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g622 ( .A(n_346), .B(n_397), .Y(n_622) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_359), .Y(n_346) );
OR2x2_ASAP7_75t_L g393 ( .A(n_347), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g407 ( .A(n_347), .Y(n_407) );
INVx2_ASAP7_75t_L g438 ( .A(n_347), .Y(n_438) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_347), .Y(n_464) );
INVx1_ASAP7_75t_L g498 ( .A(n_347), .Y(n_498) );
INVx1_ASAP7_75t_L g544 ( .A(n_347), .Y(n_544) );
AO31x2_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .A3(n_353), .B(n_357), .Y(n_347) );
INVx1_ASAP7_75t_L g632 ( .A(n_354), .Y(n_632) );
OR2x2_ASAP7_75t_L g443 ( .A(n_359), .B(n_398), .Y(n_443) );
AND2x2_ASAP7_75t_L g499 ( .A(n_359), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g567 ( .A(n_359), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g590 ( .A(n_359), .B(n_435), .Y(n_590) );
AO21x2_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B(n_376), .Y(n_359) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_361), .A2(n_376), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_370), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B1(n_366), .B2(n_368), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_372), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_390), .B1(n_399), .B2(n_402), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_380), .B(n_387), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_380), .A2(n_520), .B1(n_585), .B2(n_588), .C(n_591), .Y(n_584) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g526 ( .A(n_381), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_381), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
INVx1_ASAP7_75t_L g450 ( .A(n_382), .Y(n_450) );
AND2x4_ASAP7_75t_L g478 ( .A(n_382), .B(n_467), .Y(n_478) );
AND2x2_ASAP7_75t_L g502 ( .A(n_387), .B(n_466), .Y(n_502) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g527 ( .A(n_388), .Y(n_527) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_389), .Y(n_479) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp67_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g493 ( .A(n_393), .B(n_458), .Y(n_493) );
AND2x2_ASAP7_75t_L g406 ( .A(n_394), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g436 ( .A(n_394), .Y(n_436) );
BUFx2_ASAP7_75t_L g470 ( .A(n_394), .Y(n_470) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g514 ( .A(n_397), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_397), .B(n_470), .Y(n_524) );
AND2x2_ASAP7_75t_L g575 ( .A(n_397), .B(n_469), .Y(n_575) );
AND2x2_ASAP7_75t_L g598 ( .A(n_397), .B(n_488), .Y(n_598) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g410 ( .A(n_401), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g452 ( .A(n_401), .Y(n_452) );
INVx2_ASAP7_75t_L g518 ( .A(n_401), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_402), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_591) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_404), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g543 ( .A(n_405), .B(n_421), .Y(n_543) );
INVx2_ASAP7_75t_L g568 ( .A(n_405), .Y(n_568) );
AND2x2_ASAP7_75t_L g601 ( .A(n_405), .B(n_421), .Y(n_601) );
AND2x4_ASAP7_75t_L g413 ( .A(n_406), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g540 ( .A(n_406), .Y(n_540) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_407), .Y(n_442) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_407), .Y(n_547) );
OAI32xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .A3(n_415), .B1(n_418), .B2(n_422), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_409), .A2(n_618), .B1(n_619), .B2(n_621), .Y(n_617) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_413), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g517 ( .A(n_414), .Y(n_517) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI311xp33_ASAP7_75t_L g503 ( .A1(n_416), .A2(n_504), .A3(n_505), .B(n_508), .C(n_519), .Y(n_503) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g496 ( .A(n_417), .B(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND5xp2_ASAP7_75t_L g462 ( .A(n_420), .B(n_463), .C(n_465), .D(n_468), .E(n_469), .Y(n_462) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_439), .C(n_461), .Y(n_424) );
AOI31xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .A3(n_429), .B(n_432), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g586 ( .A(n_431), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g602 ( .A(n_431), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g620 ( .A(n_431), .B(n_447), .Y(n_620) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_437), .Y(n_433) );
AND2x4_ASAP7_75t_L g609 ( .A(n_434), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_435), .Y(n_522) );
BUFx2_ASAP7_75t_L g535 ( .A(n_435), .Y(n_535) );
AND2x4_ASAP7_75t_L g488 ( .A(n_436), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g548 ( .A(n_436), .B(n_500), .Y(n_548) );
AND2x2_ASAP7_75t_L g589 ( .A(n_437), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g595 ( .A(n_437), .B(n_459), .Y(n_595) );
INVx1_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_444), .B1(n_451), .B2(n_456), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g475 ( .A(n_441), .Y(n_475) );
OAI322xp33_ASAP7_75t_L g480 ( .A1(n_441), .A2(n_481), .A3(n_482), .B1(n_485), .B2(n_486), .C1(n_487), .C2(n_490), .Y(n_480) );
OR2x6_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVxp67_ASAP7_75t_L g460 ( .A(n_443), .Y(n_460) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_443), .Y(n_523) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g506 ( .A(n_447), .Y(n_506) );
AND2x2_ASAP7_75t_L g593 ( .A(n_447), .B(n_466), .Y(n_593) );
INVx1_ASAP7_75t_L g481 ( .A(n_448), .Y(n_481) );
AND2x4_ASAP7_75t_SL g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g491 ( .A(n_453), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x2_ASAP7_75t_L g564 ( .A(n_455), .B(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
AND2x2_ASAP7_75t_L g463 ( .A(n_458), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g474 ( .A(n_458), .Y(n_474) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_466), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI211xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_476), .B(n_480), .C(n_492), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OR2x2_ASAP7_75t_L g605 ( .A(n_479), .B(n_578), .Y(n_605) );
OAI211xp5_ASAP7_75t_L g596 ( .A1(n_481), .A2(n_597), .B(n_599), .C(n_606), .Y(n_596) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g572 ( .A(n_484), .Y(n_572) );
INVx1_ASAP7_75t_L g504 ( .A(n_488), .Y(n_504) );
AND2x2_ASAP7_75t_L g554 ( .A(n_488), .B(n_535), .Y(n_554) );
AND2x4_ASAP7_75t_L g581 ( .A(n_488), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g600 ( .A(n_488), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_501), .Y(n_492) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
INVxp67_ASAP7_75t_L g515 ( .A(n_497), .Y(n_515) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_497), .Y(n_557) );
AND2x2_ASAP7_75t_L g616 ( .A(n_497), .B(n_611), .Y(n_616) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g509 ( .A(n_499), .Y(n_509) );
AND2x2_ASAP7_75t_L g552 ( .A(n_500), .B(n_544), .Y(n_552) );
INVx1_ASAP7_75t_L g582 ( .A(n_500), .Y(n_582) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B1(n_513), .B2(n_516), .Y(n_508) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_524), .B(n_525), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g580 ( .A(n_522), .Y(n_580) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_583), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_550), .C(n_569), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_533), .B1(n_536), .B2(n_537), .C(n_541), .Y(n_530) );
OAI211xp5_ASAP7_75t_L g550 ( .A1(n_531), .A2(n_551), .B(n_553), .C(n_559), .Y(n_550) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g539 ( .A(n_535), .Y(n_539) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
NOR2x1p5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B1(n_546), .B2(n_549), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_543), .B(n_557), .Y(n_556) );
NOR2xp67_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g566 ( .A(n_552), .B(n_567), .Y(n_566) );
OAI21xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_558), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_562), .B(n_566), .Y(n_559) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_563), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI22xp33_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_573), .B1(n_576), .B2(n_579), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_575), .A2(n_600), .B1(n_602), .B2(n_604), .Y(n_599) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_596), .C(n_617), .Y(n_583) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g615 ( .A(n_590), .B(n_616), .Y(n_615) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g618 ( .A(n_600), .Y(n_618) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B1(n_612), .B2(n_615), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OA21x2_ASAP7_75t_L g639 ( .A1(n_625), .A2(n_640), .B(n_641), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
CKINVDCx16_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B1(n_635), .B2(n_636), .C1(n_638), .C2(n_642), .Y(n_630) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
endmodule