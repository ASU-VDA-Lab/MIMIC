module fake_jpeg_10278_n_63 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_10),
.B1(n_23),
.B2(n_22),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_9),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_8),
.B1(n_21),
.B2(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_2),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_44),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_47),
.B(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_5),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_49),
.Y(n_50)
);

FAx1_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_26),
.CI(n_11),
.CON(n_47),
.SN(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_4),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_12),
.B1(n_15),
.B2(n_17),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_6),
.B(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_53),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_58),
.Y(n_61)
);

OAI321xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_56),
.A3(n_55),
.B1(n_43),
.B2(n_50),
.C(n_42),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.C(n_24),
.Y(n_63)
);


endmodule