module fake_jpeg_15166_n_108 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_2),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_23),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_40),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_51),
.B1(n_47),
.B2(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_20),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_48),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_6),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_16),
.B1(n_22),
.B2(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_50),
.B(n_51),
.Y(n_71)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_63),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_16),
.B(n_22),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_37),
.B1(n_51),
.B2(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_3),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_68),
.C(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_8),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_77),
.B(n_55),
.C(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_68),
.C(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_81),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_41),
.B(n_11),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_87),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_53),
.B1(n_63),
.B2(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_88),
.B1(n_90),
.B2(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_61),
.C(n_53),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_53),
.B1(n_67),
.B2(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_71),
.B1(n_74),
.B2(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_78),
.B1(n_60),
.B2(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_78),
.B1(n_65),
.B2(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_102),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_90),
.C(n_83),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_91),
.C(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_10),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_100),
.B(n_11),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_103),
.B1(n_104),
.B2(n_12),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_12),
.Y(n_108)
);


endmodule