module real_jpeg_33543_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_0),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_0),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g333 ( 
.A1(n_1),
.A2(n_334),
.B1(n_336),
.B2(n_337),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_1),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_4),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_49),
.B1(n_76),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_49),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_5),
.B(n_176),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_5),
.A2(n_203),
.A3(n_205),
.B1(n_208),
.B2(n_214),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_5),
.B(n_53),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_5),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_192),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_6),
.Y(n_219)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_9),
.A2(n_302),
.B1(n_304),
.B2(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_9),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

INVx2_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

AOI22x1_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_72),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_11),
.A2(n_72),
.B1(n_152),
.B2(n_155),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_11),
.A2(n_72),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_320),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_293),
.B(n_318),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_226),
.B(n_292),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_184),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_18),
.B(n_184),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_19),
.B(n_126),
.C(n_168),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_90),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_50),
.B1(n_51),
.B2(n_89),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_21),
.B(n_51),
.C(n_92),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_42),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

NAND2x1p5_ASAP7_75t_L g200 ( 
.A(n_24),
.B(n_34),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_30),
.B2(n_32),
.Y(n_24)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_26),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_26),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_26),
.Y(n_261)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_33),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_34),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_34),
.B(n_194),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_36),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_39),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_40),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_40),
.Y(n_335)
);

AO22x2_ASAP7_75t_L g191 ( 
.A1(n_42),
.A2(n_192),
.B1(n_193),
.B2(n_199),
.Y(n_191)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_43),
.B(n_200),
.Y(n_233)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

OAI21x1_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_49),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_49),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_49),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_50),
.A2(n_51),
.B1(n_232),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_50),
.B(n_280),
.C(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_78),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_67),
.Y(n_52)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_53),
.Y(n_172)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_80),
.Y(n_79)
);

AOI22x1_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_65),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_67),
.B(n_79),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_73),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_79),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_85),
.Y(n_213)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g343 ( 
.A1(n_93),
.A2(n_344),
.B1(n_345),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_93),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_102),
.B(n_110),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g313 ( 
.A1(n_94),
.A2(n_102),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_117),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_111),
.Y(n_315)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_128),
.A3(n_133),
.B1(n_136),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_116),
.Y(n_314)
);

AOI22x1_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_168),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_143),
.B1(n_166),
.B2(n_167),
.Y(n_126)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_127),
.B(n_167),
.Y(n_317)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_143),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_143),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_143),
.B(n_273),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_151),
.B1(n_158),
.B2(n_161),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_154),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_167),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.C(n_177),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_170),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g312 ( 
.A1(n_169),
.A2(n_170),
.B1(n_313),
.B2(n_316),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_170),
.B(n_317),
.C(n_327),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B(n_173),
.Y(n_170)
);

AOI21x1_ASAP7_75t_L g345 ( 
.A1(n_171),
.A2(n_172),
.B(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_242),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_177),
.B(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_178),
.B(n_267),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_182),
.B(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_183),
.A2(n_301),
.B(n_308),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.C(n_201),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_185),
.A2(n_186),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_237),
.C(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_190),
.A2(n_201),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI22x1_ASAP7_75t_L g329 ( 
.A1(n_190),
.A2(n_286),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_238),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_201),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_220),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_220),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx4f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

OAI22x1_ASAP7_75t_L g331 ( 
.A1(n_222),
.A2(n_301),
.B1(n_332),
.B2(n_340),
.Y(n_331)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_283),
.B(n_291),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_239),
.B(n_282),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_236),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_232),
.B(n_300),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_232),
.B(n_300),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_276),
.B(n_281),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_265),
.B(n_275),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_249),
.B1(n_257),
.B2(n_262),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_272),
.B(n_274),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_279),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_289),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2x1_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_297),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_311),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_310),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_SL g323 ( 
.A(n_299),
.B(n_310),
.C(n_311),
.Y(n_323)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_303),
.Y(n_339)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_348),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_323),
.B(n_324),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_341),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);


endmodule