module real_aes_433_n_13 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_13);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_13;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
AOI322xp5_ASAP7_75t_SL g13 ( .A1(n_0), .A2(n_12), .A3(n_14), .B1(n_15), .B2(n_28), .C1(n_39), .C2(n_45), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_1), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_2), .B(n_5), .C(n_21), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_3), .Y(n_21) );
NAND3xp33_ASAP7_75t_SL g24 ( .A(n_4), .B(n_25), .C(n_26), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_4), .B(n_19), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_6), .Y(n_27) );
NOR2xp33_ASAP7_75t_R g38 ( .A(n_6), .B(n_8), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_7), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g36 ( .A(n_7), .B(n_37), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_9), .B(n_27), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_9), .Y(n_34) );
INVx3_ASAP7_75t_L g44 ( .A(n_10), .Y(n_44) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_11), .Y(n_23) );
NAND2xp33_ASAP7_75t_SL g48 ( .A(n_11), .B(n_18), .Y(n_48) );
NAND2xp33_ASAP7_75t_SL g46 ( .A(n_14), .B(n_47), .Y(n_46) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_17), .B(n_24), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g17 ( .A(n_18), .B(n_23), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g19 ( .A(n_20), .B(n_22), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g31 ( .A(n_23), .B(n_32), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g47 ( .A(n_24), .B(n_48), .Y(n_47) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_29), .Y(n_28) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_30), .B(n_33), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_31), .Y(n_30) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_34), .B(n_35), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
CKINVDCx14_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_41), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
INVx2_ASAP7_75t_L g42 ( .A(n_43), .Y(n_42) );
HB1xp67_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
INVx1_ASAP7_75t_SL g45 ( .A(n_46), .Y(n_45) );
endmodule