module fake_jpeg_13885_n_198 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_1),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_SL g76 ( 
.A(n_12),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_19),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_22),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_62),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_76),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_91),
.Y(n_97)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_92),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_107),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_103),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_78),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_69),
.B(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_82),
.B1(n_65),
.B2(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_59),
.B1(n_66),
.B2(n_82),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_114),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_83),
.B1(n_24),
.B2(n_25),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_93),
.B1(n_70),
.B2(n_71),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_131),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_133),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_94),
.B1(n_65),
.B2(n_59),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_139),
.B1(n_150),
.B2(n_27),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_66),
.B1(n_63),
.B2(n_73),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_113),
.CI(n_119),
.CON(n_142),
.SN(n_142)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_152),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_75),
.B(n_67),
.C(n_60),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_147),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_85),
.B1(n_64),
.B2(n_80),
.Y(n_145)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_10),
.B(n_11),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_83),
.C(n_80),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_17),
.C(n_21),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_9),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_156),
.B1(n_159),
.B2(n_164),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_145),
.B1(n_149),
.B2(n_34),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_9),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_145),
.B1(n_144),
.B2(n_149),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_136),
.C(n_137),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_171),
.C(n_178),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_164),
.B1(n_160),
.B2(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_184),
.B1(n_176),
.B2(n_173),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_164),
.B1(n_169),
.B2(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_28),
.B(n_33),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_181),
.A2(n_170),
.B1(n_177),
.B2(n_173),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_188),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_181),
.B1(n_182),
.B2(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_35),
.C(n_39),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_40),
.B(n_43),
.C(n_45),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_47),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_48),
.C(n_52),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_53),
.Y(n_198)
);


endmodule