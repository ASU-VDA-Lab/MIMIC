module fake_jpeg_26634_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_38),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_23),
.B(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_24),
.B1(n_28),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_54),
.B1(n_28),
.B2(n_21),
.Y(n_71)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_21),
.B2(n_16),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_62),
.Y(n_72)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_46),
.B(n_40),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_18),
.B(n_30),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_71),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_83),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_45),
.C(n_42),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_65),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_44),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_18),
.B1(n_27),
.B2(n_32),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_31),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_42),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_64),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_29),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_94),
.Y(n_108)
);

CKINVDCx9p33_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_43),
.B1(n_37),
.B2(n_20),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_25),
.B1(n_20),
.B2(n_58),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_37),
.B1(n_43),
.B2(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_145)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_103),
.Y(n_127)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_104),
.A2(n_118),
.B1(n_101),
.B2(n_32),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_53),
.B1(n_49),
.B2(n_25),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_86),
.C(n_70),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_53),
.B1(n_25),
.B2(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_125),
.Y(n_129)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_64),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_17),
.CI(n_33),
.CON(n_118),
.SN(n_118)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_45),
.Y(n_152)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_27),
.B1(n_19),
.B2(n_34),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_123),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_74),
.A2(n_19),
.B1(n_34),
.B2(n_17),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_86),
.Y(n_132)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_151),
.Y(n_169)
);

AO21x2_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_86),
.B(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_143),
.B1(n_121),
.B2(n_92),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_138),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_45),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_72),
.A3(n_84),
.B1(n_96),
.B2(n_88),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_118),
.B(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_89),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_139),
.B(n_142),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_144),
.Y(n_164)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_77),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_106),
.B1(n_124),
.B2(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_155),
.Y(n_180)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_26),
.CI(n_19),
.CON(n_185),
.SN(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_34),
.Y(n_155)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_91),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_162),
.B1(n_148),
.B2(n_141),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_130),
.B1(n_154),
.B2(n_131),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_160),
.A2(n_178),
.B1(n_189),
.B2(n_61),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_171),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_114),
.B(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_167),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_117),
.B(n_113),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_173),
.B(n_170),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_133),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_103),
.B1(n_75),
.B2(n_80),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_175),
.B1(n_179),
.B2(n_144),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_113),
.B(n_2),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_26),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_176),
.C(n_132),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_75),
.B1(n_97),
.B2(n_66),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_26),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_91),
.B1(n_77),
.B2(n_26),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_66),
.B1(n_50),
.B2(n_57),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_77),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_133),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_186),
.Y(n_207)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_57),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_150),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_135),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_180),
.Y(n_239)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_192),
.A2(n_196),
.B1(n_217),
.B2(n_206),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_203),
.B1(n_205),
.B2(n_214),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_129),
.B1(n_149),
.B2(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_137),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_209),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_141),
.B1(n_129),
.B2(n_138),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_162),
.A2(n_151),
.B1(n_156),
.B2(n_57),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_64),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_1),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_9),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_50),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_61),
.B1(n_64),
.B2(n_8),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_172),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_171),
.C(n_174),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_237),
.C(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_235),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_161),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_238),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_204),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_176),
.C(n_159),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_159),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_206),
.Y(n_261)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_211),
.B1(n_192),
.B2(n_218),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_254),
.B1(n_260),
.B2(n_262),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_181),
.B1(n_200),
.B2(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_226),
.C(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_267),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_215),
.C(n_216),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_259),
.C(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_180),
.C(n_206),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_175),
.B1(n_179),
.B2(n_187),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_264),
.Y(n_280)
);

AOI211xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_195),
.B(n_185),
.C(n_193),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_217),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_265),
.Y(n_272)
);

XNOR2x2_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_219),
.Y(n_266)
);

XOR2x2_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_220),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_223),
.B(n_6),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_232),
.A2(n_1),
.B(n_2),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_226),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_278),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_238),
.C(n_246),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_283),
.C(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_268),
.B(n_10),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_263),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_279),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_230),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_281),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_263),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_224),
.C(n_233),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_224),
.C(n_8),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_8),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_6),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_259),
.C(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_287),
.C(n_298),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_252),
.B1(n_253),
.B2(n_266),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_262),
.B1(n_251),
.B2(n_249),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_280),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_300),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_301),
.B(n_307),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_270),
.B(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_290),
.B(n_296),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_269),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_308),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_6),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_10),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_10),
.B(n_13),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_299),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_4),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_298),
.C(n_294),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_320),
.C(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_317),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_286),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_302),
.B(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_4),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_292),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_5),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_311),
.C(n_308),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_303),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_327),
.B1(n_322),
.B2(n_321),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_4),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_329),
.B1(n_12),
.B2(n_15),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_330),
.B1(n_324),
.B2(n_314),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_323),
.B(n_331),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_331),
.Y(n_337)
);

OAI21x1_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_12),
.B(n_1),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_3),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_3),
.C(n_333),
.Y(n_340)
);


endmodule