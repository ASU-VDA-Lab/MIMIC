module fake_jpeg_2799_n_221 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_33),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_34),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_24),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_86),
.Y(n_101)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx12f_ASAP7_75t_SL g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_0),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_72),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_56),
.C(n_57),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_88),
.C(n_64),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_102),
.C(n_66),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_65),
.B1(n_71),
.B2(n_74),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_85),
.B1(n_88),
.B2(n_82),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_79),
.B(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_59),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_70),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_108),
.B1(n_77),
.B2(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_104),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_65),
.B1(n_59),
.B2(n_74),
.Y(n_108)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_1),
.C(n_3),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_119),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_76),
.B(n_58),
.C(n_54),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_84),
.B1(n_87),
.B2(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_92),
.B(n_109),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_1),
.B(n_5),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_101),
.C(n_2),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_26),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_71),
.B1(n_59),
.B2(n_55),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_128),
.B1(n_134),
.B2(n_136),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_63),
.B1(n_87),
.B2(n_83),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_84),
.B1(n_90),
.B2(n_63),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_77),
.B1(n_55),
.B2(n_67),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_55),
.B1(n_75),
.B2(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_6),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_75),
.B1(n_3),
.B2(n_5),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_153)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_27),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_29),
.B(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_7),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_7),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_8),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_165),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_16),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_16),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_18),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_40),
.B1(n_51),
.B2(n_49),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_166),
.B(n_41),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_21),
.B(n_52),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_25),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_36),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_129),
.Y(n_173)
);

OAI322xp33_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_183),
.A3(n_188),
.B1(n_47),
.B2(n_48),
.C1(n_169),
.C2(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_157),
.C(n_147),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_189),
.C(n_171),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_141),
.B1(n_38),
.B2(n_39),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_186),
.B1(n_163),
.B2(n_189),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_42),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_43),
.C(n_44),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_45),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_162),
.B1(n_153),
.B2(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_193),
.B1(n_182),
.B2(n_190),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_187),
.C(n_184),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_182),
.B1(n_190),
.B2(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_194),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_199),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_198),
.B(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_205),
.B(n_206),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_204),
.C(n_208),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_216),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_201),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_201),
.Y(n_221)
);


endmodule