module fake_jpeg_2006_n_103 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_41),
.C(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_6),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_34),
.B1(n_42),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_62),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_31),
.B(n_33),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_63),
.B(n_0),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_29),
.B1(n_12),
.B2(n_13),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_53),
.B1(n_1),
.B2(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_3),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_67),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_70),
.B(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_86),
.B1(n_85),
.B2(n_76),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_20),
.B(n_10),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_22),
.B(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_7),
.B1(n_11),
.B2(n_15),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_91),
.C(n_92),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_83),
.Y(n_91)
);

AOI21x1_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_87),
.B(n_90),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_92),
.C(n_91),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_79),
.B(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_93),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_7),
.C(n_18),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_21),
.B(n_26),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_27),
.Y(n_103)
);


endmodule