module fake_jpeg_29019_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx8_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_3),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_6),
.B(n_0),
.C(n_1),
.Y(n_7)
);

MAJIxp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_8),
.C(n_1),
.Y(n_10)
);

XNOR2x1_ASAP7_75t_L g8 ( 
.A(n_6),
.B(n_0),
.Y(n_8)
);

BUFx24_ASAP7_75t_SL g9 ( 
.A(n_8),
.Y(n_9)
);

AOI322xp5_ASAP7_75t_L g11 ( 
.A1(n_9),
.A2(n_10),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_8),
.C2(n_7),
.Y(n_11)
);


endmodule