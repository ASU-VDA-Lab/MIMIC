module fake_jpeg_730_n_523 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_523);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_523;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_57),
.Y(n_156)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_58),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_60),
.Y(n_185)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_62),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_17),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_63),
.A2(n_69),
.B(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_17),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_84),
.Y(n_203)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_118),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_111),
.Y(n_126)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_32),
.B(n_18),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_107),
.Y(n_124)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_103),
.Y(n_208)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_110),
.B(n_116),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_15),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_50),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_50),
.Y(n_127)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_20),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_121),
.Y(n_148)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_20),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_127),
.A2(n_158),
.B(n_202),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_32),
.B1(n_48),
.B2(n_27),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_131),
.A2(n_141),
.B1(n_150),
.B2(n_170),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_63),
.B(n_22),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_132),
.B(n_147),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_59),
.A2(n_32),
.B1(n_27),
.B2(n_55),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_144),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_145),
.B(n_146),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_54),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_19),
.B1(n_51),
.B2(n_40),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_60),
.A2(n_27),
.B1(n_54),
.B2(n_36),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_91),
.B(n_51),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_64),
.B(n_40),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_164),
.A2(n_174),
.B(n_198),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_62),
.B(n_36),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_166),
.B(n_168),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_35),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_95),
.A2(n_43),
.B1(n_28),
.B2(n_35),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_28),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_26),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_187),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_72),
.A2(n_26),
.B1(n_22),
.B2(n_53),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_181),
.A2(n_83),
.B1(n_62),
.B2(n_32),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_78),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_79),
.A2(n_53),
.B1(n_31),
.B2(n_23),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_81),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_200),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_82),
.A2(n_53),
.B1(n_23),
.B2(n_3),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_196),
.B1(n_206),
.B2(n_4),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_86),
.A2(n_112),
.B1(n_94),
.B2(n_92),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_195),
.A2(n_197),
.B1(n_193),
.B2(n_156),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_88),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_90),
.A2(n_23),
.B1(n_2),
.B2(n_4),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_75),
.B(n_1),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_63),
.B(n_1),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_63),
.B(n_2),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_205),
.B(n_161),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_63),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_209),
.Y(n_320)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_211),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_212),
.A2(n_237),
.B1(n_280),
.B2(n_260),
.Y(n_310)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_213),
.Y(n_301)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_214),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_215),
.A2(n_223),
.B1(n_231),
.B2(n_233),
.Y(n_293)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_216),
.Y(n_309)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx4_ASAP7_75t_SL g315 ( 
.A(n_217),
.Y(n_315)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_218),
.Y(n_302)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

FAx1_ASAP7_75t_L g220 ( 
.A(n_139),
.B(n_6),
.CI(n_8),
.CON(n_220),
.SN(n_220)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_220),
.B(n_268),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_221),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_124),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_150),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_225),
.A2(n_227),
.B1(n_252),
.B2(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_141),
.A2(n_195),
.B1(n_131),
.B2(n_181),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_228),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_229),
.B(n_247),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_124),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_230),
.B(n_262),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_186),
.A2(n_143),
.B1(n_172),
.B2(n_159),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_186),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_139),
.B(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_235),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_126),
.A2(n_14),
.B1(n_15),
.B2(n_137),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_154),
.B(n_15),
.Y(n_239)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_182),
.B(n_138),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_267),
.Y(n_284)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_245),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_130),
.A2(n_142),
.B1(n_207),
.B2(n_169),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_246),
.A2(n_269),
.B(n_253),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_125),
.Y(n_249)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_250),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_170),
.A2(n_188),
.B1(n_197),
.B2(n_135),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_259),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_123),
.B(n_136),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_256),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_163),
.B1(n_201),
.B2(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_149),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g260 ( 
.A(n_140),
.Y(n_260)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_157),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_167),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_264),
.Y(n_328)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_173),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_175),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_265),
.Y(n_325)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_266),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_162),
.B(n_179),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_149),
.B(n_152),
.CI(n_162),
.CON(n_269),
.SN(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_152),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_130),
.B(n_178),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_203),
.A2(n_191),
.B1(n_178),
.B2(n_183),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_275),
.B1(n_277),
.B2(n_218),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_175),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_153),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_278),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_203),
.A2(n_185),
.B1(n_165),
.B2(n_204),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_171),
.B(n_185),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_274),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_163),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_312),
.C(n_262),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_291),
.A2(n_305),
.B1(n_307),
.B2(n_324),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_230),
.B(n_201),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_310),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_220),
.A2(n_201),
.B(n_240),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_217),
.B(n_238),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_240),
.A2(n_267),
.B1(n_220),
.B2(n_257),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_234),
.B1(n_250),
.B2(n_254),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_242),
.B(n_248),
.C(n_256),
.Y(n_312)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_239),
.B(n_251),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_232),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_322),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_212),
.A2(n_278),
.B1(n_237),
.B2(n_236),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_283),
.A2(n_236),
.B1(n_224),
.B2(n_246),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_332),
.A2(n_361),
.B1(n_366),
.B2(n_370),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_335),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_334),
.B(n_350),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_275),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_269),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_339),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_269),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_290),
.B(n_256),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_341),
.B(n_357),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_328),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_342),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_343),
.A2(n_348),
.B(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_300),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_303),
.B(n_316),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_285),
.B(n_235),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_351),
.B(n_329),
.Y(n_402)
);

AOI22x1_ASAP7_75t_L g353 ( 
.A1(n_283),
.A2(n_279),
.B1(n_268),
.B2(n_245),
.Y(n_353)
);

AO21x2_ASAP7_75t_SL g379 ( 
.A1(n_353),
.A2(n_368),
.B(n_302),
.Y(n_379)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_291),
.A2(n_324),
.B1(n_281),
.B2(n_303),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_355),
.A2(n_359),
.B1(n_363),
.B2(n_296),
.Y(n_392)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_216),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_281),
.A2(n_211),
.B1(n_264),
.B2(n_263),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_210),
.B(n_243),
.C(n_213),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_360),
.B(n_362),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_282),
.A2(n_228),
.B1(n_265),
.B2(n_266),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_282),
.B(n_209),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_287),
.A2(n_241),
.B1(n_292),
.B2(n_318),
.Y(n_363)
);

A2O1A1O1Ixp25_ASAP7_75t_L g364 ( 
.A1(n_298),
.A2(n_294),
.B(n_313),
.C(n_323),
.D(n_308),
.Y(n_364)
);

O2A1O1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_319),
.B(n_321),
.C(n_317),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_365),
.A2(n_301),
.B(n_327),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_293),
.A2(n_294),
.B1(n_298),
.B2(n_286),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_298),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_367),
.B(n_335),
.Y(n_393)
);

AO21x2_ASAP7_75t_L g368 ( 
.A1(n_306),
.A2(n_289),
.B(n_309),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_325),
.A2(n_286),
.B1(n_315),
.B2(n_299),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_355),
.A2(n_315),
.B1(n_330),
.B2(n_297),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_383),
.B1(n_392),
.B2(n_361),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_366),
.A2(n_301),
.B1(n_330),
.B2(n_331),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_391),
.B(n_399),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_379),
.A2(n_368),
.B1(n_353),
.B2(n_358),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_354),
.A2(n_304),
.B1(n_296),
.B2(n_329),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_359),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_369),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_334),
.B(n_302),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_386),
.B(n_396),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_345),
.A2(n_321),
.B1(n_327),
.B2(n_289),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_390),
.A2(n_385),
.B1(n_368),
.B2(n_373),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_339),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_343),
.A2(n_348),
.B(n_365),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_395),
.A2(n_337),
.B(n_338),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_356),
.B(n_309),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_397),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_352),
.A2(n_320),
.B(n_331),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_340),
.C(n_367),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_403),
.A2(n_379),
.B1(n_392),
.B2(n_382),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_351),
.C(n_363),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_409),
.C(n_418),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_408),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_407),
.A2(n_426),
.B(n_401),
.Y(n_433)
);

AO21x1_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_337),
.B(n_352),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_337),
.C(n_341),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_393),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_414),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_383),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_419),
.A2(n_422),
.B1(n_379),
.B2(n_390),
.Y(n_440)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_395),
.B(n_360),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_420),
.B(n_389),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_424),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_389),
.A2(n_332),
.B1(n_333),
.B2(n_342),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_375),
.C(n_394),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_428),
.C(n_409),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_381),
.B(n_357),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_387),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_429),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_391),
.A2(n_364),
.B(n_362),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_427),
.A2(n_379),
.B1(n_401),
.B2(n_372),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_353),
.C(n_370),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_434),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_382),
.B1(n_384),
.B2(n_373),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_436),
.B1(n_437),
.B2(n_440),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_384),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_377),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_443),
.C(n_409),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_452),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_403),
.A2(n_379),
.B1(n_377),
.B2(n_381),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_441),
.A2(n_444),
.B1(n_446),
.B2(n_414),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_399),
.C(n_397),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_379),
.B1(n_400),
.B2(n_374),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_413),
.A2(n_374),
.B1(n_371),
.B2(n_376),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_422),
.A2(n_371),
.B1(n_368),
.B2(n_380),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_423),
.B(n_388),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_451),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_459),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_461),
.C(n_466),
.Y(n_474)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_456),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_SL g458 ( 
.A(n_435),
.B(n_423),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_463),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_451),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_407),
.C(n_406),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_441),
.A2(n_405),
.B1(n_419),
.B2(n_412),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_462),
.A2(n_467),
.B1(n_431),
.B2(n_445),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_408),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_449),
.B(n_424),
.Y(n_464)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_464),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_398),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_426),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_434),
.C(n_439),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_437),
.A2(n_415),
.B1(n_420),
.B2(n_408),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_420),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_443),
.C(n_450),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_468),
.A2(n_447),
.B1(n_433),
.B2(n_436),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_477),
.B1(n_480),
.B2(n_484),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_476),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_460),
.A2(n_447),
.B1(n_444),
.B2(n_445),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_435),
.C(n_430),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_479),
.Y(n_494)
);

XOR2x2_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_449),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_462),
.A2(n_448),
.B1(n_446),
.B2(n_428),
.Y(n_480)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_482),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_468),
.A2(n_415),
.B1(n_427),
.B2(n_442),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_471),
.A2(n_470),
.B(n_467),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_487),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_455),
.C(n_457),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_457),
.C(n_463),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_490),
.B(n_491),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_472),
.B(n_464),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_458),
.C(n_453),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_493),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_481),
.A2(n_470),
.B(n_479),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_453),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_469),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_473),
.C(n_483),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_498),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_473),
.C(n_483),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_485),
.A2(n_484),
.B1(n_456),
.B2(n_486),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_489),
.Y(n_507)
);

NOR2x1_ASAP7_75t_SL g500 ( 
.A(n_492),
.B(n_482),
.Y(n_500)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_500),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_475),
.C(n_477),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_489),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_495),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_510),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_505),
.B(n_496),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_513),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_508),
.A2(n_499),
.B1(n_503),
.B2(n_480),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_514),
.A2(n_506),
.B(n_497),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_512),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_517),
.A2(n_518),
.B(n_501),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_512),
.C(n_507),
.Y(n_518)
);

AOI321xp33_ASAP7_75t_L g520 ( 
.A1(n_519),
.A2(n_498),
.A3(n_490),
.B1(n_442),
.B2(n_416),
.C(n_410),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_416),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_521),
.A2(n_410),
.B(n_417),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_417),
.B(n_411),
.Y(n_523)
);


endmodule