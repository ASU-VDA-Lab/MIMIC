module real_aes_13670_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_235;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_951;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_928;
wire n_155;
wire n_637;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_922;
wire n_679;
wire n_482;
wire n_520;
wire n_926;
wire n_633;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g567 ( .A(n_0), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g684 ( .A(n_1), .Y(n_684) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_2), .A2(n_48), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g193 ( .A(n_2), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_3), .B(n_251), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_4), .B(n_245), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_5), .B(n_170), .Y(n_169) );
NAND2xp33_ASAP7_75t_L g225 ( .A(n_6), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g633 ( .A(n_7), .B(n_231), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_7), .A2(n_97), .B1(n_948), .B2(n_949), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_7), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_8), .B(n_268), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_9), .B(n_206), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_10), .A2(n_66), .B1(n_922), .B2(n_923), .Y(n_921) );
INVx1_ASAP7_75t_L g923 ( .A(n_10), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_11), .B(n_173), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_12), .Y(n_190) );
INVx1_ASAP7_75t_L g158 ( .A(n_13), .Y(n_158) );
BUFx3_ASAP7_75t_L g162 ( .A(n_13), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_14), .B(n_230), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_15), .A2(n_297), .B(n_347), .C(n_349), .Y(n_346) );
BUFx10_ASAP7_75t_L g143 ( .A(n_16), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_17), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_18), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_19), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_20), .B(n_253), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_21), .A2(n_227), .B(n_338), .C(n_339), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_22), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_23), .B(n_291), .C(n_611), .Y(n_613) );
AND2x2_ASAP7_75t_L g241 ( .A(n_24), .B(n_240), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_25), .B(n_170), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_26), .B(n_230), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_27), .A2(n_75), .B1(n_207), .B2(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g185 ( .A(n_28), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_29), .A2(n_76), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_29), .Y(n_940) );
INVx1_ASAP7_75t_L g176 ( .A(n_30), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_31), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_32), .B(n_207), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_33), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g123 ( .A(n_34), .Y(n_123) );
AND3x2_ASAP7_75t_L g932 ( .A(n_34), .B(n_115), .C(n_141), .Y(n_932) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_35), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_36), .B(n_297), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_37), .B(n_230), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_38), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_39), .B(n_156), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_40), .Y(n_348) );
AND2x4_ASAP7_75t_L g184 ( .A(n_41), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_42), .B(n_230), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_43), .B(n_240), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_44), .B(n_230), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_45), .A2(n_88), .B1(n_206), .B2(n_207), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_46), .A2(n_919), .B1(n_925), .B2(n_926), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_46), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_47), .A2(n_920), .B1(n_921), .B2(n_924), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_47), .Y(n_924) );
INVx1_ASAP7_75t_L g192 ( .A(n_48), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_49), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_50), .A2(n_565), .B(n_566), .C(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g179 ( .A(n_51), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_52), .B(n_230), .Y(n_688) );
AND2x4_ASAP7_75t_L g120 ( .A(n_53), .B(n_121), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_54), .Y(n_929) );
INVx3_ASAP7_75t_L g651 ( .A(n_55), .Y(n_651) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_56), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g136 ( .A(n_56), .B(n_78), .Y(n_136) );
AND2x2_ASAP7_75t_L g284 ( .A(n_57), .B(n_231), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_58), .Y(n_957) );
INVx1_ASAP7_75t_L g121 ( .A(n_59), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_60), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_61), .B(n_578), .Y(n_583) );
NAND2x1_ASAP7_75t_L g296 ( .A(n_62), .B(n_297), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_63), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_64), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g663 ( .A(n_65), .Y(n_663) );
INVx1_ASAP7_75t_L g922 ( .A(n_66), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_67), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_68), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_70), .B(n_206), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_71), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_72), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_73), .B(n_291), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_74), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g941 ( .A(n_76), .Y(n_941) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_77), .B(n_276), .Y(n_283) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_79), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_80), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_81), .B(n_268), .Y(n_292) );
NAND2xp33_ASAP7_75t_SL g167 ( .A(n_82), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_83), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g558 ( .A(n_84), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_85), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_86), .B(n_160), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_87), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g165 ( .A(n_89), .Y(n_165) );
BUFx3_ASAP7_75t_L g173 ( .A(n_89), .Y(n_173) );
INVx1_ASAP7_75t_L g202 ( .A(n_89), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_90), .B(n_282), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_91), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_92), .B(n_206), .Y(n_682) );
INVx1_ASAP7_75t_L g649 ( .A(n_93), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_94), .B(n_266), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_95), .B(n_231), .Y(n_599) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_96), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g949 ( .A(n_97), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_98), .B(n_582), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_99), .Y(n_645) );
INVx1_ASAP7_75t_L g641 ( .A(n_100), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_101), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_102), .B(n_156), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_103), .B(n_578), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_124), .B(n_956), .Y(n_104) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx10_ASAP7_75t_R g958 ( .A(n_108), .Y(n_958) );
OR2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_114), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
AND2x2_ASAP7_75t_L g140 ( .A(n_115), .B(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g134 ( .A(n_116), .Y(n_134) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g544 ( .A(n_122), .Y(n_544) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_123), .B(n_136), .Y(n_135) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_933), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_137), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI21xp33_ASAP7_75t_L g950 ( .A1(n_127), .A2(n_937), .B(n_951), .Y(n_950) );
NOR2xp67_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx3_ASAP7_75t_L g955 ( .A(n_132), .Y(n_955) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_SL g945 ( .A(n_133), .Y(n_945) );
NOR2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_928), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_143), .B(n_932), .Y(n_931) );
CKINVDCx11_ASAP7_75t_R g934 ( .A(n_143), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_917), .B1(n_918), .B2(n_927), .Y(n_144) );
INVx2_ASAP7_75t_L g927 ( .A(n_145), .Y(n_927) );
AO22x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_541), .B1(n_542), .B2(n_545), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_146), .A2(n_938), .B1(n_939), .B2(n_942), .Y(n_937) );
INVx2_ASAP7_75t_L g942 ( .A(n_146), .Y(n_942) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_424), .Y(n_146) );
NOR4xp25_ASAP7_75t_L g147 ( .A(n_148), .B(n_324), .C(n_370), .D(n_410), .Y(n_147) );
OAI21xp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_233), .B(n_301), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_186), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_150), .B(n_401), .Y(n_444) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g504 ( .A(n_151), .B(n_401), .Y(n_504) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_152), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_152), .B(n_317), .Y(n_515) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g311 ( .A(n_153), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g315 ( .A(n_153), .Y(n_315) );
AND2x2_ASAP7_75t_L g386 ( .A(n_153), .B(n_213), .Y(n_386) );
AND2x2_ASAP7_75t_L g414 ( .A(n_153), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g438 ( .A(n_153), .B(n_353), .Y(n_438) );
AND2x2_ASAP7_75t_L g468 ( .A(n_153), .B(n_353), .Y(n_468) );
AO31x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_166), .A3(n_174), .B(n_180), .Y(n_153) );
AO21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_159), .B(n_163), .Y(n_154) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g168 ( .A(n_157), .Y(n_168) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
INVx2_ASAP7_75t_L g251 ( .A(n_157), .Y(n_251) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g247 ( .A(n_158), .Y(n_247) );
INVx2_ASAP7_75t_L g295 ( .A(n_160), .Y(n_295) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
INVx2_ASAP7_75t_L g218 ( .A(n_161), .Y(n_218) );
INVx2_ASAP7_75t_L g282 ( .A(n_161), .Y(n_282) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_162), .Y(n_171) );
INVx2_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_163), .A2(n_250), .B(n_252), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_163), .A2(n_265), .B(n_267), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_163), .A2(n_290), .B(n_292), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_163), .A2(n_596), .B(n_597), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_163), .A2(n_665), .B(n_666), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_163), .A2(n_681), .B(n_682), .Y(n_680) );
BUFx10_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g611 ( .A(n_164), .Y(n_611) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g569 ( .A(n_165), .Y(n_569) );
AO21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_172), .Y(n_166) );
INVx2_ASAP7_75t_L g268 ( .A(n_168), .Y(n_268) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
INVx2_ASAP7_75t_L g224 ( .A(n_171), .Y(n_224) );
INVx2_ASAP7_75t_L g253 ( .A(n_171), .Y(n_253) );
INVx3_ASAP7_75t_L g557 ( .A(n_171), .Y(n_557) );
INVx3_ASAP7_75t_L g623 ( .A(n_171), .Y(n_623) );
INVx2_ASAP7_75t_L g686 ( .A(n_171), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_172), .A2(n_262), .B(n_263), .Y(n_261) );
O2A1O1Ixp5_ASAP7_75t_L g683 ( .A1(n_172), .A2(n_684), .B(n_685), .C(n_687), .Y(n_683) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
INVx2_ASAP7_75t_L g228 ( .A(n_173), .Y(n_228) );
AOI211x1_ASAP7_75t_L g242 ( .A1(n_173), .A2(n_241), .B(n_243), .C(n_249), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_173), .B(n_643), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_173), .B(n_643), .C(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_175), .A2(n_181), .B(n_183), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVxp33_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx2_ASAP7_75t_L g182 ( .A(n_178), .Y(n_182) );
INVx1_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_178), .Y(n_240) );
INVx1_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx3_ASAP7_75t_L g214 ( .A(n_182), .Y(n_214) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_183), .A2(n_216), .B(n_222), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_183), .A2(n_239), .B(n_241), .Y(n_238) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_183), .A2(n_261), .B(n_264), .Y(n_260) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_183), .A2(n_592), .B(n_595), .Y(n_591) );
OAI21x1_ASAP7_75t_L g657 ( .A1(n_183), .A2(n_658), .B(n_664), .Y(n_657) );
BUFx6f_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
INVx1_ASAP7_75t_L g273 ( .A(n_184), .Y(n_273) );
INVx2_ASAP7_75t_L g299 ( .A(n_184), .Y(n_299) );
INVx3_ASAP7_75t_L g643 ( .A(n_184), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_186), .B(n_414), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_186), .B(n_359), .Y(n_441) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_213), .Y(n_186) );
AND2x2_ASAP7_75t_L g314 ( .A(n_187), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g310 ( .A(n_188), .Y(n_310) );
AND2x2_ASAP7_75t_L g352 ( .A(n_188), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g360 ( .A(n_188), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g381 ( .A(n_188), .Y(n_381) );
AND2x2_ASAP7_75t_L g401 ( .A(n_188), .B(n_213), .Y(n_401) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_188), .Y(n_437) );
INVxp67_ASAP7_75t_L g467 ( .A(n_188), .Y(n_467) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_195), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_191), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g344 ( .A(n_191), .Y(n_344) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
AOI21x1_ASAP7_75t_L g204 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_205), .B1(n_209), .B2(n_211), .Y(n_195) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .C(n_203), .Y(n_196) );
NAND3xp33_ASAP7_75t_L g209 ( .A(n_197), .B(n_203), .C(n_210), .Y(n_209) );
BUFx2_ASAP7_75t_L g632 ( .A(n_197), .Y(n_632) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_198), .A2(n_344), .B(n_563), .Y(n_570) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_200), .B(n_643), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_200), .B(n_643), .C(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g349 ( .A(n_201), .Y(n_349) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx3_ASAP7_75t_L g210 ( .A(n_202), .Y(n_210) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_203), .Y(n_637) );
NOR2xp33_ASAP7_75t_SL g652 ( .A(n_203), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_207), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g226 ( .A(n_208), .Y(n_226) );
INVx1_ASAP7_75t_L g291 ( .A(n_208), .Y(n_291) );
INVx2_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_L g293 ( .A1(n_210), .A2(n_294), .B(n_295), .C(n_296), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_210), .A2(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g312 ( .A(n_213), .Y(n_312) );
INVx1_ASAP7_75t_L g317 ( .A(n_213), .Y(n_317) );
INVx1_ASAP7_75t_L g361 ( .A(n_213), .Y(n_361) );
AND2x2_ASAP7_75t_L g539 ( .A(n_213), .B(n_448), .Y(n_539) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_229), .Y(n_213) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_214), .A2(n_657), .B(n_667), .Y(n_656) );
OAI21x1_ASAP7_75t_L g678 ( .A1(n_214), .A2(n_679), .B(n_688), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_219), .B(n_221), .Y(n_216) );
INVx2_ASAP7_75t_L g578 ( .A(n_218), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_218), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g582 ( .A(n_220), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_221), .A2(n_281), .B(n_283), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_225), .B(n_227), .Y(n_222) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_228), .B(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_230), .Y(n_604) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_254), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g382 ( .A(n_235), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g388 ( .A(n_235), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_235), .B(n_374), .Y(n_409) );
AND2x2_ASAP7_75t_L g433 ( .A(n_235), .B(n_319), .Y(n_433) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g356 ( .A(n_236), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g510 ( .A(n_236), .B(n_454), .Y(n_510) );
AND2x2_ASAP7_75t_L g516 ( .A(n_236), .B(n_335), .Y(n_516) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
AND2x2_ASAP7_75t_L g328 ( .A(n_237), .B(n_306), .Y(n_328) );
INVx2_ASAP7_75t_L g365 ( .A(n_237), .Y(n_365) );
INVx1_ASAP7_75t_L g397 ( .A(n_237), .Y(n_397) );
AND2x2_ASAP7_75t_L g404 ( .A(n_237), .B(n_357), .Y(n_404) );
AND2x2_ASAP7_75t_L g440 ( .A(n_237), .B(n_396), .Y(n_440) );
BUFx2_ASAP7_75t_L g479 ( .A(n_237), .Y(n_479) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_237), .Y(n_502) );
OR2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
NOR2xp67_ASAP7_75t_SL g272 ( .A(n_240), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g695 ( .A(n_240), .Y(n_695) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_248), .Y(n_243) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g266 ( .A(n_246), .Y(n_266) );
INVx2_ASAP7_75t_L g297 ( .A(n_246), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_246), .B(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_246), .Y(n_560) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_247), .Y(n_276) );
INVx2_ASAP7_75t_L g565 ( .A(n_251), .Y(n_565) );
INVxp67_ASAP7_75t_L g628 ( .A(n_253), .Y(n_628) );
INVxp67_ASAP7_75t_L g659 ( .A(n_253), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_254), .A2(n_358), .B1(n_399), .B2(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_285), .Y(n_255) );
INVx4_ASAP7_75t_L g319 ( .A(n_256), .Y(n_319) );
NAND2xp33_ASAP7_75t_SL g372 ( .A(n_256), .B(n_373), .Y(n_372) );
OAI32xp33_ASAP7_75t_L g517 ( .A1(n_256), .A2(n_402), .A3(n_518), .B1(n_519), .B2(n_521), .Y(n_517) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_270), .Y(n_256) );
INVx2_ASAP7_75t_L g369 ( .A(n_257), .Y(n_369) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_269), .Y(n_257) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_288), .B(n_300), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_258), .A2(n_260), .B(n_269), .Y(n_306) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_258), .A2(n_591), .B(n_599), .Y(n_590) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_258), .A2(n_620), .B(n_700), .Y(n_699) );
OAI21x1_ASAP7_75t_L g725 ( .A1(n_258), .A2(n_591), .B(n_599), .Y(n_725) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2x1_ASAP7_75t_SL g584 ( .A(n_259), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g625 ( .A(n_266), .Y(n_625) );
AND2x4_ASAP7_75t_L g307 ( .A(n_270), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g327 ( .A(n_270), .Y(n_327) );
INVx2_ASAP7_75t_L g357 ( .A(n_270), .Y(n_357) );
AND2x2_ASAP7_75t_L g383 ( .A(n_270), .B(n_369), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_270), .B(n_286), .Y(n_389) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_279), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_272), .A2(n_280), .B(n_284), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g338 ( .A(n_276), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_276), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g598 ( .A(n_276), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_276), .B(n_641), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_278), .A2(n_581), .B(n_583), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_282), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g471 ( .A(n_285), .B(n_404), .Y(n_471) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_285), .Y(n_520) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_286), .Y(n_331) );
AND2x2_ASAP7_75t_L g374 ( .A(n_286), .B(n_369), .Y(n_374) );
AND2x2_ASAP7_75t_L g453 ( .A(n_286), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g323 ( .A(n_287), .Y(n_323) );
INVx1_ASAP7_75t_L g368 ( .A(n_287), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_293), .B(n_298), .Y(n_288) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_SL g342 ( .A(n_299), .Y(n_342) );
INVx1_ASAP7_75t_L g614 ( .A(n_299), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_309), .B1(n_313), .B2(n_318), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_304), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g499 ( .A(n_304), .Y(n_499) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g406 ( .A(n_305), .B(n_322), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_305), .A2(n_412), .B1(n_492), .B2(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g464 ( .A(n_306), .B(n_357), .Y(n_464) );
AND2x2_ASAP7_75t_L g427 ( .A(n_307), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g449 ( .A(n_307), .B(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_307), .Y(n_508) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_308), .Y(n_495) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_310), .Y(n_391) );
AND2x2_ASAP7_75t_L g446 ( .A(n_310), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g456 ( .A(n_310), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g496 ( .A(n_310), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_310), .B(n_497), .Y(n_512) );
AND2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g475 ( .A(n_311), .Y(n_475) );
AOI33xp33_ASAP7_75t_L g509 ( .A1(n_311), .A2(n_319), .A3(n_392), .B1(n_510), .B2(n_511), .B3(n_516), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_313), .B(n_333), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_313), .A2(n_372), .B1(n_375), .B2(n_382), .Y(n_371) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AND2x2_ASAP7_75t_L g470 ( .A(n_314), .B(n_447), .Y(n_470) );
AND2x4_ASAP7_75t_L g538 ( .A(n_314), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g400 ( .A(n_315), .B(n_335), .Y(n_400) );
INVx1_ASAP7_75t_L g497 ( .A(n_315), .Y(n_497) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_317), .Y(n_378) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_318), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g493 ( .A(n_318), .Y(n_493) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_319), .A2(n_500), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g355 ( .A(n_321), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g418 ( .A(n_321), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_321), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_329), .B(n_332), .C(n_350), .Y(n_324) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_326), .A2(n_534), .B1(n_536), .B2(n_540), .Y(n_533) );
INVx4_ASAP7_75t_R g326 ( .A(n_327), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g498 ( .A1(n_327), .A2(n_499), .A3(n_500), .B1(n_501), .B2(n_503), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_327), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g330 ( .A(n_328), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g500 ( .A(n_333), .B(n_475), .Y(n_500) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_335), .Y(n_359) );
BUFx2_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
INVx1_ASAP7_75t_L g415 ( .A(n_335), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_336), .B(n_345), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_336), .B(n_345), .Y(n_353) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B(n_343), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_338), .A2(n_578), .B1(n_648), .B2(n_650), .Y(n_647) );
OR2x2_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g585 ( .A(n_342), .Y(n_585) );
INVxp67_ASAP7_75t_L g631 ( .A(n_344), .Y(n_631) );
INVx1_ASAP7_75t_L g561 ( .A(n_349), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_349), .A2(n_577), .B(n_579), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B1(n_358), .B2(n_362), .Y(n_350) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_351), .A2(n_443), .B1(n_449), .B2(n_451), .C1(n_456), .C2(n_458), .Y(n_442) );
AND2x2_ASAP7_75t_L g385 ( .A(n_352), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g380 ( .A(n_353), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g448 ( .A(n_353), .Y(n_448) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_355), .A2(n_435), .B1(n_439), .B2(n_441), .Y(n_434) );
INVx2_ASAP7_75t_L g455 ( .A(n_356), .Y(n_455) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_357), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x4_ASAP7_75t_SL g407 ( .A(n_360), .B(n_400), .Y(n_407) );
INVx1_ASAP7_75t_L g492 ( .A(n_360), .Y(n_492) );
AND2x2_ASAP7_75t_L g447 ( .A(n_361), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
INVx1_ASAP7_75t_L g459 ( .A(n_364), .Y(n_459) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_SL g428 ( .A(n_367), .Y(n_428) );
INVx1_ASAP7_75t_L g484 ( .A(n_367), .Y(n_484) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
BUFx2_ASAP7_75t_L g514 ( .A(n_368), .Y(n_514) );
INVx1_ASAP7_75t_L g454 ( .A(n_369), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_384), .C(n_398), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_374), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
OR2x2_ASAP7_75t_L g474 ( .A(n_379), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g487 ( .A(n_380), .B(n_386), .Y(n_487) );
INVx1_ASAP7_75t_L g413 ( .A(n_381), .Y(n_413) );
AND2x2_ASAP7_75t_L g394 ( .A(n_383), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_383), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g485 ( .A(n_383), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B1(n_390), .B2(n_394), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g423 ( .A(n_389), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g511 ( .A1(n_389), .A2(n_512), .B1(n_513), .B2(n_515), .Y(n_511) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_396), .Y(n_450) );
OR2x2_ASAP7_75t_L g535 ( .A(n_396), .B(n_397), .Y(n_535) );
AOI32xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .A3(n_405), .B1(n_407), .B2(n_408), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx2_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_401), .B(n_414), .Y(n_518) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g529 ( .A(n_405), .B(n_485), .C(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g482 ( .A(n_407), .Y(n_482) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_416), .B(n_420), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_418), .A2(n_491), .B1(n_493), .B2(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_488), .Y(n_424) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_426), .B(n_442), .C(n_460), .D(n_472), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g532 ( .A(n_430), .B(n_438), .Y(n_532) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
OR2x2_ASAP7_75t_L g521 ( .A(n_436), .B(n_475), .Y(n_521) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g457 ( .A(n_438), .Y(n_457) );
OR2x2_ASAP7_75t_L g491 ( .A(n_438), .B(n_492), .Y(n_491) );
OR2x2_ASAP7_75t_L g528 ( .A(n_438), .B(n_502), .Y(n_528) );
INVx1_ASAP7_75t_L g461 ( .A(n_439), .Y(n_461) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_441), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g540 ( .A(n_446), .B(n_497), .Y(n_540) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g526 ( .A(n_453), .Y(n_526) );
OAI32xp33_ASAP7_75t_L g481 ( .A1(n_458), .A2(n_482), .A3(n_483), .B1(n_485), .B2(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_465), .C(n_469), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g480 ( .A(n_464), .Y(n_480) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g530 ( .A(n_471), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_476), .B(n_481), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_489), .B(n_505), .C(n_522), .D(n_533), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .C(n_497), .Y(n_494) );
AOI322xp5_ASAP7_75t_L g522 ( .A1(n_499), .A2(n_523), .A3(n_524), .B1(n_525), .B2(n_527), .C1(n_529), .C2(n_531), .Y(n_522) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_500), .A2(n_507), .B(n_509), .Y(n_506) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_502), .Y(n_524) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_SL g505 ( .A(n_506), .B(n_517), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
BUFx8_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND3x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_821), .C(n_867), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_765), .Y(n_546) );
NAND3xp33_ASAP7_75t_SL g547 ( .A(n_548), .B(n_702), .C(n_737), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_586), .B1(n_689), .B2(n_696), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_571), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g817 ( .A(n_552), .B(n_589), .Y(n_817) );
AND2x4_ASAP7_75t_L g830 ( .A(n_552), .B(n_725), .Y(n_830) );
AND2x2_ASAP7_75t_L g861 ( .A(n_552), .B(n_746), .Y(n_861) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_552), .Y(n_894) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x6_ASAP7_75t_L g714 ( .A(n_553), .B(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_SL g726 ( .A(n_553), .B(n_693), .Y(n_726) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g692 ( .A(n_554), .Y(n_692) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_562), .B(n_570), .Y(n_554) );
AOI21x1_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_559), .B(n_561), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AOI22x1_ASAP7_75t_L g620 ( .A1(n_561), .A2(n_569), .B1(n_621), .B2(n_627), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_565), .A2(n_628), .B1(n_629), .B2(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI21x1_ASAP7_75t_L g606 ( .A1(n_569), .A2(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g806 ( .A(n_571), .B(n_807), .Y(n_806) );
OR2x2_ASAP7_75t_L g827 ( .A(n_571), .B(n_714), .Y(n_827) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g734 ( .A(n_572), .Y(n_734) );
AND2x2_ASAP7_75t_L g741 ( .A(n_572), .B(n_693), .Y(n_741) );
INVx2_ASAP7_75t_L g746 ( .A(n_572), .Y(n_746) );
AND2x2_ASAP7_75t_L g761 ( .A(n_572), .B(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g771 ( .A(n_572), .B(n_601), .Y(n_771) );
OR2x2_ASAP7_75t_L g787 ( .A(n_572), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g816 ( .A(n_572), .Y(n_816) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OAI21x1_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_580), .B(n_584), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_616), .B1(n_668), .B2(n_672), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g854 ( .A(n_588), .B(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_600), .Y(n_588) );
BUFx3_ASAP7_75t_L g670 ( .A(n_589), .Y(n_670) );
AND2x2_ASAP7_75t_L g759 ( .A(n_589), .B(n_734), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_589), .Y(n_762) );
AND2x2_ASAP7_75t_L g876 ( .A(n_589), .B(n_692), .Y(n_876) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_590), .Y(n_798) );
INVxp67_ASAP7_75t_L g612 ( .A(n_598), .Y(n_612) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_600), .Y(n_774) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_601), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_601), .B(n_692), .Y(n_807) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g715 ( .A(n_602), .Y(n_715) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_602), .Y(n_788) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_615), .Y(n_603) );
OA21x2_ASAP7_75t_L g693 ( .A1(n_605), .A2(n_615), .B(n_694), .Y(n_693) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B(n_614), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B(n_613), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g679 ( .A1(n_614), .A2(n_680), .B(n_683), .Y(n_679) );
INVx2_ASAP7_75t_L g767 ( .A(n_616), .Y(n_767) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_634), .Y(n_616) );
INVx1_ASAP7_75t_L g732 ( .A(n_617), .Y(n_732) );
INVx1_ASAP7_75t_L g764 ( .A(n_617), .Y(n_764) );
BUFx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g750 ( .A(n_618), .Y(n_750) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_631), .A3(n_632), .B(n_633), .Y(n_618) );
AO31x2_ASAP7_75t_L g782 ( .A1(n_619), .A2(n_631), .A3(n_632), .B(n_633), .Y(n_782) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22x1_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g700 ( .A(n_633), .Y(n_700) );
INVx1_ASAP7_75t_L g900 ( .A(n_634), .Y(n_900) );
INVxp67_ASAP7_75t_SL g911 ( .A(n_634), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_654), .Y(n_634) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_635), .B(n_676), .Y(n_675) );
BUFx2_ASAP7_75t_L g736 ( .A(n_635), .Y(n_736) );
INVx1_ASAP7_75t_L g778 ( .A(n_635), .Y(n_778) );
AND2x2_ASAP7_75t_L g837 ( .A(n_635), .B(n_655), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_635), .B(n_701), .Y(n_859) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g697 ( .A(n_636), .B(n_655), .Y(n_697) );
AO21x2_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B(n_652), .Y(n_636) );
AO21x1_ASAP7_75t_L g710 ( .A1(n_637), .A2(n_638), .B(n_652), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_647), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_644), .B2(n_646), .Y(n_639) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_655), .Y(n_674) );
INVx3_ASAP7_75t_L g706 ( .A(n_655), .Y(n_706) );
INVx2_ASAP7_75t_L g719 ( .A(n_655), .Y(n_719) );
AND2x2_ASAP7_75t_L g723 ( .A(n_655), .B(n_699), .Y(n_723) );
INVx1_ASAP7_75t_L g747 ( .A(n_655), .Y(n_747) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_661), .Y(n_658) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_670), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g785 ( .A(n_670), .Y(n_785) );
OR2x2_ASAP7_75t_L g826 ( .A(n_670), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
OR2x2_ASAP7_75t_L g906 ( .A(n_673), .B(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g722 ( .A(n_676), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_676), .B(n_706), .Y(n_755) );
NOR2xp67_ASAP7_75t_L g865 ( .A(n_676), .B(n_705), .Y(n_865) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g701 ( .A(n_677), .Y(n_701) );
AND2x2_ASAP7_75t_L g708 ( .A(n_677), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g820 ( .A(n_677), .B(n_699), .Y(n_820) );
INVx1_ASAP7_75t_L g843 ( .A(n_677), .Y(n_843) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_691), .A2(n_703), .B(n_711), .C(n_727), .Y(n_702) );
AND2x2_ASAP7_75t_L g851 ( .A(n_691), .B(n_815), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g904 ( .A(n_691), .B(n_746), .Y(n_904) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g730 ( .A(n_692), .Y(n_730) );
AND2x4_ASAP7_75t_L g740 ( .A(n_692), .B(n_725), .Y(n_740) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
AOI32xp33_ASAP7_75t_L g828 ( .A1(n_696), .A2(n_770), .A3(n_829), .B1(n_831), .B2(n_833), .Y(n_828) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
AND2x2_ASAP7_75t_L g819 ( .A(n_697), .B(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g720 ( .A(n_698), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_698), .B(n_778), .Y(n_794) );
AND2x2_ASAP7_75t_L g847 ( .A(n_698), .B(n_736), .Y(n_847) );
AND2x2_ASAP7_75t_L g910 ( .A(n_698), .B(n_911), .Y(n_910) );
AND2x4_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g757 ( .A(n_699), .Y(n_757) );
OR2x2_ASAP7_75t_L g781 ( .A(n_701), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
AOI21xp33_ASAP7_75t_SL g800 ( .A1(n_704), .A2(n_758), .B(n_799), .Y(n_800) );
OR2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
BUFx2_ASAP7_75t_L g845 ( .A(n_705), .Y(n_845) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_706), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g810 ( .A(n_706), .B(n_782), .Y(n_810) );
INVx1_ASAP7_75t_L g744 ( .A(n_707), .Y(n_744) );
OR2x2_ASAP7_75t_L g790 ( .A(n_707), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g749 ( .A(n_708), .Y(n_749) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_708), .Y(n_811) );
AND2x2_ASAP7_75t_L g852 ( .A(n_708), .B(n_750), .Y(n_852) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g718 ( .A(n_710), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_710), .B(n_757), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_716), .B1(n_721), .B2(n_724), .Y(n_711) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2x1p5_ASAP7_75t_L g760 ( .A(n_713), .B(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_713), .A2(n_883), .B1(n_885), .B2(n_887), .Y(n_882) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g803 ( .A(n_714), .B(n_746), .Y(n_803) );
AND2x2_ASAP7_75t_L g731 ( .A(n_715), .B(n_725), .Y(n_731) );
INVx2_ASAP7_75t_L g916 ( .A(n_716), .Y(n_916) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g824 ( .A(n_718), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g833 ( .A(n_718), .B(n_820), .Y(n_833) );
AND2x2_ASAP7_75t_L g872 ( .A(n_718), .B(n_764), .Y(n_872) );
AND2x2_ASAP7_75t_L g891 ( .A(n_718), .B(n_855), .Y(n_891) );
INVx1_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
OAI321xp33_ASAP7_75t_L g908 ( .A1(n_721), .A2(n_797), .A3(n_831), .B1(n_909), .B2(n_912), .C(n_915), .Y(n_908) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_722), .B(n_864), .Y(n_907) );
INVx1_ASAP7_75t_L g791 ( .A(n_723), .Y(n_791) );
AND2x4_ASAP7_75t_L g857 ( .A(n_723), .B(n_858), .Y(n_857) );
INVx3_ASAP7_75t_L g878 ( .A(n_724), .Y(n_878) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AND2x4_ASAP7_75t_L g770 ( .A(n_725), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g752 ( .A(n_726), .Y(n_752) );
NOR4xp25_ASAP7_75t_L g727 ( .A(n_728), .B(n_732), .C(n_733), .D(n_735), .Y(n_727) );
NAND2x1_ASAP7_75t_L g768 ( .A(n_728), .B(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_729), .A2(n_804), .B1(n_851), .B2(n_852), .Y(n_850) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
OAI322xp33_ASAP7_75t_L g889 ( .A1(n_732), .A2(n_890), .A3(n_892), .B1(n_898), .B2(n_901), .C1(n_902), .C2(n_906), .Y(n_889) );
AND2x2_ASAP7_75t_L g849 ( .A(n_733), .B(n_817), .Y(n_849) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g832 ( .A(n_734), .B(n_788), .Y(n_832) );
INVx1_ASAP7_75t_L g855 ( .A(n_734), .Y(n_855) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NOR2x1_ASAP7_75t_L g804 ( .A(n_736), .B(n_781), .Y(n_804) );
AOI211xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B(n_742), .C(n_753), .Y(n_737) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g813 ( .A(n_740), .Y(n_813) );
NOR2x1_ASAP7_75t_L g913 ( .A(n_740), .B(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g799 ( .A(n_741), .Y(n_799) );
O2A1O1Ixp33_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_745), .B(n_748), .C(n_751), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
AND2x2_ASAP7_75t_L g905 ( .A(n_746), .B(n_876), .Y(n_905) );
INVx2_ASAP7_75t_L g780 ( .A(n_747), .Y(n_780) );
OR2x6_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx2_ASAP7_75t_L g825 ( .A(n_750), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_750), .B(n_837), .Y(n_836) );
NAND2xp33_ASAP7_75t_SL g887 ( .A(n_751), .B(n_888), .Y(n_887) );
INVx2_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
OAI32xp33_ASAP7_75t_L g753 ( .A1(n_752), .A2(n_754), .A3(n_758), .B1(n_760), .B2(n_763), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_752), .B(n_855), .Y(n_901) );
OR2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g864 ( .A(n_756), .Y(n_864) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g835 ( .A(n_762), .B(n_807), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_783), .C(n_801), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_772), .B2(n_775), .Y(n_766) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
O2A1O1Ixp5_ASAP7_75t_L g812 ( .A1(n_771), .A2(n_813), .B(n_814), .C(n_818), .Y(n_812) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_771), .Y(n_870) );
INVx1_ASAP7_75t_L g914 ( .A(n_771), .Y(n_914) );
INVxp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g881 ( .A(n_777), .Y(n_881) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g886 ( .A(n_778), .B(n_843), .Y(n_886) );
INVx1_ASAP7_75t_L g793 ( .A(n_779), .Y(n_793) );
NOR2x1p5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g844 ( .A(n_782), .Y(n_844) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_789), .B1(n_792), .B2(n_795), .C(n_800), .Y(n_783) );
INVx1_ASAP7_75t_L g839 ( .A(n_784), .Y(n_839) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
OR2x2_ASAP7_75t_L g874 ( .A(n_787), .B(n_875), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_789), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AND2x2_ASAP7_75t_L g866 ( .A(n_798), .B(n_832), .Y(n_866) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_804), .B1(n_805), .B2(n_808), .C(n_812), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
AND2x4_ASAP7_75t_L g885 ( .A(n_809), .B(n_886), .Y(n_885) );
INVx2_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
OR2x2_ASAP7_75t_L g884 ( .A(n_810), .B(n_859), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx3_ASAP7_75t_R g888 ( .A(n_817), .Y(n_888) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR4xp25_ASAP7_75t_L g821 ( .A(n_822), .B(n_834), .C(n_838), .D(n_853), .Y(n_821) );
OAI21xp33_ASAP7_75t_SL g822 ( .A1(n_823), .A2(n_826), .B(n_828), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AOI21xp33_ASAP7_75t_SL g834 ( .A1(n_826), .A2(n_835), .B(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g915 ( .A1(n_830), .A2(n_866), .B(n_916), .Y(n_915) );
BUFx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI221xp5_ASAP7_75t_SL g838 ( .A1(n_839), .A2(n_840), .B1(n_846), .B2(n_848), .C(n_850), .Y(n_838) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_840), .A2(n_854), .B1(n_856), .B2(n_860), .C(n_862), .Y(n_853) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_842), .B(n_845), .Y(n_841) );
INVx1_ASAP7_75t_L g880 ( .A(n_842), .Y(n_880) );
AND2x4_ASAP7_75t_L g899 ( .A(n_842), .B(n_900), .Y(n_899) );
AND2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
INVx1_ASAP7_75t_L g896 ( .A(n_843), .Y(n_896) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVxp67_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_855), .B(n_878), .C(n_879), .D(n_881), .Y(n_877) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVxp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_866), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
NOR3xp33_ASAP7_75t_L g867 ( .A(n_868), .B(n_889), .C(n_908), .Y(n_867) );
NAND4xp25_ASAP7_75t_L g868 ( .A(n_869), .B(n_871), .C(n_877), .D(n_882), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_876), .Y(n_897) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NOR2xp33_ASAP7_75t_SL g892 ( .A(n_893), .B(n_897), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g926 ( .A(n_919), .Y(n_926) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
BUFx3_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
AND2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
OAI21xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_946), .B(n_950), .Y(n_935) );
OR2x2_ASAP7_75t_L g936 ( .A(n_937), .B(n_943), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_939), .Y(n_938) );
HB1xp67_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_SL g946 ( .A(n_947), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_947), .B(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
HB1xp67_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
BUFx3_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .Y(n_956) );
endmodule