module fake_ariane_392_n_1995 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1995);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1995;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1865;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_47),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_98),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_2),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_25),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_20),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_36),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_38),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_29),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_116),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_9),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_66),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_165),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_93),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_7),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_23),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_32),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_106),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_4),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_148),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_188),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_130),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_44),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_127),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_190),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_70),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_88),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_6),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_149),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_123),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_23),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_112),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_104),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_162),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_199),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_119),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_50),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_58),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_109),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_67),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_29),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_142),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_70),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_69),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_85),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_122),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_74),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_87),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_171),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_55),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_99),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_128),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_167),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_115),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_63),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_191),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_7),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_134),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_192),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_105),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_79),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_19),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_28),
.Y(n_296)
);

BUFx2_ASAP7_75t_SL g297 ( 
.A(n_176),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_69),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_8),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_103),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_154),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_193),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_45),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_82),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_37),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_152),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_94),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_95),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_178),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_83),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_51),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_67),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_145),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_44),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_175),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_12),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_22),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_139),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_56),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_27),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_17),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_170),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_59),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_202),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_60),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_133),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_33),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_68),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_28),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_8),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_10),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_77),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_73),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_5),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_100),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_131),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_111),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_113),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_38),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_50),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_184),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_129),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_60),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_62),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_56),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_49),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_27),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_30),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_164),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_91),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_48),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_58),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_78),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_66),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_32),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_89),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_159),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_53),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_177),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_120),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_42),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_19),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_151),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_71),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_117),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_75),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_124),
.Y(n_370)
);

BUFx8_ASAP7_75t_SL g371 ( 
.A(n_185),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_61),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_195),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_90),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_169),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_72),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_80),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_59),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_30),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_54),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_21),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_6),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_36),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_160),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_26),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_138),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_39),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_43),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_42),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_136),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_37),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_157),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_135),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_96),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_186),
.Y(n_396)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_3),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_57),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_97),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_161),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_40),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_64),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_114),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_121),
.Y(n_404)
);

INVx4_ASAP7_75t_R g405 ( 
.A(n_214),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_216),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_216),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_210),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_241),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_241),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_210),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_236),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_236),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_220),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_220),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_371),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_288),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_227),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_R g419 ( 
.A(n_261),
.B(n_76),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_269),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_269),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_334),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_285),
.B(n_0),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_349),
.B(n_1),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_354),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_269),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_213),
.B(n_1),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_371),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_229),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_226),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_226),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_269),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_233),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_233),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_228),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_271),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_271),
.Y(n_438)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_207),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_228),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_389),
.B(n_3),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_269),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_214),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_209),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_211),
.B(n_9),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_300),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_269),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_269),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_300),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_321),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_314),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_314),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_229),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_321),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_228),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_217),
.B(n_10),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_224),
.B(n_11),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_352),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_243),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_321),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_321),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_257),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_321),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_352),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_205),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_321),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_223),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_212),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_360),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_360),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_225),
.B(n_11),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_366),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_321),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_366),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_367),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_367),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_390),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_374),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

BUFx6f_ASAP7_75t_SL g483 ( 
.A(n_244),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_228),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_R g487 ( 
.A(n_315),
.B(n_201),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_374),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_209),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_209),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_255),
.B(n_14),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_258),
.B(n_259),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_234),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_391),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_391),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_396),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_223),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_218),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_213),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_396),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_208),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_219),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_239),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_239),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_273),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_235),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_409),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_409),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_420),
.A2(n_274),
.B(n_262),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_491),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_414),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_410),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_421),
.A2(n_280),
.B(n_275),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_410),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_416),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_459),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_416),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_489),
.A2(n_442),
.B(n_426),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_428),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_415),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_459),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_428),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_406),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_431),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_448),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_450),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_454),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_432),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_461),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_432),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_468),
.B(n_238),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_485),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_466),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_473),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_413),
.B(n_282),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_476),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_478),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_481),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_449),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_485),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_439),
.B(n_234),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_443),
.B(n_284),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_434),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_504),
.B(n_234),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_290),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_435),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_418),
.B(n_204),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_494),
.B(n_244),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_484),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_406),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_486),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_492),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_443),
.B(n_291),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_419),
.B(n_372),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_493),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_422),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_R g581 ( 
.A(n_468),
.B(n_315),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_429),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_458),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_507),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_462),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_435),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_436),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_437),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_437),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_503),
.B(n_244),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_440),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_483),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_438),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_438),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_483),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_477),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_497),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_462),
.B(n_301),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_559),
.B(n_250),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_503),
.Y(n_602)
);

OAI22x1_ASAP7_75t_SL g603 ( 
.A1(n_519),
.A2(n_407),
.B1(n_511),
.B2(n_510),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_522),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_465),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_587),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_587),
.B(n_444),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_498),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_529),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_591),
.B(n_596),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_585),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_544),
.B(n_453),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_596),
.B(n_445),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_565),
.B(n_441),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_532),
.Y(n_616)
);

AND2x6_ASAP7_75t_L g617 ( 
.A(n_559),
.B(n_250),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_530),
.B(n_456),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_522),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_529),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_568),
.B(n_453),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_515),
.B(n_215),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_572),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_585),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_584),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_515),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_523),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_555),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_523),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_427),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_583),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_549),
.B(n_427),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_584),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_530),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_584),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_592),
.B(n_423),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_585),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_585),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_584),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_537),
.B(n_457),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_584),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_560),
.Y(n_644)
);

AND3x1_ASAP7_75t_L g645 ( 
.A(n_564),
.B(n_424),
.C(n_471),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_538),
.B(n_495),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_592),
.B(n_373),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_595),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_564),
.B(n_303),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_539),
.B(n_408),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_580),
.B(n_483),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_539),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_597),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_536),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_540),
.B(n_411),
.Y(n_657)
);

INVx4_ASAP7_75t_SL g658 ( 
.A(n_542),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_592),
.B(n_373),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_517),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_563),
.Y(n_662)
);

BUFx8_ASAP7_75t_SL g663 ( 
.A(n_535),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_546),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_546),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_547),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_548),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_514),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_548),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_550),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_517),
.A2(n_425),
.B1(n_328),
.B2(n_290),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_581),
.A2(n_487),
.B1(n_348),
.B2(n_379),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_550),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_552),
.B(n_303),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_595),
.B(n_404),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_527),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_552),
.B(n_412),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_575),
.B(n_508),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_553),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_590),
.A2(n_348),
.B1(n_379),
.B2(n_273),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_595),
.B(n_417),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_554),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_563),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_570),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_599),
.B(n_430),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_570),
.B(n_573),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_580),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_576),
.A2(n_401),
.B1(n_265),
.B2(n_231),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_569),
.B(n_573),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_574),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_574),
.B(n_509),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_577),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_577),
.A2(n_401),
.B1(n_230),
.B2(n_245),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_516),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_517),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_520),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_525),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_578),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_527),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_578),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_517),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_545),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_545),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_533),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_527),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_545),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_527),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_526),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_561),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_558),
.B(n_513),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_528),
.B(n_531),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_558),
.B(n_446),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_521),
.Y(n_716)
);

BUFx4f_ASAP7_75t_L g717 ( 
.A(n_521),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_527),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_SL g719 ( 
.A(n_534),
.B(n_372),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_518),
.B(n_502),
.Y(n_720)
);

BUFx8_ASAP7_75t_SL g721 ( 
.A(n_535),
.Y(n_721)
);

NOR2x1p5_ASAP7_75t_L g722 ( 
.A(n_541),
.B(n_543),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_521),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_521),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_518),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_561),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_551),
.B(n_203),
.Y(n_728)
);

BUFx4f_ASAP7_75t_L g729 ( 
.A(n_551),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_551),
.B(n_292),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_571),
.A2(n_328),
.B1(n_249),
.B2(n_267),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_557),
.B(n_404),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_557),
.B(n_252),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_594),
.B(n_446),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_557),
.B(n_252),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_557),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_571),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_562),
.A2(n_341),
.B1(n_338),
.B2(n_340),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_566),
.B(n_297),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_586),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_593),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_738),
.A2(n_452),
.B1(n_464),
.B2(n_451),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_644),
.B(n_451),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_634),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_602),
.B(n_588),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_589),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_662),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_632),
.B(n_464),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_601),
.B(n_469),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_634),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_662),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_647),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_737),
.B(n_469),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_632),
.B(n_470),
.Y(n_754)
);

AOI221xp5_ASAP7_75t_L g755 ( 
.A1(n_645),
.A2(n_488),
.B1(n_505),
.B2(n_501),
.C(n_500),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_662),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_612),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_647),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_613),
.B(n_346),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_737),
.B(n_472),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_600),
.A2(n_270),
.B1(n_296),
.B2(n_254),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_672),
.A2(n_474),
.B1(n_475),
.B2(n_472),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_691),
.B(n_605),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_650),
.A2(n_499),
.B1(n_505),
.B2(n_501),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_601),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_616),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_606),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_685),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_659),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_659),
.Y(n_770)
);

O2A1O1Ixp5_ASAP7_75t_L g771 ( 
.A1(n_653),
.A2(n_339),
.B(n_344),
.C(n_362),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_716),
.B(n_320),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_606),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_650),
.B(n_488),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_600),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_600),
.A2(n_357),
.B1(n_330),
.B2(n_351),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_616),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_655),
.B(n_500),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_715),
.B(n_232),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_600),
.B(n_251),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_666),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_630),
.B(n_298),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_720),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_630),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_630),
.B(n_299),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_600),
.B(n_266),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_272),
.Y(n_787)
);

OAI21xp33_ASAP7_75t_L g788 ( 
.A1(n_618),
.A2(n_281),
.B(n_278),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_600),
.B(n_295),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_685),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_628),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_649),
.B(n_372),
.Y(n_793)
);

NOR2x1p5_ASAP7_75t_L g794 ( 
.A(n_696),
.B(n_302),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_655),
.B(n_479),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_720),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_617),
.B(n_304),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_617),
.B(n_306),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_741),
.B(n_312),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_627),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_609),
.B(n_313),
.Y(n_801)
);

BUFx12f_ASAP7_75t_L g802 ( 
.A(n_668),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_607),
.B(n_316),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_617),
.B(n_678),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_617),
.B(n_678),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_741),
.B(n_318),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_617),
.B(n_322),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_617),
.B(n_323),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_678),
.B(n_324),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_643),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_689),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_688),
.A2(n_341),
.B(n_311),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_668),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_687),
.B(n_326),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_643),
.B(n_332),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_666),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_621),
.B(n_512),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_687),
.B(n_337),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_631),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_641),
.B(n_342),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_673),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_656),
.B(n_343),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_725),
.B(n_319),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_740),
.B(n_350),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_734),
.B(n_355),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_669),
.B(n_358),
.Y(n_826)
);

INVx8_ASAP7_75t_L g827 ( 
.A(n_739),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_669),
.B(n_361),
.Y(n_828)
);

BUFx8_ASAP7_75t_L g829 ( 
.A(n_725),
.Y(n_829)
);

INVx8_ASAP7_75t_L g830 ( 
.A(n_739),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_646),
.B(n_615),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_670),
.B(n_364),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_696),
.B(n_310),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_658),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_671),
.A2(n_331),
.B1(n_347),
.B2(n_333),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_612),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_700),
.B(n_381),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_694),
.A2(n_380),
.B(n_386),
.C(n_365),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_694),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_615),
.A2(n_327),
.B1(n_335),
.B2(n_336),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_698),
.B(n_376),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_700),
.A2(n_377),
.B1(n_394),
.B2(n_395),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_668),
.B(n_382),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_703),
.A2(n_383),
.B1(n_384),
.B2(n_402),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_703),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_623),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_614),
.B(n_388),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_611),
.B(n_392),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_681),
.A2(n_400),
.B1(n_403),
.B2(n_206),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_739),
.B(n_257),
.Y(n_850)
);

AOI22x1_ASAP7_75t_L g851 ( 
.A1(n_626),
.A2(n_320),
.B1(n_399),
.B2(n_338),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_679),
.B(n_682),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_684),
.B(n_15),
.Y(n_853)
);

AND2x2_ASAP7_75t_SL g854 ( 
.A(n_622),
.B(n_340),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_738),
.A2(n_674),
.B1(n_717),
.B2(n_716),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_681),
.B(n_372),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_626),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_652),
.B(n_221),
.Y(n_858)
);

NAND2x1_ASAP7_75t_L g859 ( 
.A(n_625),
.B(n_405),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_714),
.B(n_222),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_654),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_629),
.B(n_398),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_629),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_693),
.B(n_398),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_653),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_664),
.B(n_665),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_664),
.B(n_237),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_675),
.B(n_17),
.Y(n_868)
);

AOI221xp5_ASAP7_75t_L g869 ( 
.A1(n_695),
.A2(n_399),
.B1(n_385),
.B2(n_240),
.C(n_393),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_665),
.A2(n_686),
.B1(n_702),
.B2(n_692),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_667),
.B(n_242),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_667),
.B(n_246),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_698),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_683),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_663),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_738),
.A2(n_293),
.B1(n_378),
.B2(n_375),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_699),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_690),
.B(n_247),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_686),
.B(n_248),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_651),
.B(n_657),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_636),
.B(n_253),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_680),
.B(n_305),
.C(n_370),
.Y(n_882)
);

BUFx6f_ASAP7_75t_SL g883 ( 
.A(n_711),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_831),
.A2(n_620),
.B(n_610),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_766),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_834),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_763),
.A2(n_709),
.B(n_705),
.C(n_706),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_866),
.A2(n_620),
.B(n_610),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_834),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_763),
.B(n_699),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_765),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_880),
.B(n_604),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_880),
.A2(n_717),
.B(n_622),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_767),
.B(n_711),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_852),
.A2(n_717),
.B(n_697),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_765),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_800),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_857),
.B(n_604),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_L g899 ( 
.A(n_825),
.B(n_731),
.C(n_719),
.Y(n_899)
);

NAND3xp33_ASAP7_75t_L g900 ( 
.A(n_779),
.B(n_719),
.C(n_677),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_863),
.B(n_619),
.Y(n_901)
);

AND2x2_ASAP7_75t_SL g902 ( 
.A(n_855),
.B(n_603),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_779),
.A2(n_801),
.B1(n_787),
.B2(n_848),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_771),
.A2(n_704),
.B(n_661),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_L g905 ( 
.A(n_802),
.B(n_713),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_791),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_745),
.A2(n_709),
.B(n_706),
.C(n_705),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_771),
.A2(n_704),
.B(n_661),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_810),
.B(n_625),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_767),
.B(n_711),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_784),
.B(n_722),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_759),
.A2(n_648),
.B(n_660),
.C(n_625),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_787),
.A2(n_738),
.B1(n_674),
.B2(n_633),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_827),
.B(n_663),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_791),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_777),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_870),
.A2(n_724),
.B(n_697),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_784),
.B(n_658),
.Y(n_918)
);

OR2x6_ASAP7_75t_SL g919 ( 
.A(n_778),
.B(n_721),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_757),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_744),
.A2(n_723),
.B1(n_704),
.B2(n_661),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_747),
.A2(n_724),
.B(n_642),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_751),
.A2(n_768),
.B(n_756),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_848),
.B(n_619),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_801),
.A2(n_732),
.B(n_635),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_773),
.B(n_721),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_750),
.A2(n_723),
.B(n_633),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_862),
.A2(n_635),
.B(n_642),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_847),
.B(n_674),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_752),
.A2(n_723),
.B(n_735),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_820),
.B(n_674),
.Y(n_931)
);

OAI321xp33_ASAP7_75t_L g932 ( 
.A1(n_762),
.A2(n_733),
.A3(n_730),
.B1(n_728),
.B2(n_712),
.C(n_707),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_815),
.B(n_674),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_758),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_773),
.B(n_624),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_743),
.B(n_624),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_769),
.A2(n_736),
.B1(n_708),
.B2(n_718),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_815),
.B(n_624),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_810),
.B(n_658),
.Y(n_939)
);

BUFx4f_ASAP7_75t_L g940 ( 
.A(n_827),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_813),
.B(n_658),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_770),
.A2(n_729),
.B(n_736),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_875),
.B(n_638),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_790),
.A2(n_638),
.B(n_639),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_792),
.A2(n_638),
.B(n_639),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_781),
.A2(n_729),
.B(n_708),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_762),
.B(n_637),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_816),
.A2(n_736),
.B(n_708),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_821),
.A2(n_718),
.B(n_637),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_819),
.B(n_718),
.Y(n_950)
);

OAI21xp33_ASAP7_75t_L g951 ( 
.A1(n_759),
.A2(n_803),
.B(n_853),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_826),
.B(n_640),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_819),
.B(n_640),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_746),
.B(n_640),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_764),
.B(n_833),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_839),
.A2(n_727),
.B(n_726),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_845),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_861),
.B(n_707),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_865),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_757),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_868),
.A2(n_853),
.B(n_869),
.C(n_881),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_874),
.A2(n_726),
.B(n_712),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_793),
.A2(n_710),
.B(n_701),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_836),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_829),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_835),
.B(n_701),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_835),
.B(n_854),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_826),
.B(n_710),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_854),
.B(n_701),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_804),
.B(n_710),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_829),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_875),
.B(n_676),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_795),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_846),
.A2(n_676),
.B(n_215),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_796),
.B(n_260),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_867),
.A2(n_676),
.B(n_309),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_805),
.B(n_676),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_871),
.A2(n_676),
.B(n_317),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_836),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_749),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_841),
.B(n_263),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_811),
.B(n_294),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_872),
.A2(n_289),
.B(n_369),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_879),
.A2(n_287),
.B(n_368),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_868),
.A2(n_307),
.B(n_363),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_864),
.A2(n_268),
.B(n_215),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_836),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_796),
.B(n_264),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_803),
.A2(n_387),
.B(n_329),
.C(n_356),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_772),
.B(n_215),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_828),
.A2(n_329),
.B(n_353),
.C(n_345),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_849),
.B(n_276),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_780),
.A2(n_359),
.B(n_325),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_783),
.B(n_18),
.Y(n_994)
);

O2A1O1Ixp5_ASAP7_75t_L g995 ( 
.A1(n_812),
.A2(n_806),
.B(n_799),
.C(n_837),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_850),
.B(n_18),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_836),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_851),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_782),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_786),
.A2(n_308),
.B(n_286),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_772),
.B(n_268),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_814),
.A2(n_283),
.B(n_279),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_782),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_772),
.B(n_268),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_877),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_828),
.A2(n_277),
.B(n_256),
.C(n_243),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_789),
.A2(n_256),
.B(n_243),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_797),
.A2(n_256),
.B(n_243),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_832),
.A2(n_256),
.B(n_25),
.C(n_26),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_775),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_785),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_755),
.B(n_24),
.C(n_31),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_798),
.A2(n_268),
.B(n_215),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_807),
.A2(n_268),
.B(n_215),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_859),
.B(n_102),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_832),
.A2(n_268),
.B1(n_215),
.B2(n_34),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_808),
.A2(n_268),
.B(n_101),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_837),
.B(n_24),
.Y(n_1018)
);

OAI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_748),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_873),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_818),
.A2(n_35),
.B(n_39),
.C(n_40),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_809),
.B(n_41),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_785),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_858),
.B(n_860),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_873),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_856),
.A2(n_775),
.B(n_788),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_775),
.A2(n_110),
.B(n_194),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_817),
.B(n_108),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_823),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_827),
.B(n_830),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_754),
.B(n_823),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_830),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_761),
.B(n_43),
.Y(n_1033)
);

INVx11_ASAP7_75t_L g1034 ( 
.A(n_883),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_838),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_L g1036 ( 
.A(n_742),
.B(n_45),
.C(n_46),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_L g1037 ( 
.A1(n_753),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_761),
.A2(n_49),
.B(n_52),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_774),
.B(n_52),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_823),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_842),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_776),
.B(n_53),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_742),
.B(n_54),
.C(n_55),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_760),
.A2(n_126),
.B(n_182),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_776),
.B(n_57),
.Y(n_1045)
);

INVxp33_ASAP7_75t_SL g1046 ( 
.A(n_843),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_822),
.A2(n_118),
.B(n_174),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_850),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_882),
.B(n_61),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_893),
.A2(n_855),
.B(n_824),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_897),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_892),
.A2(n_878),
.B(n_850),
.Y(n_1052)
);

O2A1O1Ixp5_ASAP7_75t_L g1053 ( 
.A1(n_961),
.A2(n_844),
.B(n_772),
.C(n_876),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_892),
.A2(n_830),
.B(n_840),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_888),
.A2(n_772),
.B(n_794),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_890),
.B(n_62),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_903),
.A2(n_883),
.B(n_64),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_1034),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_884),
.A2(n_140),
.B(n_163),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_934),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_951),
.B(n_65),
.C(n_68),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_957),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_959),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_986),
.A2(n_86),
.B(n_92),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_980),
.B(n_107),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_974),
.A2(n_141),
.B(n_144),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_SL g1067 ( 
.A1(n_1024),
.A2(n_146),
.B(n_156),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_891),
.B(n_896),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_927),
.A2(n_930),
.B(n_921),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_924),
.A2(n_938),
.B(n_968),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_921),
.A2(n_908),
.B(n_904),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_929),
.A2(n_931),
.B(n_952),
.Y(n_1072)
);

AOI211x1_ASAP7_75t_L g1073 ( 
.A1(n_1038),
.A2(n_1019),
.B(n_1012),
.C(n_985),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_917),
.A2(n_928),
.B(n_922),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1041),
.B(n_1031),
.Y(n_1075)
);

CKINVDCx10_ASAP7_75t_R g1076 ( 
.A(n_914),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_999),
.B(n_1003),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_1010),
.Y(n_1078)
);

OAI22x1_ASAP7_75t_L g1079 ( 
.A1(n_1036),
.A2(n_1043),
.B1(n_996),
.B2(n_1040),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_1010),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_904),
.A2(n_887),
.B(n_900),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_1038),
.A2(n_942),
.B(n_1018),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_894),
.B(n_910),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_1032),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_936),
.A2(n_933),
.B(n_946),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_902),
.A2(n_967),
.B1(n_899),
.B2(n_985),
.Y(n_1086)
);

OA21x2_ASAP7_75t_L g1087 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1007),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_906),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_923),
.A2(n_956),
.B(n_949),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_947),
.B(n_975),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1002),
.A2(n_1009),
.B1(n_1022),
.B2(n_991),
.C(n_1021),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_898),
.A2(n_901),
.B(n_937),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_948),
.A2(n_901),
.B(n_898),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1008),
.A2(n_962),
.B(n_1017),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_989),
.A2(n_1001),
.A3(n_990),
.B(n_1004),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_998),
.A2(n_963),
.B(n_937),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_988),
.B(n_1011),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_990),
.A2(n_1004),
.B(n_1001),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1049),
.A2(n_1016),
.B(n_1002),
.C(n_967),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_1033),
.A2(n_1042),
.B(n_1035),
.C(n_995),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_925),
.A2(n_945),
.B(n_944),
.Y(n_1101)
);

BUFx2_ASAP7_75t_SL g1102 ( 
.A(n_916),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_907),
.A2(n_1006),
.B(n_1039),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1046),
.B(n_1020),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_885),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_969),
.A2(n_978),
.B(n_976),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_SL g1107 ( 
.A1(n_912),
.A2(n_1044),
.B(n_1026),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_970),
.A2(n_969),
.B(n_935),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_966),
.A2(n_970),
.A3(n_977),
.B(n_987),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_932),
.A2(n_913),
.B(n_966),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_993),
.A2(n_1000),
.B(n_977),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1015),
.A2(n_1027),
.B(n_909),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_955),
.A2(n_915),
.B(n_973),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1023),
.B(n_950),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_994),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1015),
.A2(n_909),
.B(n_939),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1025),
.B(n_1029),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_994),
.B(n_953),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_920),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_914),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_911),
.B(n_1005),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_983),
.A2(n_984),
.B(n_954),
.Y(n_1122)
);

NAND2x1_ASAP7_75t_L g1123 ( 
.A(n_886),
.B(n_889),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1037),
.A2(n_979),
.B(n_992),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_911),
.B(n_926),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1028),
.A2(n_1045),
.B(n_1047),
.C(n_996),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_943),
.B(n_958),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_981),
.A2(n_997),
.B(n_889),
.Y(n_1128)
);

AOI21x1_ASAP7_75t_L g1129 ( 
.A1(n_972),
.A2(n_982),
.B(n_1048),
.Y(n_1129)
);

CKINVDCx8_ASAP7_75t_R g1130 ( 
.A(n_914),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_960),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_940),
.B(n_982),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_960),
.B(n_964),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_905),
.A2(n_964),
.B(n_941),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1030),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1030),
.B(n_965),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_971),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_919),
.A2(n_903),
.B(n_951),
.C(n_961),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1030),
.A2(n_893),
.B(n_892),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_890),
.B(n_796),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_890),
.B(n_796),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_890),
.B(n_763),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_903),
.A2(n_890),
.B1(n_961),
.B2(n_951),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_903),
.A2(n_890),
.B1(n_961),
.B2(n_951),
.Y(n_1146)
);

NAND2x1p5_ASAP7_75t_L g1147 ( 
.A(n_1010),
.B(n_918),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_897),
.Y(n_1148)
);

AOI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_903),
.A2(n_825),
.B(n_581),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_1030),
.B(n_775),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1151)
);

OAI22x1_ASAP7_75t_L g1152 ( 
.A1(n_1036),
.A2(n_672),
.B1(n_680),
.B2(n_1043),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_890),
.B(n_763),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_903),
.A2(n_961),
.B(n_763),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_890),
.B(n_763),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_890),
.A2(n_763),
.B1(n_951),
.B2(n_755),
.C(n_762),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_903),
.A2(n_961),
.B(n_763),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_916),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_903),
.A2(n_961),
.B(n_763),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_906),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_SL g1163 ( 
.A(n_903),
.B(n_951),
.C(n_961),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_921),
.A2(n_961),
.A3(n_895),
.B(n_870),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_890),
.B(n_763),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1036),
.A2(n_1043),
.B1(n_902),
.B2(n_951),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_888),
.A2(n_884),
.B(n_986),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1034),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_888),
.A2(n_884),
.B(n_986),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1030),
.B(n_1032),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_896),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_934),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1034),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_890),
.B(n_903),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_903),
.A2(n_961),
.B(n_763),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_893),
.A2(n_892),
.B(n_903),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1155),
.A2(n_1161),
.B(n_1159),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1142),
.B(n_1153),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1157),
.A2(n_1179),
.B1(n_1149),
.B2(n_1146),
.C(n_1145),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1143),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1060),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1180),
.B(n_1090),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1189)
);

BUFx8_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1156),
.A2(n_1167),
.B1(n_1138),
.B2(n_1169),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1150),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1068),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1160),
.Y(n_1194)
);

NAND2xp33_ASAP7_75t_L g1195 ( 
.A(n_1083),
.B(n_1138),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1058),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1104),
.B(n_1141),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1086),
.B(n_1163),
.Y(n_1198)
);

AOI211xp5_ASAP7_75t_L g1199 ( 
.A1(n_1163),
.A2(n_1057),
.B(n_1056),
.C(n_1099),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1086),
.B(n_1144),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1174),
.B(n_1104),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1076),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1144),
.B(n_1151),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1088),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1151),
.B(n_1158),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1121),
.B(n_1125),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1099),
.A2(n_1053),
.B(n_1054),
.C(n_1169),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1174),
.B(n_1162),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1073),
.A2(n_1152),
.B1(n_1079),
.B2(n_1057),
.C(n_1053),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1058),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1097),
.B(n_1117),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1160),
.Y(n_1212)
);

NOR2x1_ASAP7_75t_L g1213 ( 
.A(n_1102),
.B(n_1105),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1154),
.B(n_1165),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1062),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1051),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1181),
.A2(n_1166),
.B(n_1168),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1176),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1171),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1118),
.A2(n_1061),
.B1(n_1075),
.B2(n_1054),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1168),
.A2(n_1177),
.B(n_1175),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1132),
.B(n_1113),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1178),
.Y(n_1223)
);

AND2x6_ASAP7_75t_L g1224 ( 
.A(n_1173),
.B(n_1135),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1175),
.A2(n_1070),
.B(n_1092),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_R g1226 ( 
.A(n_1130),
.B(n_1120),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1115),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1136),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1071),
.A2(n_1069),
.B1(n_1093),
.B2(n_1126),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1150),
.B(n_1084),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1091),
.B(n_1081),
.C(n_1050),
.Y(n_1231)
);

INVx3_ASAP7_75t_SL g1232 ( 
.A(n_1084),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1077),
.B(n_1065),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1134),
.B(n_1078),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1052),
.A2(n_1050),
.B(n_1100),
.C(n_1139),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1078),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1063),
.A2(n_1052),
.B1(n_1114),
.B2(n_1100),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1108),
.B(n_1110),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_1078),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1078),
.B(n_1080),
.Y(n_1240)
);

NAND3xp33_ASAP7_75t_L g1241 ( 
.A(n_1103),
.B(n_1124),
.C(n_1085),
.Y(n_1241)
);

AND2x6_ASAP7_75t_L g1242 ( 
.A(n_1080),
.B(n_1131),
.Y(n_1242)
);

AOI21xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1133),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1080),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1080),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1123),
.B(n_1129),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1072),
.A2(n_1101),
.B(n_1111),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1089),
.B(n_1101),
.C(n_1122),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1110),
.A2(n_1119),
.B1(n_1133),
.B2(n_1128),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1148),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_1067),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1082),
.B(n_1107),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1055),
.A2(n_1112),
.B(n_1116),
.C(n_1094),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1095),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1109),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1095),
.B(n_1164),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_SL g1257 ( 
.A(n_1095),
.Y(n_1257)
);

NOR3xp33_ASAP7_75t_L g1258 ( 
.A(n_1106),
.B(n_1096),
.C(n_1059),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1164),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1098),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_1066),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1064),
.B(n_1074),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1087),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1087),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1087),
.B(n_1170),
.Y(n_1265)
);

AOI221x1_ASAP7_75t_L g1266 ( 
.A1(n_1172),
.A2(n_1179),
.B1(n_1146),
.B2(n_1145),
.C(n_1163),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1076),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1150),
.B(n_1030),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1142),
.B(n_1153),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1150),
.B(n_1030),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1060),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1150),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1060),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1179),
.A2(n_902),
.B1(n_432),
.B2(n_434),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1076),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1068),
.Y(n_1280)
);

CKINVDCx6p67_ASAP7_75t_R g1281 ( 
.A(n_1076),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1155),
.A2(n_1180),
.B(n_1161),
.Y(n_1282)
);

AND2x2_ASAP7_75t_SL g1283 ( 
.A(n_1169),
.B(n_902),
.Y(n_1283)
);

INVx3_ASAP7_75t_SL g1284 ( 
.A(n_1171),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1155),
.A2(n_1180),
.B(n_1161),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1171),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1088),
.B(n_891),
.Y(n_1288)
);

OR2x6_ASAP7_75t_SL g1289 ( 
.A(n_1171),
.B(n_431),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1179),
.A2(n_903),
.B(n_1155),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1068),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1060),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1060),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1150),
.B(n_1030),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1155),
.A2(n_1180),
.B(n_1161),
.Y(n_1296)
);

INVx4_ASAP7_75t_SL g1297 ( 
.A(n_1160),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1150),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1142),
.B(n_1153),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1088),
.B(n_891),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1160),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1171),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1155),
.A2(n_1180),
.B(n_1161),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1104),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1155),
.B(n_1159),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1179),
.B(n_1140),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1150),
.Y(n_1310)
);

AOI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1142),
.A2(n_1156),
.B(n_1153),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1143),
.B(n_1154),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1155),
.B(n_1159),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1068),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1149),
.A2(n_903),
.B(n_1179),
.C(n_951),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1179),
.B(n_890),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1160),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1160),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1088),
.B(n_891),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1186),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1187),
.B(n_1271),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1215),
.Y(n_1322)
);

INVx4_ASAP7_75t_SL g1323 ( 
.A(n_1224),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1256),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1316),
.A2(n_1184),
.B(n_1315),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1268),
.B(n_1273),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1283),
.A2(n_1191),
.B1(n_1198),
.B2(n_1195),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1191),
.A2(n_1198),
.B1(n_1257),
.B2(n_1233),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1255),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1218),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1263),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1318),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1274),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1276),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1260),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1290),
.A2(n_1199),
.B1(n_1307),
.B2(n_1313),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1292),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1290),
.A2(n_1277),
.B1(n_1209),
.B2(n_1254),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1234),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1293),
.Y(n_1340)
);

CKINVDCx6p67_ASAP7_75t_R g1341 ( 
.A(n_1281),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1257),
.A2(n_1251),
.B1(n_1307),
.B2(n_1313),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1194),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1264),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1306),
.B(n_1183),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1234),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1259),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_1202),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1279),
.B(n_1286),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1258),
.A2(n_1247),
.B(n_1207),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1291),
.A2(n_1182),
.B1(n_1282),
.B2(n_1285),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1294),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1302),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1216),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1246),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1296),
.A2(n_1304),
.B1(n_1197),
.B2(n_1211),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1298),
.B(n_1305),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1227),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1272),
.B(n_1300),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1208),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1288),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1193),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1280),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1314),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1246),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1188),
.A2(n_1289),
.B1(n_1266),
.B2(n_1301),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1250),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1309),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_SL g1369 ( 
.A(n_1241),
.B(n_1231),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1217),
.A2(n_1221),
.B(n_1225),
.Y(n_1370)
);

AO21x1_ASAP7_75t_SL g1371 ( 
.A1(n_1200),
.A2(n_1205),
.B(n_1203),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1200),
.B(n_1238),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1238),
.B(n_1188),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1319),
.Y(n_1374)
);

INVx6_ASAP7_75t_L g1375 ( 
.A(n_1273),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1239),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1199),
.B(n_1201),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1228),
.Y(n_1378)
);

AO21x1_ASAP7_75t_L g1379 ( 
.A1(n_1229),
.A2(n_1237),
.B(n_1220),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1239),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1235),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1229),
.A2(n_1222),
.B1(n_1224),
.B2(n_1237),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1220),
.Y(n_1383)
);

AOI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1265),
.A2(n_1203),
.B(n_1262),
.Y(n_1384)
);

BUFx2_ASAP7_75t_SL g1385 ( 
.A(n_1287),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1204),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1249),
.A2(n_1253),
.B(n_1248),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1204),
.A2(n_1273),
.B1(n_1295),
.B2(n_1206),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1261),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1192),
.B(n_1299),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1224),
.A2(n_1231),
.B1(n_1294),
.B2(n_1241),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1317),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1248),
.A2(n_1249),
.B(n_1311),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1192),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1224),
.A2(n_1294),
.B1(n_1226),
.B2(n_1185),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1236),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1236),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1212),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1244),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1275),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1232),
.A2(n_1213),
.B1(n_1295),
.B2(n_1230),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1244),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1267),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1245),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1214),
.B(n_1312),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1245),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1275),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1310),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1252),
.A2(n_1308),
.B(n_1189),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1240),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1230),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1269),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1242),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1270),
.B(n_1189),
.Y(n_1415)
);

AO21x1_ASAP7_75t_L g1416 ( 
.A1(n_1252),
.A2(n_1243),
.B(n_1308),
.Y(n_1416)
);

BUFx2_ASAP7_75t_SL g1417 ( 
.A(n_1223),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1196),
.Y(n_1418)
);

CKINVDCx8_ASAP7_75t_R g1419 ( 
.A(n_1297),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1278),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1297),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1196),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1210),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1210),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1223),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1284),
.B(n_1219),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1190),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1190),
.A2(n_1283),
.B1(n_902),
.B2(n_742),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1303),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1283),
.A2(n_414),
.B1(n_449),
.B2(n_415),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1208),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1316),
.A2(n_1179),
.B1(n_903),
.B2(n_1153),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1219),
.Y(n_1433)
);

BUFx10_ASAP7_75t_L g1434 ( 
.A(n_1219),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1318),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1256),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1208),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1268),
.B(n_1273),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1256),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1316),
.A2(n_1090),
.B1(n_1179),
.B2(n_1146),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1283),
.A2(n_902),
.B1(n_742),
.B2(n_1179),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1187),
.B(n_1271),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1258),
.A2(n_1247),
.B(n_1207),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1316),
.A2(n_1179),
.B1(n_1120),
.B2(n_223),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1316),
.B(n_890),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1283),
.A2(n_902),
.B1(n_742),
.B2(n_1179),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1187),
.B(n_1271),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1260),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1316),
.B(n_890),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1319),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1186),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1186),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1202),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1186),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1256),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1348),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1331),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1445),
.B(n_1449),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1372),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1373),
.Y(n_1460)
);

BUFx5_ASAP7_75t_L g1461 ( 
.A(n_1383),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1389),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1343),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1384),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1343),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1373),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1335),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1381),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1398),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1389),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1381),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1360),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1345),
.B(n_1432),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1387),
.A2(n_1393),
.B(n_1379),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1384),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1320),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1332),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1377),
.B(n_1371),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_SL g1479 ( 
.A(n_1419),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1322),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1330),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1333),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1334),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1337),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1377),
.B(n_1371),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1340),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1325),
.A2(n_1440),
.B(n_1336),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1350),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1321),
.B(n_1349),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1453),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1324),
.B(n_1455),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1431),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1350),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1321),
.B(n_1349),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1436),
.B(n_1455),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1454),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1451),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1436),
.B(n_1439),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1389),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1439),
.B(n_1339),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1452),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1347),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1350),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1443),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1379),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1344),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1443),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1437),
.B(n_1362),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1335),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1352),
.B(n_1326),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1369),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1430),
.A2(n_1446),
.B1(n_1441),
.B2(n_1327),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1369),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1357),
.B(n_1442),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1410),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1339),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1359),
.B(n_1453),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1346),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1346),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1357),
.B(n_1442),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1443),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1447),
.B(n_1368),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1386),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1366),
.A2(n_1329),
.B(n_1388),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1394),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1400),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1447),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1356),
.B(n_1450),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1363),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1400),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1407),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1335),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1364),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1351),
.A2(n_1416),
.B(n_1409),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1358),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1409),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1407),
.B(n_1382),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1378),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1448),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1332),
.Y(n_1540)
);

AND2x4_ASAP7_75t_SL g1541 ( 
.A(n_1352),
.B(n_1326),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1326),
.B(n_1438),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1370),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1353),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1354),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1353),
.B(n_1412),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1361),
.B(n_1374),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1396),
.A2(n_1404),
.B(n_1397),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1392),
.B(n_1412),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1435),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1355),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1399),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1355),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1391),
.B(n_1402),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1406),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1448),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1365),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1448),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1414),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1428),
.A2(n_1338),
.B1(n_1328),
.B2(n_1342),
.Y(n_1560)
);

INVx11_ASAP7_75t_L g1561 ( 
.A(n_1341),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1458),
.B(n_1385),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1473),
.B(n_1460),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1517),
.B(n_1426),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1460),
.B(n_1435),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1457),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1457),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1548),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1478),
.B(n_1425),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1478),
.B(n_1485),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1485),
.B(n_1438),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1466),
.B(n_1367),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1476),
.Y(n_1573)
);

OAI211xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1487),
.A2(n_1423),
.B(n_1429),
.C(n_1427),
.Y(n_1574)
);

INVx5_ASAP7_75t_L g1575 ( 
.A(n_1515),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1476),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1510),
.B(n_1323),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1480),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1468),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1480),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1491),
.B(n_1495),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1481),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1491),
.B(n_1438),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1495),
.B(n_1411),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1481),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1505),
.B(n_1444),
.C(n_1401),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1466),
.B(n_1413),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1472),
.B(n_1417),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1492),
.B(n_1422),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1469),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1459),
.B(n_1390),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1502),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1498),
.B(n_1408),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1482),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1482),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1510),
.B(n_1323),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1483),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1514),
.B(n_1408),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1514),
.B(n_1405),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1459),
.B(n_1405),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1483),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1512),
.A2(n_1395),
.B1(n_1419),
.B2(n_1418),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1484),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1560),
.A2(n_1528),
.B1(n_1505),
.B2(n_1556),
.C(n_1468),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1484),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1486),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1471),
.B(n_1522),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1467),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1524),
.A2(n_1554),
.B1(n_1506),
.B2(n_1545),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1527),
.A2(n_1418),
.B1(n_1422),
.B2(n_1424),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1511),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1535),
.B(n_1376),
.Y(n_1613)
);

NOR2x1_ASAP7_75t_SL g1614 ( 
.A(n_1542),
.B(n_1418),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1464),
.B(n_1424),
.Y(n_1615)
);

NAND2xp33_ASAP7_75t_L g1616 ( 
.A(n_1461),
.B(n_1418),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1502),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1531),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1456),
.B(n_1426),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1523),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1531),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1529),
.B(n_1533),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1462),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1496),
.B(n_1415),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1496),
.B(n_1415),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1497),
.B(n_1501),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1563),
.B(n_1620),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1587),
.A2(n_1537),
.B1(n_1479),
.B2(n_1513),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1591),
.B(n_1513),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1608),
.B(n_1538),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1581),
.B(n_1470),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1605),
.B(n_1521),
.C(n_1506),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1574),
.B(n_1583),
.C(n_1612),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1622),
.B(n_1508),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1626),
.B(n_1508),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1493),
.C(n_1488),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1570),
.B(n_1499),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1587),
.A2(n_1501),
.B1(n_1497),
.B2(n_1507),
.C(n_1503),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1603),
.A2(n_1524),
.B1(n_1537),
.B2(n_1461),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1570),
.B(n_1461),
.Y(n_1640)
);

OAI221xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1610),
.A2(n_1549),
.B1(n_1554),
.B2(n_1494),
.C(n_1489),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1593),
.B(n_1617),
.C(n_1590),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1601),
.B(n_1463),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1463),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1465),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1600),
.B(n_1465),
.Y(n_1646)
);

NOR3xp33_ASAP7_75t_L g1647 ( 
.A(n_1589),
.B(n_1488),
.C(n_1493),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1619),
.B(n_1561),
.C(n_1543),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1562),
.A2(n_1520),
.B1(n_1565),
.B2(n_1564),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1565),
.B(n_1546),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1572),
.A2(n_1532),
.B1(n_1539),
.B2(n_1509),
.C(n_1558),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1569),
.B(n_1477),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1584),
.B(n_1461),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1584),
.B(n_1461),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1569),
.B(n_1461),
.Y(n_1655)
);

OAI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1579),
.A2(n_1488),
.B(n_1493),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1568),
.B(n_1550),
.C(n_1540),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1624),
.B(n_1552),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1577),
.B(n_1490),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1624),
.B(n_1555),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1625),
.B(n_1474),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1474),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1568),
.B(n_1475),
.C(n_1464),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1618),
.B(n_1474),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1618),
.B(n_1621),
.C(n_1534),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1573),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1573),
.B(n_1548),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1594),
.B(n_1461),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1576),
.B(n_1548),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1576),
.B(n_1461),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1578),
.B(n_1547),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1578),
.B(n_1509),
.Y(n_1672)
);

NAND4xp25_ASAP7_75t_L g1673 ( 
.A(n_1623),
.B(n_1539),
.C(n_1532),
.D(n_1509),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_L g1674 ( 
.A(n_1572),
.B(n_1534),
.C(n_1504),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1592),
.B(n_1534),
.C(n_1504),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1615),
.A2(n_1534),
.B(n_1551),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1577),
.A2(n_1524),
.B1(n_1375),
.B2(n_1559),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1592),
.B(n_1507),
.C(n_1503),
.Y(n_1678)
);

NAND4xp25_ASAP7_75t_L g1679 ( 
.A(n_1623),
.B(n_1532),
.C(n_1539),
.D(n_1558),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1588),
.A2(n_1558),
.B1(n_1421),
.B2(n_1429),
.C(n_1516),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1566),
.A2(n_1525),
.B1(n_1536),
.B2(n_1530),
.C(n_1526),
.Y(n_1681)
);

NOR3xp33_ASAP7_75t_L g1682 ( 
.A(n_1611),
.B(n_1475),
.C(n_1464),
.Y(n_1682)
);

AND2x2_ASAP7_75t_SL g1683 ( 
.A(n_1616),
.B(n_1500),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1567),
.A2(n_1421),
.B1(n_1519),
.B2(n_1516),
.C(n_1518),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1599),
.B(n_1571),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1580),
.B(n_1518),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1580),
.B(n_1519),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1582),
.B(n_1551),
.C(n_1553),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1582),
.B(n_1557),
.C(n_1553),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1599),
.B(n_1500),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1585),
.B(n_1500),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1586),
.B(n_1525),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1586),
.B(n_1557),
.C(n_1475),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1595),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1667),
.Y(n_1695)
);

INVx6_ASAP7_75t_L g1696 ( 
.A(n_1683),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1669),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1670),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1640),
.B(n_1614),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1664),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1640),
.B(n_1614),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1631),
.B(n_1691),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1686),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1687),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1692),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1674),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1666),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1671),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1688),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1685),
.B(n_1475),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1627),
.B(n_1595),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1642),
.B(n_1596),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1683),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1689),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1635),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1637),
.B(n_1655),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1693),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1629),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1672),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1634),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1630),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1658),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1628),
.A2(n_1597),
.B1(n_1577),
.B2(n_1541),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1653),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1660),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1678),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1665),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1647),
.B(n_1596),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1676),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1681),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1633),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1638),
.B(n_1598),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1654),
.B(n_1575),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1690),
.B(n_1668),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1682),
.B(n_1598),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1675),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1684),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1698),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1724),
.B(n_1652),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1696),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1724),
.B(n_1734),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1713),
.B(n_1636),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1709),
.B(n_1650),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1698),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1705),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1712),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1712),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1649),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1714),
.B(n_1652),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1705),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1703),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1703),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1714),
.B(n_1602),
.Y(n_1753)
);

NAND2x1_ASAP7_75t_SL g1754 ( 
.A(n_1736),
.B(n_1668),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1731),
.B(n_1602),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1731),
.B(n_1673),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1713),
.B(n_1679),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1696),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1717),
.B(n_1604),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1717),
.B(n_1604),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1724),
.B(n_1645),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1704),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1724),
.B(n_1646),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1696),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1737),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1718),
.B(n_1606),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1706),
.B(n_1643),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1734),
.B(n_1644),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1735),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1734),
.B(n_1609),
.Y(n_1771)
);

OAI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1727),
.A2(n_1639),
.B(n_1648),
.C(n_1651),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1711),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1737),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1732),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1706),
.B(n_1606),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1716),
.B(n_1609),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1711),
.Y(n_1778)
);

NOR2xp67_ASAP7_75t_L g1779 ( 
.A(n_1713),
.B(n_1736),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1699),
.B(n_1663),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1699),
.B(n_1597),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1706),
.B(n_1607),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1716),
.B(n_1609),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1708),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1770),
.B(n_1736),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1716),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1746),
.B(n_1730),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1776),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1753),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1741),
.B(n_1729),
.Y(n_1791)
);

AOI211xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1772),
.A2(n_1727),
.B(n_1659),
.C(n_1723),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1776),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1747),
.B(n_1730),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1783),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1748),
.B(n_1718),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1754),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1754),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1781),
.B(n_1720),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1755),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1782),
.B(n_1702),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1783),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1775),
.B(n_1743),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1775),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1749),
.B(n_1720),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1782),
.B(n_1702),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1760),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1743),
.B(n_1735),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1756),
.B(n_1597),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1782),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1738),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1757),
.A2(n_1729),
.B1(n_1696),
.B2(n_1723),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1773),
.B(n_1707),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1778),
.B(n_1707),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1766),
.A2(n_1726),
.B(n_1632),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1761),
.B(n_1721),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1739),
.B(n_1702),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1767),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1768),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1774),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1750),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1779),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1740),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1780),
.B(n_1699),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1740),
.A2(n_1726),
.B(n_1700),
.Y(n_1825)
);

NAND2x2_ASAP7_75t_L g1826 ( 
.A(n_1768),
.B(n_1561),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1751),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1758),
.B(n_1726),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1752),
.B(n_1721),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1785),
.B(n_1694),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1785),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1769),
.B(n_1722),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1791),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1792),
.A2(n_1728),
.B(n_1742),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1798),
.B(n_1739),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1817),
.B(n_1780),
.Y(n_1836)
);

AO22x1_ASAP7_75t_L g1837 ( 
.A1(n_1822),
.A2(n_1742),
.B1(n_1758),
.B2(n_1765),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1820),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1821),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1791),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1827),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1819),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1802),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1803),
.B(n_1808),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1804),
.B(n_1745),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1796),
.B(n_1808),
.Y(n_1846)
);

NOR2xp67_ASAP7_75t_L g1847 ( 
.A(n_1797),
.B(n_1758),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1803),
.B(n_1745),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1831),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1790),
.B(n_1759),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1802),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1786),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1791),
.Y(n_1853)
);

HB1xp67_ASAP7_75t_L g1854 ( 
.A(n_1823),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1817),
.B(n_1780),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1815),
.A2(n_1639),
.B1(n_1765),
.B2(n_1742),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1828),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1828),
.A2(n_1728),
.B(n_1759),
.Y(n_1858)
);

INVx4_ASAP7_75t_L g1859 ( 
.A(n_1809),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1800),
.B(n_1763),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1809),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1801),
.B(n_1769),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1801),
.B(n_1771),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1789),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1805),
.B(n_1816),
.Y(n_1865)
);

NOR3x1_ASAP7_75t_SL g1866 ( 
.A(n_1809),
.B(n_1403),
.C(n_1348),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1789),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1797),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1807),
.B(n_1763),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1788),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1793),
.Y(n_1871)
);

NAND3xp33_ASAP7_75t_L g1872 ( 
.A(n_1834),
.B(n_1825),
.C(n_1794),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1834),
.A2(n_1812),
.B(n_1799),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1839),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1838),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1839),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1841),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1844),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1841),
.Y(n_1879)
);

NAND3x1_ASAP7_75t_L g1880 ( 
.A(n_1866),
.B(n_1810),
.C(n_1806),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1843),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1857),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1844),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1870),
.A2(n_1852),
.B1(n_1846),
.B2(n_1856),
.C(n_1858),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1870),
.B(n_1818),
.Y(n_1885)
);

INVxp67_ASAP7_75t_L g1886 ( 
.A(n_1854),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1843),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1833),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1857),
.A2(n_1829),
.B(n_1814),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1870),
.A2(n_1793),
.B1(n_1795),
.B2(n_1765),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1851),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1862),
.B(n_1787),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1851),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1865),
.B(n_1832),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1849),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1859),
.B(n_1847),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1852),
.B(n_1787),
.Y(n_1897)
);

AOI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1858),
.A2(n_1795),
.B1(n_1641),
.B2(n_1813),
.C(n_1700),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1842),
.B(n_1830),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1842),
.B(n_1830),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1882),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1875),
.B(n_1865),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1875),
.B(n_1859),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1882),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1881),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1886),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1886),
.B(n_1859),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1878),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1892),
.B(n_1862),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1883),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1887),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1884),
.B(n_1833),
.Y(n_1912)
);

INVx3_ASAP7_75t_SL g1913 ( 
.A(n_1888),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1895),
.B(n_1833),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1891),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1893),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1889),
.B(n_1840),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1894),
.B(n_1840),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1897),
.B(n_1848),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1896),
.B(n_1840),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1896),
.B(n_1853),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1874),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1876),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1913),
.B(n_1885),
.Y(n_1924)
);

NAND4xp25_ASAP7_75t_L g1925 ( 
.A(n_1910),
.B(n_1872),
.C(n_1900),
.D(n_1899),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1912),
.A2(n_1873),
.B1(n_1880),
.B2(n_1898),
.Y(n_1926)
);

OAI211xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1917),
.A2(n_1868),
.B(n_1879),
.C(n_1877),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1913),
.A2(n_1868),
.B1(n_1835),
.B2(n_1890),
.Y(n_1928)
);

AOI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1901),
.A2(n_1868),
.B(n_1871),
.Y(n_1929)
);

A2O1A1Ixp33_ASAP7_75t_L g1930 ( 
.A1(n_1902),
.A2(n_1866),
.B(n_1861),
.C(n_1847),
.Y(n_1930)
);

OR3x1_ASAP7_75t_L g1931 ( 
.A(n_1907),
.B(n_1867),
.C(n_1864),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1913),
.A2(n_1837),
.B1(n_1871),
.B2(n_1867),
.C(n_1864),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1908),
.A2(n_1853),
.B1(n_1826),
.B2(n_1859),
.Y(n_1933)
);

AOI321xp33_ASAP7_75t_L g1934 ( 
.A1(n_1904),
.A2(n_1853),
.A3(n_1835),
.B1(n_1871),
.B2(n_1861),
.C(n_1845),
.Y(n_1934)
);

NAND3xp33_ASAP7_75t_L g1935 ( 
.A(n_1904),
.B(n_1837),
.C(n_1845),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1918),
.A2(n_1914),
.B1(n_1909),
.B2(n_1920),
.Y(n_1936)
);

OAI32xp33_ASAP7_75t_L g1937 ( 
.A1(n_1906),
.A2(n_1861),
.A3(n_1848),
.B1(n_1810),
.B2(n_1826),
.Y(n_1937)
);

INVx5_ASAP7_75t_L g1938 ( 
.A(n_1920),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1919),
.B(n_1918),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1934),
.B(n_1906),
.C(n_1903),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1938),
.B(n_1909),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_L g1942 ( 
.A(n_1924),
.B(n_1914),
.C(n_1921),
.Y(n_1942)
);

NOR2x1_ASAP7_75t_L g1943 ( 
.A(n_1931),
.B(n_1403),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1938),
.B(n_1921),
.Y(n_1944)
);

AOI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1926),
.A2(n_1923),
.B1(n_1916),
.B2(n_1915),
.C(n_1911),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1930),
.B(n_1938),
.Y(n_1946)
);

NOR3xp33_ASAP7_75t_L g1947 ( 
.A(n_1929),
.B(n_1923),
.C(n_1922),
.Y(n_1947)
);

NOR3xp33_ASAP7_75t_L g1948 ( 
.A(n_1925),
.B(n_1927),
.C(n_1935),
.Y(n_1948)
);

AO22x2_ASAP7_75t_L g1949 ( 
.A1(n_1939),
.A2(n_1911),
.B1(n_1915),
.B2(n_1916),
.Y(n_1949)
);

AOI211xp5_ASAP7_75t_L g1950 ( 
.A1(n_1932),
.A2(n_1919),
.B(n_1905),
.C(n_1855),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1936),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1937),
.A2(n_1860),
.B(n_1850),
.Y(n_1952)
);

OAI31xp33_ASAP7_75t_SL g1953 ( 
.A1(n_1933),
.A2(n_1836),
.A3(n_1855),
.B(n_1863),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1928),
.Y(n_1954)
);

NOR2x1_ASAP7_75t_L g1955 ( 
.A(n_1931),
.B(n_1420),
.Y(n_1955)
);

NAND4xp25_ASAP7_75t_L g1956 ( 
.A(n_1948),
.B(n_1836),
.C(n_1824),
.D(n_1863),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1940),
.A2(n_1869),
.B(n_1860),
.C(n_1850),
.Y(n_1957)
);

OAI21xp33_ASAP7_75t_L g1958 ( 
.A1(n_1953),
.A2(n_1869),
.B(n_1824),
.Y(n_1958)
);

AOI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1945),
.A2(n_1811),
.B1(n_1810),
.B2(n_1695),
.C(n_1697),
.Y(n_1959)
);

AOI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1949),
.A2(n_1811),
.B1(n_1695),
.B2(n_1697),
.C(n_1824),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1943),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1944),
.B(n_1420),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1941),
.B(n_1806),
.Y(n_1963)
);

NOR3x1_ASAP7_75t_L g1964 ( 
.A(n_1946),
.B(n_1951),
.C(n_1954),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_L g1965 ( 
.A(n_1955),
.B(n_1433),
.Y(n_1965)
);

INVxp67_ASAP7_75t_SL g1966 ( 
.A(n_1964),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1961),
.A2(n_1942),
.B1(n_1949),
.B2(n_1947),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1963),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1962),
.A2(n_1950),
.B1(n_1952),
.B2(n_1490),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1965),
.Y(n_1970)
);

AO22x2_ASAP7_75t_L g1971 ( 
.A1(n_1957),
.A2(n_1744),
.B1(n_1738),
.B2(n_1697),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1958),
.A2(n_1696),
.B1(n_1744),
.B2(n_1433),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1956),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1967),
.A2(n_1959),
.B(n_1960),
.Y(n_1974)
);

AOI221xp5_ASAP7_75t_SL g1975 ( 
.A1(n_1966),
.A2(n_1771),
.B1(n_1784),
.B2(n_1777),
.C(n_1764),
.Y(n_1975)
);

NOR3x1_ASAP7_75t_L g1976 ( 
.A(n_1970),
.B(n_1434),
.C(n_1433),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1969),
.B(n_1762),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1972),
.A2(n_1694),
.B1(n_1657),
.B2(n_1698),
.C(n_1680),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1968),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1973),
.B(n_1777),
.Y(n_1980)
);

XOR2xp5_ASAP7_75t_L g1981 ( 
.A(n_1980),
.B(n_1971),
.Y(n_1981)
);

XOR2xp5_ASAP7_75t_L g1982 ( 
.A(n_1979),
.B(n_1434),
.Y(n_1982)
);

AOI31xp33_ASAP7_75t_L g1983 ( 
.A1(n_1975),
.A2(n_1434),
.A3(n_1784),
.B(n_1762),
.Y(n_1983)
);

XNOR2xp5_ASAP7_75t_L g1984 ( 
.A(n_1982),
.B(n_1977),
.Y(n_1984)
);

NAND4xp25_ASAP7_75t_SL g1985 ( 
.A(n_1984),
.B(n_1976),
.C(n_1981),
.D(n_1983),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1974),
.B1(n_1978),
.B2(n_1708),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1985),
.A2(n_1418),
.B1(n_1725),
.B2(n_1722),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1986),
.A2(n_1764),
.B(n_1725),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1987),
.A2(n_1715),
.B(n_1719),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1988),
.Y(n_1990)
);

AOI21xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1989),
.A2(n_1380),
.B(n_1376),
.Y(n_1991)
);

AO21x2_ASAP7_75t_L g1992 ( 
.A1(n_1990),
.A2(n_1991),
.B(n_1715),
.Y(n_1992)
);

AOI322xp5_ASAP7_75t_L g1993 ( 
.A1(n_1992),
.A2(n_1710),
.A3(n_1719),
.B1(n_1677),
.B2(n_1733),
.C1(n_1656),
.C2(n_1701),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1993),
.A2(n_1710),
.B1(n_1733),
.B2(n_1424),
.C(n_1699),
.Y(n_1994)
);

AOI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1380),
.B(n_1701),
.C(n_1699),
.Y(n_1995)
);


endmodule