module real_aes_10929_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_402;
wire n_733;
wire n_602;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1699;
wire n_730;
wire n_1023;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_1772;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1679;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_0), .A2(n_391), .B1(n_1056), .B2(n_1058), .C(n_1063), .Y(n_1055) );
AOI21xp33_ASAP7_75t_L g1094 ( .A1(n_0), .A2(n_1095), .B(n_1096), .Y(n_1094) );
INVxp67_ASAP7_75t_L g399 ( .A(n_1), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_1), .A2(n_184), .B1(n_461), .B2(n_490), .C(n_495), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g1117 ( .A1(n_2), .A2(n_682), .B1(n_869), .B2(n_1118), .C(n_1123), .Y(n_1117) );
INVx1_ASAP7_75t_L g1137 ( .A(n_2), .Y(n_1137) );
XNOR2x2_ASAP7_75t_L g847 ( .A(n_3), .B(n_848), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g1430 ( .A1(n_3), .A2(n_301), .B1(n_1404), .B2(n_1412), .Y(n_1430) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_4), .A2(n_72), .B1(n_911), .B2(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1021 ( .A(n_4), .Y(n_1021) );
INVxp33_ASAP7_75t_L g940 ( .A(n_5), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_5), .A2(n_92), .B1(n_975), .B2(n_976), .C(n_977), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_6), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g340 ( .A1(n_7), .A2(n_238), .B1(n_341), .B2(n_352), .C(n_359), .Y(n_340) );
INVx1_ASAP7_75t_L g476 ( .A(n_7), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_8), .A2(n_103), .B1(n_355), .B2(n_695), .C(n_1018), .Y(n_1115) );
INVx1_ASAP7_75t_L g1142 ( .A(n_8), .Y(n_1142) );
INVx1_ASAP7_75t_L g956 ( .A(n_9), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1701 ( .A1(n_10), .A2(n_172), .B1(n_463), .B2(n_795), .Y(n_1701) );
OAI22xp5_ASAP7_75t_L g1718 ( .A1(n_10), .A2(n_172), .B1(n_1719), .B2(n_1721), .Y(n_1718) );
OAI221xp5_ASAP7_75t_L g1068 ( .A1(n_11), .A2(n_177), .B1(n_376), .B2(n_385), .C(n_388), .Y(n_1068) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_11), .Y(n_1101) );
AO22x1_ASAP7_75t_L g1106 ( .A1(n_12), .A2(n_1107), .B1(n_1144), .B2(n_1145), .Y(n_1106) );
INVx1_ASAP7_75t_L g1145 ( .A(n_12), .Y(n_1145) );
INVx1_ASAP7_75t_L g566 ( .A(n_13), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_14), .Y(n_420) );
INVx1_ASAP7_75t_L g1015 ( .A(n_15), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_15), .A2(n_82), .B1(n_713), .B2(n_1042), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g1753 ( .A(n_16), .Y(n_1753) );
AOI22xp33_ASAP7_75t_SL g1360 ( .A1(n_17), .A2(n_145), .B1(n_1361), .B2(n_1362), .Y(n_1360) );
AOI221xp5_ASAP7_75t_L g1385 ( .A1(n_17), .A2(n_234), .B1(n_900), .B2(n_1386), .C(n_1387), .Y(n_1385) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_18), .A2(n_151), .B1(n_640), .B2(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1284 ( .A(n_18), .Y(n_1284) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_19), .A2(n_109), .B1(n_374), .B2(n_383), .C(n_388), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_19), .A2(n_109), .B1(n_444), .B2(n_455), .Y(n_443) );
INVx1_ASAP7_75t_L g1003 ( .A(n_20), .Y(n_1003) );
OAI221xp5_ASAP7_75t_L g1026 ( .A1(n_20), .A2(n_869), .B1(n_881), .B2(n_1027), .C(n_1031), .Y(n_1026) );
OAI221xp5_ASAP7_75t_L g1779 ( .A1(n_21), .A2(n_76), .B1(n_455), .B2(n_1780), .C(n_1781), .Y(n_1779) );
INVx1_ASAP7_75t_L g1784 ( .A(n_21), .Y(n_1784) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_22), .A2(n_23), .B1(n_854), .B2(n_856), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_22), .A2(n_267), .B1(n_712), .B2(n_713), .Y(n_920) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_23), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g1431 ( .A1(n_24), .A2(n_271), .B1(n_1420), .B2(n_1426), .Y(n_1431) );
CKINVDCx16_ASAP7_75t_R g1457 ( .A(n_25), .Y(n_1457) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_26), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_27), .A2(n_91), .B1(n_492), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g698 ( .A(n_27), .Y(n_698) );
INVx1_ASAP7_75t_L g879 ( .A(n_28), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g890 ( .A1(n_28), .A2(n_170), .B1(n_891), .B2(n_893), .C(n_895), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_29), .A2(n_73), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
INVx1_ASAP7_75t_L g1092 ( .A(n_29), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_30), .A2(n_54), .B1(n_609), .B2(n_638), .Y(n_637) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_30), .A2(n_392), .B(n_676), .Y(n_675) );
INVxp33_ASAP7_75t_L g726 ( .A(n_31), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_31), .A2(n_90), .B1(n_634), .B2(n_756), .C(n_758), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g1164 ( .A1(n_32), .A2(n_94), .B1(n_374), .B2(n_384), .C(n_1165), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_32), .A2(n_94), .B1(n_579), .B2(n_800), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g802 ( .A1(n_33), .A2(n_225), .B1(n_496), .B2(n_768), .C(n_771), .Y(n_802) );
INVx1_ASAP7_75t_L g833 ( .A(n_33), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_34), .A2(n_162), .B1(n_738), .B2(n_739), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_34), .A2(n_162), .B1(n_776), .B2(n_778), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_35), .A2(n_40), .B1(n_688), .B2(n_743), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_35), .A2(n_103), .B1(n_713), .B2(n_1042), .Y(n_1143) );
INVx1_ASAP7_75t_L g318 ( .A(n_36), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g1677 ( .A1(n_37), .A2(n_223), .B1(n_1678), .B2(n_1679), .C(n_1680), .Y(n_1677) );
AOI22xp33_ASAP7_75t_L g1697 ( .A1(n_37), .A2(n_223), .B1(n_463), .B2(n_636), .Y(n_1697) );
INVx1_ASAP7_75t_L g928 ( .A(n_38), .Y(n_928) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_39), .Y(n_981) );
INVx1_ASAP7_75t_L g1141 ( .A(n_40), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_41), .A2(n_178), .B1(n_634), .B2(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1035 ( .A(n_41), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_42), .A2(n_157), .B1(n_1404), .B2(n_1412), .Y(n_1403) );
INVx1_ASAP7_75t_L g884 ( .A(n_43), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_44), .A2(n_203), .B1(n_1416), .B2(n_1445), .Y(n_1444) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_45), .A2(n_280), .B1(n_742), .B2(n_744), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_45), .A2(n_280), .B1(n_768), .B2(n_769), .C(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g1180 ( .A(n_46), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g1370 ( .A(n_47), .Y(n_1370) );
INVx1_ASAP7_75t_L g1302 ( .A(n_48), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_48), .A2(n_273), .B1(n_693), .B2(n_1325), .Y(n_1324) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_49), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g1116 ( .A1(n_50), .A2(n_100), .B1(n_700), .B2(n_702), .Y(n_1116) );
OAI22xp5_ASAP7_75t_SL g1130 ( .A1(n_50), .A2(n_100), .B1(n_648), .B2(n_654), .Y(n_1130) );
AO221x2_ASAP7_75t_L g1432 ( .A1(n_51), .A2(n_235), .B1(n_1420), .B2(n_1426), .C(n_1433), .Y(n_1432) );
XOR2x2_ASAP7_75t_L g1344 ( .A(n_52), .B(n_1345), .Y(n_1344) );
AOI22xp5_ASAP7_75t_L g1424 ( .A1(n_52), .A2(n_124), .B1(n_1404), .B2(n_1412), .Y(n_1424) );
CKINVDCx16_ASAP7_75t_R g1458 ( .A(n_53), .Y(n_1458) );
INVx1_ASAP7_75t_L g674 ( .A(n_54), .Y(n_674) );
INVx1_ASAP7_75t_L g605 ( .A(n_55), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_55), .A2(n_270), .B1(n_616), .B2(n_617), .C(n_619), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_56), .A2(n_122), .B1(n_739), .B2(n_742), .Y(n_745) );
INVxp67_ASAP7_75t_SL g753 ( .A(n_56), .Y(n_753) );
INVx1_ASAP7_75t_L g1204 ( .A(n_57), .Y(n_1204) );
AOI22xp5_ASAP7_75t_SL g1462 ( .A1(n_58), .A2(n_219), .B1(n_1416), .B2(n_1420), .Y(n_1462) );
INVxp33_ASAP7_75t_L g927 ( .A(n_59), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_59), .A2(n_113), .B1(n_964), .B2(n_967), .C(n_968), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_60), .Y(n_1357) );
INVxp33_ASAP7_75t_SL g1358 ( .A(n_61), .Y(n_1358) );
AOI221xp5_ASAP7_75t_L g1377 ( .A1(n_61), .A2(n_228), .B1(n_1378), .B2(n_1380), .C(n_1381), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_62), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_63), .A2(n_171), .B1(n_676), .B2(n_863), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_63), .A2(n_171), .B1(n_514), .B2(n_1080), .Y(n_1079) );
INVxp33_ASAP7_75t_L g939 ( .A(n_64), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_64), .A2(n_265), .B1(n_636), .B2(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g1699 ( .A(n_65), .Y(n_1699) );
OAI211xp5_ASAP7_75t_L g1653 ( .A1(n_66), .A2(n_1654), .B(n_1657), .C(n_1660), .Y(n_1653) );
INVx1_ASAP7_75t_L g1692 ( .A(n_66), .Y(n_1692) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_67), .A2(n_215), .B1(n_540), .B2(n_821), .C(n_934), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_67), .A2(n_215), .B1(n_455), .B2(n_962), .Y(n_961) );
CKINVDCx14_ASAP7_75t_R g1506 ( .A(n_68), .Y(n_1506) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_69), .A2(n_869), .B1(n_871), .B2(n_877), .C(n_881), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_69), .A2(n_221), .B1(n_499), .B2(n_900), .C(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g1128 ( .A(n_70), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1364 ( .A1(n_71), .A2(n_234), .B1(n_742), .B2(n_1365), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_71), .A2(n_145), .B1(n_1390), .B2(n_1391), .Y(n_1389) );
INVx1_ASAP7_75t_L g1024 ( .A(n_72), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_73), .A2(n_115), .B1(n_437), .B2(n_1090), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1761 ( .A1(n_74), .A2(n_285), .B1(n_526), .B2(n_1074), .Y(n_1761) );
INVx1_ASAP7_75t_L g1782 ( .A(n_74), .Y(n_1782) );
INVxp67_ASAP7_75t_SL g1352 ( .A(n_75), .Y(n_1352) );
OAI22xp33_ASAP7_75t_L g1374 ( .A1(n_75), .A2(n_274), .B1(n_1375), .B2(n_1376), .Y(n_1374) );
INVx1_ASAP7_75t_L g1785 ( .A(n_76), .Y(n_1785) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_77), .A2(n_112), .B1(n_738), .B2(n_744), .Y(n_746) );
INVxp67_ASAP7_75t_L g766 ( .A(n_77), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_78), .Y(n_797) );
INVx1_ASAP7_75t_L g1355 ( .A(n_79), .Y(n_1355) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_80), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_81), .A2(n_196), .B1(n_1404), .B2(n_1443), .Y(n_1442) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_82), .A2(n_304), .B1(n_1017), .B2(n_1018), .C(n_1019), .Y(n_1016) );
INVx1_ASAP7_75t_L g1006 ( .A(n_83), .Y(n_1006) );
OAI211xp5_ASAP7_75t_L g1011 ( .A1(n_83), .A2(n_851), .B(n_1012), .C(n_1020), .Y(n_1011) );
INVx1_ASAP7_75t_L g1160 ( .A(n_84), .Y(n_1160) );
OAI222xp33_ASAP7_75t_L g537 ( .A1(n_85), .A2(n_137), .B1(n_278), .B2(n_526), .C1(n_538), .C2(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g583 ( .A(n_85), .Y(n_583) );
OAI211xp5_ASAP7_75t_SL g1309 ( .A1(n_86), .A2(n_1078), .B(n_1310), .C(n_1313), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_86), .A2(n_181), .B1(n_1327), .B2(n_1331), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_87), .A2(n_211), .B1(n_462), .B2(n_643), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_87), .A2(n_211), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1214 ( .A1(n_88), .A2(n_218), .B1(n_794), .B2(n_1215), .C(n_1216), .Y(n_1214) );
INVx1_ASAP7_75t_L g1234 ( .A(n_88), .Y(n_1234) );
CKINVDCx14_ASAP7_75t_R g1434 ( .A(n_89), .Y(n_1434) );
INVxp33_ASAP7_75t_SL g730 ( .A(n_90), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_91), .A2(n_96), .B1(n_665), .B2(n_683), .Y(n_704) );
INVxp67_ASAP7_75t_L g943 ( .A(n_92), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_93), .A2(n_107), .B1(n_634), .B2(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g681 ( .A(n_93), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_95), .A2(n_303), .B1(n_800), .B2(n_1268), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1279 ( .A1(n_95), .A2(n_303), .B1(n_374), .B2(n_384), .C(n_821), .Y(n_1279) );
OAI222xp33_ASAP7_75t_L g706 ( .A1(n_96), .A2(n_129), .B1(n_210), .B2(n_527), .C1(n_707), .C2(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g349 ( .A(n_97), .Y(n_349) );
OR2x2_ASAP7_75t_L g381 ( .A(n_97), .B(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g394 ( .A(n_97), .Y(n_394) );
BUFx2_ASAP7_75t_L g529 ( .A(n_97), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_98), .A2(n_134), .B1(n_676), .B2(n_863), .Y(n_1062) );
INVx1_ASAP7_75t_L g1086 ( .A(n_98), .Y(n_1086) );
INVx1_ASAP7_75t_L g1122 ( .A(n_99), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_99), .A2(n_208), .B1(n_795), .B2(n_966), .Y(n_1135) );
INVx1_ASAP7_75t_L g656 ( .A(n_101), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_101), .A2(n_189), .B1(n_700), .B2(n_702), .C(n_703), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g1367 ( .A1(n_102), .A2(n_191), .B1(n_742), .B2(n_1365), .Y(n_1367) );
INVxp33_ASAP7_75t_SL g1394 ( .A(n_102), .Y(n_1394) );
INVx1_ASAP7_75t_L g1112 ( .A(n_104), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_104), .A2(n_250), .B1(n_436), .B2(n_795), .Y(n_1139) );
CKINVDCx5p33_ASAP7_75t_R g1218 ( .A(n_105), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g1667 ( .A1(n_106), .A2(n_232), .B1(n_1668), .B2(n_1670), .Y(n_1667) );
AOI221xp5_ASAP7_75t_L g1685 ( .A1(n_106), .A2(n_232), .B1(n_1686), .B2(n_1688), .C(n_1690), .Y(n_1685) );
INVx1_ASAP7_75t_L g679 ( .A(n_107), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g1258 ( .A1(n_108), .A2(n_183), .B1(n_595), .B2(n_597), .C(n_771), .Y(n_1258) );
INVxp67_ASAP7_75t_SL g1288 ( .A(n_108), .Y(n_1288) );
AOI22xp33_ASAP7_75t_SL g1368 ( .A1(n_110), .A2(n_246), .B1(n_1361), .B2(n_1362), .Y(n_1368) );
INVxp33_ASAP7_75t_L g1393 ( .A(n_110), .Y(n_1393) );
INVxp33_ASAP7_75t_L g1159 ( .A(n_111), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1191 ( .A1(n_111), .A2(n_311), .B1(n_794), .B2(n_1192), .C(n_1193), .Y(n_1191) );
INVxp33_ASAP7_75t_L g780 ( .A(n_112), .Y(n_780) );
INVxp33_ASAP7_75t_L g931 ( .A(n_113), .Y(n_931) );
INVx1_ASAP7_75t_L g1681 ( .A(n_114), .Y(n_1681) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_115), .A2(n_131), .B1(n_526), .B2(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g729 ( .A(n_116), .Y(n_729) );
INVx1_ASAP7_75t_L g360 ( .A(n_117), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_118), .A2(n_154), .B1(n_500), .B2(n_771), .C(n_972), .Y(n_1263) );
INVx1_ASAP7_75t_L g1277 ( .A(n_118), .Y(n_1277) );
INVx1_ASAP7_75t_L g984 ( .A(n_119), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_120), .Y(n_1225) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_121), .Y(n_808) );
INVxp33_ASAP7_75t_L g781 ( .A(n_122), .Y(n_781) );
INVx1_ASAP7_75t_L g1666 ( .A(n_123), .Y(n_1666) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_125), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1312 ( .A(n_126), .Y(n_1312) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_127), .A2(n_240), .B1(n_595), .B2(n_1199), .C(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1241 ( .A(n_127), .Y(n_1241) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_128), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_129), .A2(n_255), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_690) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_130), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g754 ( .A1(n_130), .A2(n_167), .B1(n_444), .B2(n_455), .Y(n_754) );
INVx1_ASAP7_75t_L g1098 ( .A(n_131), .Y(n_1098) );
INVx1_ASAP7_75t_L g1257 ( .A(n_132), .Y(n_1257) );
XNOR2xp5_ASAP7_75t_L g1206 ( .A(n_133), .B(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1083 ( .A(n_134), .Y(n_1083) );
AOI21xp33_ASAP7_75t_L g1307 ( .A1(n_135), .A2(n_496), .B(n_966), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_135), .A2(n_166), .B1(n_1327), .B2(n_1329), .Y(n_1326) );
INVxp33_ASAP7_75t_L g1168 ( .A(n_136), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_136), .A2(n_148), .B1(n_1201), .B2(n_1202), .Y(n_1200) );
INVx1_ASAP7_75t_L g602 ( .A(n_137), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g1751 ( .A(n_138), .Y(n_1751) );
AOI22xp5_ASAP7_75t_SL g1461 ( .A1(n_139), .A2(n_164), .B1(n_1404), .B2(n_1412), .Y(n_1461) );
OAI22xp33_ASAP7_75t_L g1318 ( .A1(n_140), .A2(n_181), .B1(n_514), .B2(n_516), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_140), .A2(n_253), .B1(n_693), .B2(n_1333), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_141), .Y(n_804) );
OAI22xp33_ASAP7_75t_SL g1212 ( .A1(n_142), .A2(n_289), .B1(n_579), .B2(n_1213), .Y(n_1212) );
OAI221xp5_ASAP7_75t_L g1235 ( .A1(n_142), .A2(n_289), .B1(n_374), .B2(n_384), .C(n_1165), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1311 ( .A(n_143), .Y(n_1311) );
INVx1_ASAP7_75t_L g874 ( .A(n_144), .Y(n_874) );
INVx1_ASAP7_75t_L g1408 ( .A(n_146), .Y(n_1408) );
AOI221xp5_ASAP7_75t_L g858 ( .A1(n_147), .A2(n_267), .B1(n_695), .B2(n_859), .C(n_861), .Y(n_858) );
INVxp67_ASAP7_75t_SL g919 ( .A(n_147), .Y(n_919) );
INVxp67_ASAP7_75t_SL g1175 ( .A(n_148), .Y(n_1175) );
INVx1_ASAP7_75t_L g1747 ( .A(n_149), .Y(n_1747) );
AOI22xp33_ASAP7_75t_SL g1775 ( .A1(n_149), .A2(n_282), .B1(n_795), .B2(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g930 ( .A(n_150), .Y(n_930) );
INVx1_ASAP7_75t_L g1289 ( .A(n_151), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_152), .A2(n_1249), .B1(n_1293), .B2(n_1294), .Y(n_1248) );
INVx1_ASAP7_75t_L g1294 ( .A(n_152), .Y(n_1294) );
INVx1_ASAP7_75t_L g1183 ( .A(n_153), .Y(n_1183) );
INVx1_ASAP7_75t_L g1275 ( .A(n_154), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1220 ( .A(n_155), .Y(n_1220) );
CKINVDCx16_ASAP7_75t_R g1454 ( .A(n_156), .Y(n_1454) );
INVx1_ASAP7_75t_L g1154 ( .A(n_157), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_158), .A2(n_198), .B1(n_1265), .B2(n_1266), .Y(n_1264) );
INVx1_ASAP7_75t_L g1274 ( .A(n_158), .Y(n_1274) );
INVx1_ASAP7_75t_L g1409 ( .A(n_159), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_159), .B(n_1407), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_160), .A2(n_185), .B1(n_587), .B2(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g813 ( .A(n_160), .Y(n_813) );
INVx1_ASAP7_75t_L g552 ( .A(n_161), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_163), .Y(n_1217) );
INVx2_ASAP7_75t_L g330 ( .A(n_165), .Y(n_330) );
INVx1_ASAP7_75t_L g1304 ( .A(n_166), .Y(n_1304) );
INVxp67_ASAP7_75t_SL g724 ( .A(n_167), .Y(n_724) );
INVxp67_ASAP7_75t_L g556 ( .A(n_168), .Y(n_556) );
OAI222xp33_ASAP7_75t_L g585 ( .A1(n_168), .A2(n_175), .B1(n_261), .B2(n_586), .C1(n_588), .C2(n_590), .Y(n_585) );
INVx1_ASAP7_75t_L g1227 ( .A(n_169), .Y(n_1227) );
AOI21xp33_ASAP7_75t_L g880 ( .A1(n_170), .A2(n_392), .B(n_859), .Y(n_880) );
BUFx3_ASAP7_75t_L g439 ( .A(n_173), .Y(n_439) );
INVx1_ASAP7_75t_L g469 ( .A(n_173), .Y(n_469) );
XNOR2x2_ASAP7_75t_L g337 ( .A(n_174), .B(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_L g564 ( .A(n_175), .Y(n_564) );
INVxp67_ASAP7_75t_L g413 ( .A(n_176), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_176), .A2(n_244), .B1(n_499), .B2(n_503), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_177), .Y(n_1102) );
INVx1_ASAP7_75t_L g1032 ( .A(n_178), .Y(n_1032) );
INVx1_ASAP7_75t_L g1742 ( .A(n_179), .Y(n_1742) );
AOI21xp33_ASAP7_75t_L g1777 ( .A1(n_179), .A2(n_436), .B(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g950 ( .A(n_180), .Y(n_950) );
INVx1_ASAP7_75t_L g876 ( .A(n_182), .Y(n_876) );
INVxp67_ASAP7_75t_SL g1285 ( .A(n_183), .Y(n_1285) );
INVxp67_ASAP7_75t_L g407 ( .A(n_184), .Y(n_407) );
INVx1_ASAP7_75t_L g817 ( .A(n_185), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g1644 ( .A1(n_186), .A2(n_264), .B1(n_1645), .B2(n_1649), .Y(n_1644) );
INVx1_ASAP7_75t_L g1711 ( .A(n_186), .Y(n_1711) );
INVx1_ASAP7_75t_L g442 ( .A(n_187), .Y(n_442) );
INVx1_ASAP7_75t_L g481 ( .A(n_187), .Y(n_481) );
INVx1_ASAP7_75t_L g1254 ( .A(n_188), .Y(n_1254) );
INVx1_ASAP7_75t_L g652 ( .A(n_189), .Y(n_652) );
INVx1_ASAP7_75t_L g727 ( .A(n_190), .Y(n_727) );
INVxp67_ASAP7_75t_SL g1373 ( .A(n_191), .Y(n_1373) );
XNOR2xp5_ASAP7_75t_L g534 ( .A(n_192), .B(n_535), .Y(n_534) );
INVxp67_ASAP7_75t_SL g1174 ( .A(n_193), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_193), .A2(n_268), .B1(n_768), .B2(n_1197), .C(n_1199), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_194), .Y(n_806) );
INVxp67_ASAP7_75t_L g543 ( .A(n_195), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_195), .A2(n_286), .B1(n_595), .B2(n_596), .C(n_597), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g1504 ( .A(n_197), .Y(n_1504) );
INVx1_ASAP7_75t_L g1278 ( .A(n_198), .Y(n_1278) );
CKINVDCx5p33_ASAP7_75t_R g1750 ( .A(n_199), .Y(n_1750) );
OA22x2_ASAP7_75t_L g786 ( .A1(n_200), .A2(n_787), .B1(n_843), .B2(n_844), .Y(n_786) );
INVx1_ASAP7_75t_L g844 ( .A(n_200), .Y(n_844) );
XOR2xp5_ASAP7_75t_L g1052 ( .A(n_201), .B(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g922 ( .A(n_202), .Y(n_922) );
CKINVDCx14_ASAP7_75t_R g1436 ( .A(n_204), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1731 ( .A1(n_204), .A2(n_1732), .B1(n_1736), .B2(n_1786), .Y(n_1731) );
INVx1_ASAP7_75t_L g1664 ( .A(n_205), .Y(n_1664) );
XNOR2xp5_ASAP7_75t_L g625 ( .A(n_206), .B(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_207), .A2(n_258), .B1(n_436), .B2(n_795), .Y(n_1316) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_207), .A2(n_306), .B1(n_1072), .B2(n_1074), .Y(n_1339) );
INVx1_ASAP7_75t_L g1120 ( .A(n_208), .Y(n_1120) );
INVx1_ASAP7_75t_L g1014 ( .A(n_209), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_209), .A2(n_304), .B1(n_707), .B2(n_710), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_210), .A2(n_300), .B1(n_687), .B2(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g957 ( .A(n_212), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1759 ( .A1(n_213), .A2(n_220), .B1(n_569), .B2(n_1760), .Y(n_1759) );
INVx1_ASAP7_75t_L g1769 ( .A(n_213), .Y(n_1769) );
OA332x1_ASAP7_75t_L g1740 ( .A1(n_214), .A2(n_391), .A3(n_1056), .B1(n_1741), .B2(n_1746), .B3(n_1749), .C1(n_1752), .C2(n_1757), .Y(n_1740) );
AOI21xp5_ASAP7_75t_L g1771 ( .A1(n_214), .A2(n_972), .B(n_1772), .Y(n_1771) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_216), .A2(n_283), .B1(n_700), .B2(n_702), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_216), .A2(n_283), .B1(n_909), .B2(n_911), .C(n_912), .Y(n_908) );
INVx1_ASAP7_75t_L g1270 ( .A(n_217), .Y(n_1270) );
INVx1_ASAP7_75t_L g1231 ( .A(n_218), .Y(n_1231) );
AOI22xp33_ASAP7_75t_SL g1770 ( .A1(n_220), .A2(n_285), .B1(n_436), .B2(n_795), .Y(n_1770) );
OAI211xp5_ASAP7_75t_L g850 ( .A1(n_221), .A2(n_851), .B(n_852), .C(n_865), .Y(n_850) );
INVx1_ASAP7_75t_L g866 ( .A(n_222), .Y(n_866) );
INVx1_ASAP7_75t_L g1683 ( .A(n_224), .Y(n_1683) );
INVx1_ASAP7_75t_L g828 ( .A(n_225), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_226), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_227), .A2(n_230), .B1(n_799), .B2(n_800), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_227), .A2(n_230), .B1(n_384), .B2(n_820), .C(n_821), .Y(n_819) );
INVxp33_ASAP7_75t_SL g1354 ( .A(n_228), .Y(n_1354) );
INVx1_ASAP7_75t_L g581 ( .A(n_229), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_231), .A2(n_251), .B1(n_604), .B2(n_640), .Y(n_1223) );
INVx1_ASAP7_75t_L g1238 ( .A(n_231), .Y(n_1238) );
CKINVDCx5p33_ASAP7_75t_R g1125 ( .A(n_233), .Y(n_1125) );
INVx1_ASAP7_75t_L g867 ( .A(n_236), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_237), .A2(n_252), .B1(n_609), .B2(n_611), .C(n_771), .Y(n_792) );
INVx1_ASAP7_75t_L g814 ( .A(n_237), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_238), .A2(n_308), .B1(n_461), .B2(n_464), .C(n_470), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_239), .Y(n_782) );
INVx1_ASAP7_75t_L g1239 ( .A(n_240), .Y(n_1239) );
INVx1_ASAP7_75t_L g438 ( .A(n_241), .Y(n_438) );
BUFx3_ASAP7_75t_L g454 ( .A(n_241), .Y(n_454) );
INVx1_ASAP7_75t_L g1700 ( .A(n_242), .Y(n_1700) );
AO221x2_ASAP7_75t_L g1501 ( .A1(n_243), .A2(n_295), .B1(n_1445), .B2(n_1502), .C(n_1503), .Y(n_1501) );
INVxp67_ASAP7_75t_L g396 ( .A(n_244), .Y(n_396) );
AOI21xp33_ASAP7_75t_L g1317 ( .A1(n_245), .A2(n_500), .B(n_972), .Y(n_1317) );
INVx1_ASAP7_75t_L g1337 ( .A(n_245), .Y(n_1337) );
INVxp67_ASAP7_75t_SL g1384 ( .A(n_246), .Y(n_1384) );
AOI22xp5_ASAP7_75t_L g1425 ( .A1(n_247), .A2(n_248), .B1(n_1420), .B2(n_1426), .Y(n_1425) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_249), .Y(n_326) );
AND2x2_ASAP7_75t_L g350 ( .A(n_249), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_249), .B(n_296), .Y(n_382) );
INVx1_ASAP7_75t_L g430 ( .A(n_249), .Y(n_430) );
INVx1_ASAP7_75t_L g1111 ( .A(n_250), .Y(n_1111) );
INVx1_ASAP7_75t_L g1242 ( .A(n_251), .Y(n_1242) );
INVx1_ASAP7_75t_L g816 ( .A(n_252), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_253), .A2(n_1080), .B1(n_1300), .B2(n_1305), .C(n_1308), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g1124 ( .A(n_254), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_255), .A2(n_300), .B1(n_712), .B2(n_713), .Y(n_711) );
OR2x2_ASAP7_75t_L g441 ( .A(n_256), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g449 ( .A(n_256), .Y(n_449) );
XNOR2xp5_ASAP7_75t_L g1737 ( .A(n_257), .B(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1338 ( .A(n_258), .Y(n_1338) );
INVx1_ASAP7_75t_L g545 ( .A(n_259), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_260), .A2(n_272), .B1(n_344), .B2(n_1065), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_260), .A2(n_272), .B1(n_516), .B2(n_1078), .Y(n_1077) );
INVxp67_ASAP7_75t_L g562 ( .A(n_261), .Y(n_562) );
INVx1_ASAP7_75t_L g1059 ( .A(n_262), .Y(n_1059) );
AOI21xp33_ASAP7_75t_L g1084 ( .A1(n_262), .A2(n_496), .B(n_595), .Y(n_1084) );
INVx1_ASAP7_75t_L g1185 ( .A(n_263), .Y(n_1185) );
INVx1_ASAP7_75t_L g1691 ( .A(n_264), .Y(n_1691) );
INVxp67_ASAP7_75t_L g946 ( .A(n_265), .Y(n_946) );
AOI22xp5_ASAP7_75t_SL g1415 ( .A1(n_266), .A2(n_269), .B1(n_1416), .B2(n_1420), .Y(n_1415) );
INVxp33_ASAP7_75t_SL g1170 ( .A(n_268), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_270), .A2(n_281), .B1(n_607), .B2(n_609), .C(n_611), .Y(n_606) );
INVx1_ASAP7_75t_L g1306 ( .A(n_273), .Y(n_1306) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_274), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_275), .A2(n_1296), .B1(n_1340), .B2(n_1341), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g1340 ( .A(n_275), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_276), .Y(n_521) );
INVx1_ASAP7_75t_L g1186 ( .A(n_277), .Y(n_1186) );
INVx1_ASAP7_75t_L g577 ( .A(n_278), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g1755 ( .A(n_279), .Y(n_1755) );
OAI332xp33_ASAP7_75t_L g541 ( .A1(n_281), .A2(n_391), .A3(n_542), .B1(n_548), .B2(n_555), .B3(n_563), .C1(n_567), .C2(n_569), .Y(n_541) );
INVx1_ASAP7_75t_L g1743 ( .A(n_282), .Y(n_1743) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_284), .A2(n_287), .B1(n_463), .B2(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g668 ( .A(n_284), .Y(n_668) );
INVx1_ASAP7_75t_L g549 ( .A(n_286), .Y(n_549) );
INVx1_ASAP7_75t_L g670 ( .A(n_287), .Y(n_670) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_288), .B(n_318), .Y(n_1411) );
AND3x2_ASAP7_75t_L g1419 ( .A(n_288), .B(n_318), .C(n_1408), .Y(n_1419) );
CKINVDCx5p33_ASAP7_75t_R g987 ( .A(n_290), .Y(n_987) );
INVx2_ASAP7_75t_L g331 ( .A(n_291), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_292), .A2(n_305), .B1(n_464), .B2(n_609), .Y(n_803) );
INVx1_ASAP7_75t_L g827 ( .A(n_292), .Y(n_827) );
OAI211xp5_ASAP7_75t_L g1109 ( .A1(n_293), .A2(n_851), .B(n_1110), .C(n_1113), .Y(n_1109) );
INVx1_ASAP7_75t_L g1138 ( .A(n_293), .Y(n_1138) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_294), .Y(n_997) );
INVx1_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
INVx2_ASAP7_75t_L g351 ( .A(n_296), .Y(n_351) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_297), .B(n_525), .Y(n_1297) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_298), .Y(n_993) );
INVx1_ASAP7_75t_L g1162 ( .A(n_299), .Y(n_1162) );
INVx1_ASAP7_75t_L g1262 ( .A(n_302), .Y(n_1262) );
INVx1_ASAP7_75t_L g835 ( .A(n_305), .Y(n_835) );
INVx1_ASAP7_75t_L g1314 ( .A(n_306), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g1748 ( .A(n_307), .Y(n_1748) );
INVxp33_ASAP7_75t_SL g366 ( .A(n_308), .Y(n_366) );
INVx1_ASAP7_75t_L g1253 ( .A(n_309), .Y(n_1253) );
INVx1_ASAP7_75t_L g954 ( .A(n_310), .Y(n_954) );
INVxp33_ASAP7_75t_L g1163 ( .A(n_311), .Y(n_1163) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_334), .B(n_1396), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1730 ( .A(n_316), .B(n_322), .Y(n_1730) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g1735 ( .A(n_317), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_317), .B(n_319), .Y(n_1789) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_319), .B(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x6_ASAP7_75t_L g1726 ( .A(n_324), .B(n_529), .Y(n_1726) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g736 ( .A(n_325), .B(n_333), .Y(n_736) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_393), .Y(n_392) );
INVx8_ASAP7_75t_L g1710 ( .A(n_327), .Y(n_1710) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
INVx1_ASAP7_75t_L g398 ( .A(n_328), .Y(n_398) );
OR2x2_ASAP7_75t_L g526 ( .A(n_328), .B(n_381), .Y(n_526) );
INVx2_ASAP7_75t_SL g554 ( .A(n_328), .Y(n_554) );
BUFx2_ASAP7_75t_L g826 ( .A(n_328), .Y(n_826) );
BUFx6f_ASAP7_75t_L g1246 ( .A(n_328), .Y(n_1246) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_328), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g1682 ( .A(n_328), .Y(n_1682) );
OR2x6_ASAP7_75t_L g1713 ( .A(n_328), .B(n_1714), .Y(n_1713) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g345 ( .A(n_330), .Y(n_345) );
INVx1_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
AND2x2_ASAP7_75t_L g365 ( .A(n_330), .B(n_331), .Y(n_365) );
AND2x4_ASAP7_75t_L g372 ( .A(n_330), .B(n_358), .Y(n_372) );
INVx1_ASAP7_75t_L g405 ( .A(n_330), .Y(n_405) );
INVx1_ASAP7_75t_L g347 ( .A(n_331), .Y(n_347) );
INVx2_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
INVx1_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
INVx1_ASAP7_75t_L g404 ( .A(n_331), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_331), .B(n_345), .Y(n_412) );
AND2x4_ASAP7_75t_L g1705 ( .A(n_332), .B(n_379), .Y(n_1705) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_1046), .B1(n_1047), .B2(n_1395), .Y(n_334) );
INVx1_ASAP7_75t_L g1395 ( .A(n_335), .Y(n_1395) );
AO22x2_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_784), .B1(n_1044), .B2(n_1045), .Y(n_335) );
INVx1_ASAP7_75t_L g1044 ( .A(n_336), .Y(n_1044) );
XNOR2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_531), .Y(n_336) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_431), .Y(n_338) );
NOR3xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_373), .C(n_389), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_342), .A2(n_353), .B1(n_726), .B2(n_727), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_342), .A2(n_362), .B1(n_1162), .B2(n_1163), .Y(n_1161) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_348), .Y(n_342) );
AND2x2_ASAP7_75t_L g539 ( .A(n_343), .B(n_348), .Y(n_539) );
AND2x2_ASAP7_75t_L g818 ( .A(n_343), .B(n_348), .Y(n_818) );
AND2x2_ASAP7_75t_L g932 ( .A(n_343), .B(n_348), .Y(n_932) );
INVx2_ASAP7_75t_SL g1689 ( .A(n_343), .Y(n_1689) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g669 ( .A(n_344), .B(n_350), .Y(n_669) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_344), .Y(n_687) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_344), .Y(n_743) );
INVx1_ASAP7_75t_L g855 ( .A(n_344), .Y(n_855) );
INVx1_ASAP7_75t_L g1328 ( .A(n_344), .Y(n_1328) );
BUFx2_ASAP7_75t_L g1678 ( .A(n_344), .Y(n_1678) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x6_ASAP7_75t_L g354 ( .A(n_348), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g362 ( .A(n_348), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g369 ( .A(n_348), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g570 ( .A(n_348), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_348), .B(n_676), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_348), .B(n_561), .Y(n_1075) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
OR2x2_ASAP7_75t_L g709 ( .A(n_349), .B(n_441), .Y(n_709) );
INVx2_ASAP7_75t_L g665 ( .A(n_350), .Y(n_665) );
AND2x4_ASAP7_75t_L g870 ( .A(n_350), .B(n_692), .Y(n_870) );
INVx1_ASAP7_75t_L g393 ( .A(n_351), .Y(n_393) );
INVx1_ASAP7_75t_L g429 ( .A(n_351), .Y(n_429) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_354), .A2(n_369), .B1(n_813), .B2(n_814), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_354), .A2(n_368), .B1(n_927), .B2(n_928), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_354), .A2(n_731), .B1(n_1159), .B2(n_1160), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_354), .A2(n_1217), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_354), .A2(n_1232), .B1(n_1354), .B2(n_1355), .Y(n_1353) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_355), .B(n_380), .Y(n_388) );
BUFx2_ASAP7_75t_L g1017 ( .A(n_355), .Y(n_1017) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_356), .Y(n_571) );
BUFx2_ASAP7_75t_L g623 ( .A(n_356), .Y(n_623) );
BUFx3_ASAP7_75t_L g694 ( .A(n_356), .Y(n_694) );
BUFx6f_ASAP7_75t_L g863 ( .A(n_356), .Y(n_863) );
AND2x4_ASAP7_75t_L g1716 ( .A(n_356), .B(n_1717), .Y(n_1716) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_366), .B2(n_367), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_360), .A2(n_471), .B1(n_476), .B2(n_477), .C(n_480), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_361), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g616 ( .A(n_362), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_362), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_362), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_362), .A2(n_818), .B1(n_1218), .B2(n_1234), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_362), .A2(n_539), .B1(n_1277), .B2(n_1278), .Y(n_1276) );
AOI221xp5_ASAP7_75t_L g1336 ( .A1(n_362), .A2(n_932), .B1(n_1337), .B2(n_1338), .C(n_1339), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_362), .A2(n_818), .B1(n_1357), .B2(n_1358), .Y(n_1356) );
INVx1_ASAP7_75t_L g860 ( .A(n_363), .Y(n_860) );
BUFx2_ASAP7_75t_L g1325 ( .A(n_363), .Y(n_1325) );
BUFx3_ASAP7_75t_L g1361 ( .A(n_363), .Y(n_1361) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g676 ( .A(n_364), .Y(n_676) );
INVx2_ASAP7_75t_L g705 ( .A(n_364), .Y(n_705) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_365), .Y(n_692) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g618 ( .A(n_369), .Y(n_618) );
BUFx2_ASAP7_75t_L g731 ( .A(n_369), .Y(n_731) );
BUFx2_ASAP7_75t_L g1232 ( .A(n_369), .Y(n_1232) );
BUFx3_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
INVx2_ASAP7_75t_L g875 ( .A(n_370), .Y(n_875) );
INVx1_ASAP7_75t_SL g1060 ( .A(n_370), .Y(n_1060) );
INVx1_ASAP7_75t_L g1121 ( .A(n_370), .Y(n_1121) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g561 ( .A(n_371), .Y(n_561) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_371), .Y(n_689) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_372), .Y(n_547) );
INVx1_ASAP7_75t_L g667 ( .A(n_372), .Y(n_667) );
INVx1_ASAP7_75t_L g1724 ( .A(n_372), .Y(n_1724) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_SL g934 ( .A(n_375), .Y(n_934) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_376), .Y(n_820) );
NAND2x1_ASAP7_75t_SL g376 ( .A(n_377), .B(n_380), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g700 ( .A(n_377), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_379), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_380), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g620 ( .A(n_380), .B(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_L g622 ( .A(n_380), .B(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g721 ( .A(n_380), .B(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g684 ( .A(n_382), .Y(n_684) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx4f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx4f_ASAP7_75t_L g540 ( .A(n_385), .Y(n_540) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x6_ASAP7_75t_L g702 ( .A(n_387), .B(n_683), .Y(n_702) );
BUFx3_ASAP7_75t_L g821 ( .A(n_388), .Y(n_821) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_388), .Y(n_1165) );
OAI33xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_395), .A3(n_406), .B1(n_416), .B2(n_419), .B3(n_424), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI33xp33_ASAP7_75t_L g822 ( .A1(n_391), .A2(n_424), .A3(n_823), .B1(n_829), .B2(n_836), .B3(n_840), .Y(n_822) );
INVx1_ASAP7_75t_L g937 ( .A(n_391), .Y(n_937) );
OAI33xp33_ASAP7_75t_L g1166 ( .A1(n_391), .A2(n_424), .A3(n_1167), .B1(n_1173), .B2(n_1178), .B3(n_1184), .Y(n_1166) );
OAI33xp33_ASAP7_75t_L g1236 ( .A1(n_391), .A2(n_424), .A3(n_1237), .B1(n_1240), .B2(n_1243), .B3(n_1245), .Y(n_1236) );
OAI33xp33_ASAP7_75t_L g1280 ( .A1(n_391), .A2(n_567), .A3(n_1281), .B1(n_1286), .B2(n_1290), .B3(n_1292), .Y(n_1280) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g1714 ( .A(n_393), .Y(n_1714) );
BUFx2_ASAP7_75t_L g520 ( .A(n_394), .Y(n_520) );
INVx2_ASAP7_75t_L g631 ( .A(n_394), .Y(n_631) );
OAI22xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B1(n_399), .B2(n_400), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_397), .A2(n_408), .B1(n_417), .B2(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g565 ( .A(n_398), .Y(n_565) );
OAI22xp5_ASAP7_75t_SL g563 ( .A1(n_400), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
OAI22xp33_ASAP7_75t_L g1184 ( .A1(n_400), .A2(n_1169), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g1028 ( .A(n_401), .Y(n_1028) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx3_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
BUFx3_ASAP7_75t_L g941 ( .A(n_402), .Y(n_941) );
OAI22xp33_ASAP7_75t_L g1749 ( .A1(n_402), .A2(n_1246), .B1(n_1750), .B2(n_1751), .Y(n_1749) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g551 ( .A(n_404), .B(n_405), .Y(n_551) );
INVx1_ASAP7_75t_L g723 ( .A(n_405), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_413), .B2(n_414), .Y(n_406) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g544 ( .A(n_410), .Y(n_544) );
INVx2_ASAP7_75t_L g1287 ( .A(n_410), .Y(n_1287) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g678 ( .A(n_411), .Y(n_678) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g559 ( .A(n_412), .Y(n_559) );
INVx1_ASAP7_75t_L g832 ( .A(n_412), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_414), .A2(n_420), .B1(n_421), .B2(n_423), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_414), .A2(n_950), .B1(n_951), .B2(n_954), .Y(n_949) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_415), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_417), .A2(n_420), .B1(n_513), .B2(n_515), .Y(n_512) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_418), .A2(n_434), .B(n_443), .C(n_460), .Y(n_433) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g823 ( .A1(n_422), .A2(n_824), .B1(n_827), .B2(n_828), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g1237 ( .A1(n_422), .A2(n_1169), .B1(n_1238), .B2(n_1239), .Y(n_1237) );
OAI22xp33_ASAP7_75t_L g1746 ( .A1(n_422), .A2(n_553), .B1(n_1747), .B2(n_1748), .Y(n_1746) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_423), .A2(n_483), .B1(n_489), .B2(n_498), .C(n_506), .Y(n_482) );
INVx1_ASAP7_75t_L g747 ( .A(n_424), .Y(n_747) );
OAI33xp33_ASAP7_75t_L g935 ( .A1(n_424), .A2(n_936), .A3(n_938), .B1(n_942), .B2(n_949), .B3(n_955), .Y(n_935) );
CKINVDCx8_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
INVx5_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx6_ASAP7_75t_L g568 ( .A(n_426), .Y(n_568) );
OR2x6_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_427), .B(n_446), .Y(n_651) );
INVx2_ASAP7_75t_L g696 ( .A(n_428), .Y(n_696) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g1708 ( .A(n_429), .Y(n_1708) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_517), .B1(n_521), .B2(n_522), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_482), .C(n_512), .Y(n_432) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_435), .A2(n_753), .B(n_754), .C(n_755), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_435), .A2(n_513), .B1(n_950), .B2(n_956), .Y(n_980) );
AOI211xp5_ASAP7_75t_SL g1189 ( .A1(n_435), .A2(n_1180), .B(n_1190), .C(n_1191), .Y(n_1189) );
AOI211xp5_ASAP7_75t_SL g1210 ( .A1(n_435), .A2(n_1211), .B(n_1212), .C(n_1214), .Y(n_1210) );
AOI211xp5_ASAP7_75t_L g1372 ( .A1(n_435), .A2(n_1373), .B(n_1374), .C(n_1377), .Y(n_1372) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_440), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g463 ( .A(n_437), .Y(n_463) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_437), .Y(n_587) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_437), .Y(n_595) );
INVx2_ASAP7_75t_SL g635 ( .A(n_437), .Y(n_635) );
BUFx2_ASAP7_75t_L g768 ( .A(n_437), .Y(n_768) );
BUFx6f_ASAP7_75t_L g966 ( .A(n_437), .Y(n_966) );
BUFx2_ASAP7_75t_L g975 ( .A(n_437), .Y(n_975) );
HB1xp67_ASAP7_75t_L g1215 ( .A(n_437), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1265 ( .A(n_437), .Y(n_1265) );
AND2x6_ASAP7_75t_L g1669 ( .A(n_437), .B(n_1647), .Y(n_1669) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
INVx2_ASAP7_75t_L g459 ( .A(n_439), .Y(n_459) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_454), .Y(n_488) );
AND2x4_ASAP7_75t_L g486 ( .A(n_440), .B(n_487), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_440), .A2(n_486), .B1(n_566), .B2(n_585), .C(n_591), .Y(n_584) );
AND2x2_ASAP7_75t_L g796 ( .A(n_440), .B(n_587), .Y(n_796) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g514 ( .A(n_441), .B(n_479), .Y(n_514) );
OR2x2_ASAP7_75t_L g516 ( .A(n_441), .B(n_467), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g1763 ( .A1(n_441), .A2(n_1764), .B(n_1765), .C(n_1766), .Y(n_1763) );
INVx1_ASAP7_75t_L g447 ( .A(n_442), .Y(n_447) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g962 ( .A(n_445), .Y(n_962) );
INVx2_ASAP7_75t_L g1375 ( .A(n_445), .Y(n_1375) );
INVx2_ASAP7_75t_SL g1780 ( .A(n_445), .Y(n_1780) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_450), .Y(n_445) );
AND2x2_ASAP7_75t_L g456 ( .A(n_446), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g510 ( .A(n_446), .Y(n_510) );
AND2x2_ASAP7_75t_L g530 ( .A(n_446), .B(n_502), .Y(n_530) );
AND2x4_ASAP7_75t_L g580 ( .A(n_446), .B(n_450), .Y(n_580) );
AND2x4_ASAP7_75t_L g582 ( .A(n_446), .B(n_457), .Y(n_582) );
BUFx2_ASAP7_75t_L g592 ( .A(n_446), .Y(n_592) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AND2x4_ASAP7_75t_L g480 ( .A(n_448), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g497 ( .A(n_449), .B(n_481), .Y(n_497) );
INVx1_ASAP7_75t_L g1648 ( .A(n_449), .Y(n_1648) );
HB1xp67_ASAP7_75t_L g1652 ( .A(n_449), .Y(n_1652) );
INVx1_ASAP7_75t_L g1673 ( .A(n_449), .Y(n_1673) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_450), .A2(n_457), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g649 ( .A(n_451), .Y(n_649) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g1663 ( .A(n_452), .Y(n_1663) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g502 ( .A(n_453), .B(n_459), .Y(n_502) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g468 ( .A(n_454), .B(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g655 ( .A(n_457), .Y(n_655) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x6_ASAP7_75t_L g1665 ( .A(n_458), .B(n_1648), .Y(n_1665) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g604 ( .A(n_465), .Y(n_604) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_466), .Y(n_1000) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g1090 ( .A(n_467), .Y(n_1090) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_468), .Y(n_505) );
INVx1_ASAP7_75t_L g644 ( .A(n_468), .Y(n_644) );
INVx1_ASAP7_75t_L g757 ( .A(n_468), .Y(n_757) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_468), .Y(n_795) );
INVx1_ASAP7_75t_L g474 ( .A(n_469), .Y(n_474) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g714 ( .A(n_473), .Y(n_714) );
INVx1_ASAP7_75t_L g761 ( .A(n_473), .Y(n_761) );
INVx1_ASAP7_75t_L g969 ( .A(n_473), .Y(n_969) );
INVx1_ASAP7_75t_L g996 ( .A(n_473), .Y(n_996) );
BUFx4f_ASAP7_75t_L g1134 ( .A(n_473), .Y(n_1134) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
OR2x2_ASAP7_75t_L g479 ( .A(n_474), .B(n_475), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_477), .A2(n_993), .B1(n_994), .B2(n_997), .C(n_998), .Y(n_992) );
OAI221xp5_ASAP7_75t_L g1695 ( .A1(n_477), .A2(n_1681), .B1(n_1683), .B2(n_1696), .C(n_1697), .Y(n_1695) );
OAI221xp5_ASAP7_75t_L g1698 ( .A1(n_477), .A2(n_1696), .B1(n_1699), .B2(n_1700), .C(n_1701), .Y(n_1698) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g708 ( .A(n_478), .Y(n_708) );
INVx2_ASAP7_75t_L g970 ( .A(n_478), .Y(n_970) );
INVx2_ASAP7_75t_L g1301 ( .A(n_478), .Y(n_1301) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g589 ( .A(n_479), .Y(n_589) );
BUFx2_ASAP7_75t_L g762 ( .A(n_479), .Y(n_762) );
INVx1_ASAP7_75t_L g1088 ( .A(n_479), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1645 ( .A(n_479), .B(n_1646), .Y(n_1645) );
INVx1_ASAP7_75t_L g611 ( .A(n_480), .Y(n_611) );
AND2x4_ASAP7_75t_L g645 ( .A(n_480), .B(n_529), .Y(n_645) );
AND2x4_ASAP7_75t_L g907 ( .A(n_480), .B(n_529), .Y(n_907) );
INVx2_ASAP7_75t_SL g972 ( .A(n_480), .Y(n_972) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_480), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_480), .A2(n_708), .B1(n_761), .B2(n_1160), .C(n_1162), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_480), .A2(n_708), .B1(n_761), .B2(n_1217), .C(n_1218), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_480), .Y(n_1382) );
INVx1_ASAP7_75t_L g1675 ( .A(n_481), .Y(n_1675) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g973 ( .A1(n_485), .A2(n_508), .B1(n_957), .B2(n_974), .C(n_978), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g1383 ( .A1(n_485), .A2(n_508), .B1(n_1384), .B2(n_1385), .C(n_1389), .Y(n_1383) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_486), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_486), .A2(n_591), .B1(n_802), .B2(n_803), .C(n_804), .Y(n_801) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_486), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_486), .Y(n_1195) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_486), .A2(n_591), .B1(n_1220), .B2(n_1221), .C(n_1223), .Y(n_1219) );
AND2x4_ASAP7_75t_L g591 ( .A(n_487), .B(n_592), .Y(n_591) );
BUFx4f_ASAP7_75t_L g596 ( .A(n_487), .Y(n_596) );
INVx1_ASAP7_75t_L g608 ( .A(n_487), .Y(n_608) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_487), .Y(n_638) );
INVx2_ASAP7_75t_SL g1198 ( .A(n_487), .Y(n_1198) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_488), .Y(n_494) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g771 ( .A(n_493), .Y(n_771) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_494), .Y(n_511) );
INVx1_ASAP7_75t_L g659 ( .A(n_494), .Y(n_659) );
BUFx6f_ASAP7_75t_L g1656 ( .A(n_494), .Y(n_1656) );
AND2x4_ASAP7_75t_L g1658 ( .A(n_494), .B(n_1659), .Y(n_1658) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g1388 ( .A(n_496), .Y(n_1388) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
BUFx3_ASAP7_75t_L g598 ( .A(n_497), .Y(n_598) );
INVx1_ASAP7_75t_L g632 ( .A(n_497), .Y(n_632) );
INVx2_ASAP7_75t_L g774 ( .A(n_497), .Y(n_774) );
INVx1_ASAP7_75t_L g1778 ( .A(n_497), .Y(n_1778) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g918 ( .A(n_500), .B(n_916), .Y(n_918) );
A2O1A1Ixp33_ASAP7_75t_L g1097 ( .A1(n_500), .A2(n_1098), .B(n_1099), .C(n_1103), .Y(n_1097) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g1390 ( .A(n_501), .Y(n_1390) );
INVx1_ASAP7_75t_L g1772 ( .A(n_501), .Y(n_1772) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx6_ASAP7_75t_L g610 ( .A(n_502), .Y(n_610) );
BUFx2_ASAP7_75t_L g777 ( .A(n_502), .Y(n_777) );
AND2x4_ASAP7_75t_L g1650 ( .A(n_502), .B(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI221xp5_ASAP7_75t_SL g593 ( .A1(n_504), .A2(n_545), .B1(n_552), .B2(n_588), .C(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g906 ( .A(n_504), .Y(n_906) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g590 ( .A(n_505), .Y(n_590) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_505), .Y(n_636) );
INVx1_ASAP7_75t_L g896 ( .A(n_505), .Y(n_896) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_505), .Y(n_1260) );
BUFx6f_ASAP7_75t_L g1391 ( .A(n_505), .Y(n_1391) );
AND2x6_ASAP7_75t_L g1671 ( .A(n_505), .B(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_508), .A2(n_765), .B1(n_766), .B2(n_767), .C(n_775), .Y(n_764) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_510), .B(n_655), .Y(n_1376) );
INVx1_ASAP7_75t_L g892 ( .A(n_511), .Y(n_892) );
BUFx6f_ASAP7_75t_L g976 ( .A(n_511), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_513), .A2(n_515), .B1(n_780), .B2(n_781), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_513), .A2(n_515), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_513), .A2(n_515), .B1(n_1183), .B2(n_1185), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_513), .A2(n_515), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_513), .A2(n_515), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_513), .A2(n_515), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
INVx6_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI211xp5_ASAP7_75t_L g960 ( .A1(n_515), .A2(n_954), .B(n_961), .C(n_963), .Y(n_960) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_SL g1039 ( .A(n_517), .Y(n_1039) );
INVx5_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g1108 ( .A1(n_518), .A2(n_1109), .B(n_1117), .Y(n_1108) );
BUFx8_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
AOI31xp33_ASAP7_75t_L g751 ( .A1(n_519), .A2(n_752), .A3(n_764), .B(n_779), .Y(n_751) );
INVx2_ASAP7_75t_L g1104 ( .A(n_519), .Y(n_1104) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g614 ( .A(n_520), .Y(n_614) );
AND2x4_ASAP7_75t_L g1674 ( .A(n_520), .B(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_524), .A2(n_614), .B1(n_959), .B2(n_981), .Y(n_958) );
AOI21xp5_ASAP7_75t_L g1369 ( .A1(n_524), .A2(n_1370), .B(n_1371), .Y(n_1369) );
INVx5_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g749 ( .A(n_525), .Y(n_749) );
INVx2_ASAP7_75t_SL g809 ( .A(n_525), .Y(n_809) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x6_ASAP7_75t_L g885 ( .A(n_528), .B(n_886), .Y(n_885) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_530), .B(n_1782), .Y(n_1781) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_716), .B2(n_783), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AO22x2_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_624), .B1(n_625), .B2(n_715), .Y(n_533) );
INVx1_ASAP7_75t_L g715 ( .A(n_534), .Y(n_715) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_572), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g1071 ( .A(n_539), .Y(n_1071) );
INVx1_ASAP7_75t_L g1760 ( .A(n_539), .Y(n_1760) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g1012 ( .A1(n_546), .A2(n_1013), .B1(n_1014), .B2(n_1015), .C(n_1016), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_546), .A2(n_1211), .B1(n_1226), .B2(n_1244), .Y(n_1243) );
INVx4_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_SL g1366 ( .A(n_547), .Y(n_1366) );
BUFx3_ASAP7_75t_L g1679 ( .A(n_547), .Y(n_1679) );
INVx2_ASAP7_75t_SL g1687 ( .A(n_547), .Y(n_1687) );
INVx2_ASAP7_75t_SL g1756 ( .A(n_547), .Y(n_1756) );
OAI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_552), .B2(n_553), .Y(n_548) );
OR2x6_ASAP7_75t_L g682 ( .A(n_550), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g842 ( .A(n_550), .Y(n_842) );
OR2x2_ASAP7_75t_L g881 ( .A(n_550), .B(n_683), .Y(n_881) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g673 ( .A(n_551), .Y(n_673) );
INVx2_ASAP7_75t_L g878 ( .A(n_551), .Y(n_878) );
BUFx2_ASAP7_75t_L g1172 ( .A(n_551), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_553), .A2(n_939), .B1(n_940), .B2(n_941), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g955 ( .A1(n_553), .A2(n_941), .B1(n_956), .B2(n_957), .Y(n_955) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_553), .A2(n_993), .B1(n_997), .B2(n_1028), .C(n_1029), .Y(n_1027) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_553), .A2(n_673), .B1(n_1124), .B2(n_1125), .C(n_1126), .Y(n_1123) );
OAI22xp33_ASAP7_75t_SL g1690 ( .A1(n_553), .A2(n_673), .B1(n_1691), .B2(n_1692), .Y(n_1690) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_560), .B2(n_562), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_557), .A2(n_1032), .B1(n_1033), .B2(n_1035), .Y(n_1031) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_559), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1719 ( .A(n_559), .B(n_1720), .Y(n_1719) );
INVx1_ASAP7_75t_L g1034 ( .A(n_560), .Y(n_1034) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g834 ( .A(n_561), .Y(n_834) );
INVx2_ASAP7_75t_L g839 ( .A(n_561), .Y(n_839) );
INVx2_ASAP7_75t_L g857 ( .A(n_561), .Y(n_857) );
HB1xp67_ASAP7_75t_L g1745 ( .A(n_561), .Y(n_1745) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI33xp33_ASAP7_75t_L g1359 ( .A1(n_568), .A2(n_733), .A3(n_1360), .B1(n_1364), .B2(n_1367), .B3(n_1368), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g1676 ( .A1(n_568), .A2(n_1677), .B1(n_1684), .B2(n_1685), .C(n_1693), .Y(n_1676) );
INVx1_ASAP7_75t_L g1757 ( .A(n_568), .Y(n_1757) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g1072 ( .A(n_570), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_570), .A2(n_1075), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
INVx2_ASAP7_75t_SL g1363 ( .A(n_571), .Y(n_1363) );
AOI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_612), .B(n_615), .Y(n_572) );
NAND4xp25_ASAP7_75t_SL g573 ( .A(n_574), .B(n_584), .C(n_593), .D(n_599), .Y(n_573) );
AOI222xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_577), .B1(n_578), .B2(n_581), .C1(n_582), .C2(n_583), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx4_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g799 ( .A(n_580), .Y(n_799) );
INVx1_ASAP7_75t_SL g1268 ( .A(n_580), .Y(n_1268) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_580), .A2(n_582), .B1(n_1311), .B2(n_1312), .Y(n_1310) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_581), .A2(n_620), .B(n_622), .Y(n_619) );
INVx2_ASAP7_75t_SL g800 ( .A(n_582), .Y(n_800) );
INVx2_ASAP7_75t_L g1213 ( .A(n_582), .Y(n_1213) );
OR2x2_ASAP7_75t_L g710 ( .A(n_586), .B(n_709), .Y(n_710) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx4f_ASAP7_75t_L g904 ( .A(n_587), .Y(n_904) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g1194 ( .A1(n_591), .A2(n_1186), .B1(n_1195), .B2(n_1196), .C(n_1200), .Y(n_1194) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_591), .A2(n_1256), .B1(n_1257), .B2(n_1258), .C(n_1259), .Y(n_1255) );
INVx1_ASAP7_75t_L g1308 ( .A(n_591), .Y(n_1308) );
INVx1_ASAP7_75t_L g1766 ( .A(n_591), .Y(n_1766) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_592), .Y(n_1103) );
BUFx3_ASAP7_75t_L g601 ( .A(n_595), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g1765 ( .A1(n_596), .A2(n_915), .B1(n_1751), .B2(n_1753), .Y(n_1765) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g977 ( .A(n_598), .Y(n_977) );
INVxp67_ASAP7_75t_L g1199 ( .A(n_598), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B1(n_603), .B2(n_605), .C(n_606), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_610), .Y(n_641) );
INVx2_ASAP7_75t_L g894 ( .A(n_610), .Y(n_894) );
INVx2_ASAP7_75t_L g1095 ( .A(n_610), .Y(n_1095) );
INVx1_ASAP7_75t_L g1776 ( .A(n_610), .Y(n_1776) );
INVx1_ASAP7_75t_L g763 ( .A(n_611), .Y(n_763) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI31xp33_ASAP7_75t_L g1371 ( .A1(n_613), .A2(n_1372), .A3(n_1383), .B(n_1392), .Y(n_1371) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI21x1_ASAP7_75t_L g661 ( .A1(n_614), .A2(n_662), .B(n_685), .Y(n_661) );
OAI31xp33_ASAP7_75t_L g1762 ( .A1(n_614), .A2(n_1763), .A3(n_1767), .B(n_1779), .Y(n_1762) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_620), .A2(n_622), .B1(n_720), .B2(n_721), .C(n_724), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_620), .A2(n_622), .B1(n_721), .B2(n_1311), .C(n_1312), .Y(n_1335) );
INVx1_ASAP7_75t_L g1351 ( .A(n_620), .Y(n_1351) );
AOI221xp5_ASAP7_75t_L g1783 ( .A1(n_620), .A2(n_622), .B1(n_721), .B2(n_1784), .C(n_1785), .Y(n_1783) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_621), .B(n_888), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1347 ( .A1(n_622), .A2(n_1348), .B1(n_1349), .B2(n_1350), .C(n_1352), .Y(n_1347) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_623), .Y(n_744) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR4xp75_ASAP7_75t_L g626 ( .A(n_627), .B(n_661), .C(n_706), .D(n_711), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_646), .Y(n_627) );
AOI33xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_633), .A3(n_637), .B1(n_639), .B2(n_642), .B3(n_645), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_SL g1131 ( .A1(n_630), .A2(n_1001), .B1(n_1132), .B2(n_1136), .Y(n_1131) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x4_ASAP7_75t_L g735 ( .A(n_631), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g789 ( .A(n_631), .Y(n_789) );
BUFx2_ASAP7_75t_L g882 ( .A(n_631), .Y(n_882) );
OR2x6_ASAP7_75t_L g898 ( .A(n_631), .B(n_774), .Y(n_898) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_631), .B(n_696), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1323 ( .A(n_631), .B(n_736), .Y(n_1323) );
OR2x2_ASAP7_75t_L g1694 ( .A(n_631), .B(n_774), .Y(n_1694) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_635), .A2(n_874), .B1(n_876), .B2(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g915 ( .A(n_635), .Y(n_915) );
INVx1_ASAP7_75t_L g1192 ( .A(n_635), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g1764 ( .A1(n_636), .A2(n_894), .B1(n_1750), .B2(n_1755), .Y(n_1764) );
INVx1_ASAP7_75t_L g901 ( .A(n_638), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_638), .B(n_660), .Y(n_912) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx4_ASAP7_75t_L g979 ( .A(n_641), .Y(n_979) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g712 ( .A(n_644), .B(n_709), .Y(n_712) );
OR2x6_ASAP7_75t_L g1042 ( .A(n_644), .B(n_709), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_652), .B1(n_653), .B2(n_656), .C(n_657), .Y(n_646) );
INVx2_ASAP7_75t_L g1009 ( .A(n_647), .Y(n_1009) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g910 ( .A(n_648), .Y(n_910) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OR2x6_ASAP7_75t_L g654 ( .A(n_651), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g660 ( .A(n_651), .Y(n_660) );
OR2x2_ASAP7_75t_L g911 ( .A(n_651), .B(n_655), .Y(n_911) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g989 ( .A(n_657), .Y(n_989) );
NOR3xp33_ASAP7_75t_L g1129 ( .A(n_657), .B(n_1130), .C(n_1131), .Y(n_1129) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI221x1_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_668), .B1(n_669), .B2(n_670), .C(n_671), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_663), .A2(n_669), .B1(n_866), .B2(n_867), .Y(n_865) );
INVx3_ASAP7_75t_L g1038 ( .A(n_663), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_663), .A2(n_669), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
AND2x4_ASAP7_75t_L g697 ( .A(n_664), .B(n_694), .Y(n_697) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g680 ( .A(n_666), .Y(n_680) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g1065 ( .A(n_667), .Y(n_1065) );
INVx3_ASAP7_75t_L g1037 ( .A(n_669), .Y(n_1037) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_677), .B(n_682), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_674), .B(n_675), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g1680 ( .A1(n_673), .A2(n_1681), .B1(n_1682), .B2(n_1683), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_676), .B(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
INVx2_ASAP7_75t_L g945 ( .A(n_678), .Y(n_945) );
INVx1_ASAP7_75t_L g1331 ( .A(n_680), .Y(n_1331) );
INVx1_ASAP7_75t_L g701 ( .A(n_683), .Y(n_701) );
INVx1_ASAP7_75t_L g888 ( .A(n_683), .Y(n_888) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI221xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_690), .B1(n_697), .B2(n_698), .C(n_699), .Y(n_685) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx3_ASAP7_75t_L g948 ( .A(n_689), .Y(n_948) );
INVx2_ASAP7_75t_L g1177 ( .A(n_689), .Y(n_1177) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx6f_ASAP7_75t_L g1018 ( .A(n_692), .Y(n_1018) );
INVx3_ASAP7_75t_L g1334 ( .A(n_692), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g1019 ( .A(n_696), .Y(n_1019) );
INVx8_ASAP7_75t_L g851 ( .A(n_697), .Y(n_851) );
CKINVDCx11_ASAP7_75t_R g1025 ( .A(n_702), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
BUFx3_ASAP7_75t_L g738 ( .A(n_705), .Y(n_738) );
OR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OR2x6_ASAP7_75t_L g713 ( .A(n_709), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g916 ( .A(n_709), .Y(n_916) );
INVx1_ASAP7_75t_L g1005 ( .A(n_714), .Y(n_1005) );
OAI21xp33_ASAP7_75t_L g1082 ( .A1(n_714), .A2(n_1083), .B(n_1084), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1381 ( .A1(n_714), .A2(n_970), .B1(n_1355), .B2(n_1357), .C(n_1382), .Y(n_1381) );
BUFx3_ASAP7_75t_L g1696 ( .A(n_714), .Y(n_1696) );
INVx2_ASAP7_75t_L g783 ( .A(n_716), .Y(n_783) );
XOR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_782), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_748), .Y(n_717) );
AND4x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_725), .C(n_728), .D(n_732), .Y(n_718) );
HB1xp67_ASAP7_75t_L g1348 ( .A(n_721), .Y(n_1348) );
AND2x4_ASAP7_75t_L g1706 ( .A(n_722), .B(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI221xp5_ASAP7_75t_L g758 ( .A1(n_727), .A2(n_729), .B1(n_759), .B2(n_762), .C(n_763), .Y(n_758) );
AOI33xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_737), .A3(n_741), .B1(n_745), .B2(n_746), .B3(n_747), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx3_ASAP7_75t_L g1684 ( .A(n_735), .Y(n_1684) );
INVx1_ASAP7_75t_L g1030 ( .A(n_736), .Y(n_1030) );
BUFx2_ASAP7_75t_SL g1126 ( .A(n_736), .Y(n_1126) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
BUFx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_751), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_749), .A2(n_1104), .B1(n_1188), .B2(n_1204), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g1208 ( .A1(n_749), .A2(n_789), .B1(n_1209), .B2(n_1227), .Y(n_1208) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g778 ( .A(n_757), .Y(n_778) );
INVx1_ASAP7_75t_L g967 ( .A(n_757), .Y(n_967) );
OAI211xp5_ASAP7_75t_L g1768 ( .A1(n_759), .A2(n_1769), .B(n_1770), .C(n_1771), .Y(n_1768) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp33_ASAP7_75t_L g1099 ( .A(n_761), .B(n_1100), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1002 ( .A1(n_762), .A2(n_1003), .B1(n_1004), .B2(n_1006), .C(n_1007), .Y(n_1002) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_782), .A2(n_1451), .B1(n_1452), .B2(n_1454), .Y(n_1450) );
INVx1_ASAP7_75t_L g1045 ( .A(n_784), .Y(n_1045) );
XNOR2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_845), .Y(n_784) );
INVx3_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g843 ( .A(n_787), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_810), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B1(n_808), .B2(n_809), .Y(n_788) );
NOR2xp67_ASAP7_75t_L g886 ( .A(n_789), .B(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g1320 ( .A(n_789), .Y(n_1320) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_801), .C(n_805), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_796), .B2(n_797), .C(n_798), .Y(n_791) );
BUFx6f_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g1303 ( .A(n_795), .Y(n_1303) );
BUFx3_ASAP7_75t_L g1380 ( .A(n_795), .Y(n_1380) );
INVx1_ASAP7_75t_L g1078 ( .A(n_796), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g1261 ( .A1(n_796), .A2(n_1262), .B1(n_1263), .B2(n_1264), .C(n_1267), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_797), .A2(n_807), .B1(n_830), .B2(n_837), .Y(n_836) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_804), .A2(n_806), .B1(n_824), .B2(n_841), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g1250 ( .A1(n_809), .A2(n_1251), .B1(n_1269), .B2(n_1270), .Y(n_1250) );
NOR3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_819), .C(n_822), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_815), .Y(n_811) );
INVx2_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g1169 ( .A(n_825), .Y(n_1169) );
INVx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_830), .A2(n_1174), .B1(n_1175), .B2(n_1176), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1240 ( .A1(n_830), .A2(n_1176), .B1(n_1241), .B2(n_1242), .Y(n_1240) );
BUFx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx2_ASAP7_75t_L g1754 ( .A(n_831), .Y(n_1754) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_832), .Y(n_873) );
INVx1_ASAP7_75t_L g953 ( .A(n_832), .Y(n_953) );
INVx2_ASAP7_75t_L g1013 ( .A(n_832), .Y(n_1013) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g1182 ( .A(n_839), .Y(n_1182) );
INVx1_ASAP7_75t_L g1329 ( .A(n_839), .Y(n_1329) );
OAI22xp33_ASAP7_75t_L g1281 ( .A1(n_841), .A2(n_1282), .B1(n_1284), .B2(n_1285), .Y(n_1281) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
XOR2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_982), .Y(n_845) );
XNOR2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_921), .Y(n_846) );
NAND4xp25_ASAP7_75t_L g848 ( .A(n_849), .B(n_883), .C(n_889), .D(n_913), .Y(n_848) );
OAI21xp5_ASAP7_75t_SL g849 ( .A1(n_850), .A2(n_868), .B(n_882), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_858), .B(n_864), .Y(n_852) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_SL g862 ( .A(n_863), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_866), .A2(n_867), .B1(n_903), .B2(n_905), .Y(n_902) );
CKINVDCx6p67_ASAP7_75t_R g869 ( .A(n_870), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_872), .A2(n_1254), .B1(n_1262), .B2(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_875), .A2(n_1287), .B1(n_1288), .B2(n_1289), .Y(n_1286) );
OAI21xp5_ASAP7_75t_SL g877 ( .A1(n_878), .A2(n_879), .B(n_880), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g1245 ( .A1(n_878), .A2(n_1220), .B1(n_1225), .B2(n_1246), .Y(n_1245) );
CKINVDCx8_ASAP7_75t_R g1269 ( .A(n_882), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_885), .B(n_987), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_885), .B(n_1128), .Y(n_1127) );
AOI221xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_897), .B1(n_899), .B2(n_907), .C(n_908), .Y(n_889) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1202 ( .A(n_896), .Y(n_1202) );
INVx1_ASAP7_75t_L g1266 ( .A(n_896), .Y(n_1266) );
INVx1_ASAP7_75t_L g991 ( .A(n_897), .Y(n_991) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx4_ASAP7_75t_L g1001 ( .A(n_907), .Y(n_1001) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_917), .B1(n_918), .B2(n_919), .C(n_920), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_914), .A2(n_918), .B1(n_1141), .B2(n_1142), .C(n_1143), .Y(n_1140) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
XNOR2x1_ASAP7_75t_SL g921 ( .A(n_922), .B(n_923), .Y(n_921) );
AND2x2_ASAP7_75t_L g923 ( .A(n_924), .B(n_958), .Y(n_923) );
NOR3xp33_ASAP7_75t_SL g924 ( .A(n_925), .B(n_933), .C(n_935), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_929), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_928), .A2(n_930), .B1(n_969), .B2(n_970), .C(n_971), .Y(n_968) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_941), .A2(n_1246), .B1(n_1253), .B2(n_1257), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .B1(n_946), .B2(n_947), .Y(n_942) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g1179 ( .A(n_945), .Y(n_1179) );
INVx2_ASAP7_75t_L g1244 ( .A(n_945), .Y(n_1244) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g1058 ( .A1(n_953), .A2(n_1059), .B1(n_1060), .B2(n_1061), .C(n_1062), .Y(n_1058) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_973), .C(n_980), .Y(n_959) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g1379 ( .A(n_966), .Y(n_1379) );
BUFx3_ASAP7_75t_L g1386 ( .A(n_966), .Y(n_1386) );
OAI211xp5_ASAP7_75t_L g1091 ( .A1(n_969), .A2(n_1092), .B(n_1093), .C(n_1094), .Y(n_1091) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_970), .A2(n_1124), .B1(n_1125), .B2(n_1133), .C(n_1135), .Y(n_1132) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
XNOR2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_985), .Y(n_983) );
AND4x1_ASAP7_75t_L g985 ( .A(n_986), .B(n_988), .C(n_1010), .D(n_1040), .Y(n_985) );
NOR3xp33_ASAP7_75t_SL g988 ( .A(n_989), .B(n_990), .C(n_1008), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B1(n_1001), .B2(n_1002), .Y(n_990) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
OAI22xp5_ASAP7_75t_SL g1693 ( .A1(n_1001), .A2(n_1694), .B1(n_1695), .B2(n_1698), .Y(n_1693) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI31xp33_ASAP7_75t_L g1010 ( .A1(n_1011), .A2(n_1026), .A3(n_1036), .B(n_1039), .Y(n_1010) );
AOI222xp33_ASAP7_75t_L g1704 ( .A1(n_1017), .A2(n_1664), .B1(n_1666), .B2(n_1700), .C1(n_1705), .C2(n_1706), .Y(n_1704) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1022), .B1(n_1024), .B2(n_1025), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1033 ( .A(n_1034), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1043), .Y(n_1040) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
XNOR2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1147), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1050), .B1(n_1105), .B2(n_1146), .Y(n_1048) );
INVxp67_ASAP7_75t_SL g1049 ( .A(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
NAND3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1069), .C(n_1076), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1068), .Y(n_1054) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_1061), .A2(n_1086), .B1(n_1087), .B2(n_1089), .Y(n_1085) );
NAND3xp33_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .C(n_1067), .Y(n_1063) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1065), .Y(n_1291) );
AOI33xp33_ASAP7_75t_L g1322 ( .A1(n_1067), .A2(n_1323), .A3(n_1324), .B1(n_1326), .B2(n_1330), .B3(n_1332), .Y(n_1322) );
NOR2xp33_ASAP7_75t_SL g1069 ( .A(n_1070), .B(n_1073), .Y(n_1069) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
OAI31xp33_ASAP7_75t_SL g1076 ( .A1(n_1077), .A2(n_1079), .A3(n_1081), .B(n_1104), .Y(n_1076) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1080), .Y(n_1256) );
OAI211xp5_ASAP7_75t_SL g1081 ( .A1(n_1082), .A2(n_1085), .B(n_1091), .C(n_1097), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_1087), .A2(n_1133), .B1(n_1137), .B2(n_1138), .C(n_1139), .Y(n_1136) );
INVx2_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
BUFx6f_ASAP7_75t_L g1201 ( .A(n_1095), .Y(n_1201) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1105), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1107), .Y(n_1144) );
NAND4xp25_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1127), .C(n_1129), .D(n_1140), .Y(n_1107) );
AOI21xp5_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1115), .B(n_1116), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1120), .B1(n_1121), .B2(n_1122), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g1741 ( .A1(n_1119), .A2(n_1742), .B1(n_1743), .B2(n_1744), .Y(n_1741) );
OAI21xp33_ASAP7_75t_L g1305 ( .A1(n_1133), .A2(n_1306), .B(n_1307), .Y(n_1305) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1134), .Y(n_1315) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1134), .Y(n_1774) );
AOI22xp5_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1149), .B1(n_1343), .B2(n_1344), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
AO22x1_ASAP7_75t_L g1149 ( .A1(n_1150), .A2(n_1151), .B1(n_1247), .B2(n_1342), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
AO22x2_ASAP7_75t_L g1151 ( .A1(n_1152), .A2(n_1153), .B1(n_1205), .B2(n_1206), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
XNOR2xp5_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1155), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1187), .Y(n_1155) );
NOR3xp33_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1164), .C(n_1166), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1161), .Y(n_1157) );
OAI22xp33_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1169), .B1(n_1170), .B2(n_1171), .Y(n_1167) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1180), .B1(n_1181), .B2(n_1183), .Y(n_1178) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1194), .C(n_1203), .Y(n_1188) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1198), .Y(n_1222) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1228), .Y(n_1207) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1219), .C(n_1224), .Y(n_1209) );
NOR3xp33_ASAP7_75t_SL g1228 ( .A(n_1229), .B(n_1235), .C(n_1236), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1233), .Y(n_1229) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1247), .Y(n_1342) );
XOR2x2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1295), .Y(n_1247) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1249), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1271), .Y(n_1249) );
NAND3xp33_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1255), .C(n_1261), .Y(n_1251) );
NOR3xp33_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1279), .C(n_1280), .Y(n_1271) );
NAND2xp5_ASAP7_75t_SL g1272 ( .A(n_1273), .B(n_1276), .Y(n_1272) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1296), .Y(n_1341) );
NAND4xp75_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .C(n_1321), .D(n_1336), .Y(n_1296) );
OAI31xp33_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1309), .A3(n_1318), .B(n_1319), .Y(n_1298) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B1(n_1303), .B2(n_1304), .Y(n_1300) );
OAI211xp5_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1315), .B(n_1316), .C(n_1317), .Y(n_1313) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_SL g1321 ( .A(n_1322), .B(n_1335), .Y(n_1321) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1369), .Y(n_1345) );
AND4x1_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1353), .C(n_1356), .D(n_1359), .Y(n_1346) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
OAI221xp5_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1637), .B1(n_1639), .B2(n_1727), .C(n_1731), .Y(n_1396) );
AOI21xp5_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1542), .B(n_1586), .Y(n_1397) );
NAND5xp2_ASAP7_75t_SL g1398 ( .A(n_1399), .B(n_1481), .C(n_1510), .D(n_1533), .E(n_1537), .Y(n_1398) );
AOI21xp5_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1438), .B(n_1459), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1421), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1401), .B(n_1448), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_1401), .B(n_1536), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1401), .B(n_1470), .Y(n_1560) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1401), .B(n_1448), .Y(n_1571) );
INVx2_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1402), .B(n_1468), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1402), .B(n_1448), .Y(n_1480) );
BUFx2_ASAP7_75t_L g1487 ( .A(n_1402), .Y(n_1487) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1402), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1402), .B(n_1421), .Y(n_1545) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1402), .B(n_1478), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1402), .B(n_1470), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1415), .Y(n_1402) );
AND2x4_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1410), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1406), .B(n_1411), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1409), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1409), .Y(n_1418) );
AND2x4_ASAP7_75t_L g1412 ( .A(n_1410), .B(n_1413), .Y(n_1412) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1437 ( .A(n_1411), .B(n_1414), .Y(n_1437) );
BUFx2_ASAP7_75t_L g1443 ( .A(n_1412), .Y(n_1443) );
HB1xp67_ASAP7_75t_L g1788 ( .A(n_1413), .Y(n_1788) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1416), .Y(n_1456) );
BUFx3_ASAP7_75t_L g1502 ( .A(n_1416), .Y(n_1502) );
AND2x4_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1419), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1417), .B(n_1419), .Y(n_1426) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_1418), .B(n_1419), .Y(n_1420) );
INVx2_ASAP7_75t_L g1446 ( .A(n_1420), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1427), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1422), .B(n_1474), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1422), .B(n_1465), .Y(n_1530) );
A2O1A1Ixp33_ASAP7_75t_L g1603 ( .A1(n_1422), .A2(n_1604), .B(n_1607), .C(n_1608), .Y(n_1603) );
INVxp67_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
BUFx2_ASAP7_75t_L g1468 ( .A(n_1423), .Y(n_1468) );
BUFx3_ASAP7_75t_L g1478 ( .A(n_1423), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1423), .B(n_1465), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1425), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1427), .B(n_1468), .Y(n_1499) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1427), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1432), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1428), .B(n_1478), .Y(n_1483) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1428), .B(n_1468), .Y(n_1549) );
INVx2_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1429), .B(n_1432), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1429), .B(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1429), .B(n_1478), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1429), .B(n_1432), .Y(n_1514) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_1429), .B(n_1478), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1431), .Y(n_1429) );
INVx2_ASAP7_75t_SL g1475 ( .A(n_1432), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1432), .B(n_1478), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g1433 ( .A1(n_1434), .A2(n_1435), .B1(n_1436), .B2(n_1437), .Y(n_1433) );
BUFx6f_ASAP7_75t_L g1451 ( .A(n_1435), .Y(n_1451) );
XNOR2xp5_ASAP7_75t_L g1641 ( .A(n_1436), .B(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1437), .Y(n_1453) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1438), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1447), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1439), .B(n_1509), .Y(n_1508) );
INVx2_ASAP7_75t_L g1525 ( .A(n_1439), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1439), .B(n_1540), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1439), .B(n_1448), .Y(n_1575) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1440), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_1440), .B(n_1460), .Y(n_1623) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1516 ( .A(n_1441), .B(n_1460), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1441), .B(n_1471), .Y(n_1518) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1441), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1444), .Y(n_1441) );
INVx2_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
OAI22xp5_ASAP7_75t_L g1455 ( .A1(n_1446), .A2(n_1456), .B1(n_1457), .B2(n_1458), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1447), .B(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1447), .Y(n_1585) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1448), .B(n_1460), .Y(n_1488) );
INVx2_ASAP7_75t_SL g1524 ( .A(n_1448), .Y(n_1524) );
AND2x4_ASAP7_75t_L g1540 ( .A(n_1448), .B(n_1471), .Y(n_1540) );
HB1xp67_ASAP7_75t_L g1577 ( .A(n_1448), .Y(n_1577) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_1449), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1449), .B(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1449), .B(n_1460), .Y(n_1532) );
OR2x2_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1455), .Y(n_1449) );
BUFx3_ASAP7_75t_L g1505 ( .A(n_1451), .Y(n_1505) );
HB1xp67_ASAP7_75t_L g1507 ( .A(n_1452), .Y(n_1507) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OAI211xp5_ASAP7_75t_SL g1459 ( .A1(n_1460), .A2(n_1463), .B(n_1469), .C(n_1476), .Y(n_1459) );
INVx3_ASAP7_75t_L g1471 ( .A(n_1460), .Y(n_1471) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1460), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1461), .B(n_1462), .Y(n_1460) );
OAI321xp33_ASAP7_75t_L g1568 ( .A1(n_1463), .A2(n_1483), .A3(n_1514), .B1(n_1562), .B2(n_1569), .C(n_1570), .Y(n_1568) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1464), .B(n_1524), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1464), .B(n_1615), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1465), .B(n_1467), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1465), .B(n_1494), .Y(n_1579) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1592 ( .A(n_1466), .B(n_1569), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1467), .B(n_1514), .Y(n_1600) );
NOR2x1_ASAP7_75t_L g1567 ( .A(n_1468), .B(n_1475), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1468), .B(n_1514), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1472), .Y(n_1469) );
AOI221xp5_ASAP7_75t_L g1543 ( .A1(n_1470), .A2(n_1544), .B1(n_1546), .B2(n_1552), .C(n_1553), .Y(n_1543) );
NOR2xp33_ASAP7_75t_L g1479 ( .A(n_1471), .B(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1471), .Y(n_1491) );
OR2x2_ASAP7_75t_L g1597 ( .A(n_1471), .B(n_1598), .Y(n_1597) );
AOI221xp5_ASAP7_75t_L g1612 ( .A1(n_1471), .A2(n_1515), .B1(n_1613), .B2(n_1616), .C(n_1619), .Y(n_1612) );
O2A1O1Ixp33_ASAP7_75t_L g1556 ( .A1(n_1472), .A2(n_1539), .B(n_1557), .C(n_1559), .Y(n_1556) );
AOI222xp33_ASAP7_75t_L g1593 ( .A1(n_1472), .A2(n_1518), .B1(n_1594), .B2(n_1596), .C1(n_1599), .C2(n_1601), .Y(n_1593) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1595 ( .A(n_1473), .B(n_1486), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1474), .B(n_1478), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1554 ( .A(n_1474), .B(n_1487), .Y(n_1554) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1474), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1475), .B(n_1478), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1479), .Y(n_1476) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1477), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1477), .B(n_1494), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_1478), .B(n_1513), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1478), .B(n_1527), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1478), .B(n_1579), .Y(n_1607) );
O2A1O1Ixp33_ASAP7_75t_L g1619 ( .A1(n_1480), .A2(n_1620), .B(n_1621), .C(n_1622), .Y(n_1619) );
A2O1A1Ixp33_ASAP7_75t_L g1481 ( .A1(n_1482), .A2(n_1484), .B(n_1489), .C(n_1508), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1511 ( .A(n_1483), .B(n_1512), .Y(n_1511) );
O2A1O1Ixp33_ASAP7_75t_L g1553 ( .A1(n_1483), .A2(n_1487), .B(n_1554), .C(n_1555), .Y(n_1553) );
NOR2xp33_ASAP7_75t_L g1559 ( .A(n_1483), .B(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1488), .Y(n_1485) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1486), .B(n_1521), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1566 ( .A(n_1486), .B(n_1567), .Y(n_1566) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
AOI321xp33_ASAP7_75t_L g1510 ( .A1(n_1487), .A2(n_1511), .A3(n_1515), .B1(n_1517), .B2(n_1519), .C(n_1528), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_1487), .B(n_1532), .Y(n_1531) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1487), .B(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_SL g1583 ( .A(n_1487), .B(n_1521), .Y(n_1583) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1488), .Y(n_1551) );
OAI211xp5_ASAP7_75t_SL g1489 ( .A1(n_1490), .A2(n_1492), .B(n_1496), .C(n_1500), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1546 ( .A1(n_1490), .A2(n_1547), .B1(n_1550), .B2(n_1551), .Y(n_1546) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
A2O1A1Ixp33_ASAP7_75t_L g1581 ( .A1(n_1491), .A2(n_1582), .B(n_1584), .C(n_1585), .Y(n_1581) );
AOI31xp33_ASAP7_75t_L g1632 ( .A1(n_1492), .A2(n_1529), .A3(n_1633), .B(n_1635), .Y(n_1632) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1494), .B(n_1514), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1494), .B(n_1524), .Y(n_1629) );
INVxp67_ASAP7_75t_L g1550 ( .A(n_1495), .Y(n_1550) );
INVxp67_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1499), .Y(n_1497) );
INVx2_ASAP7_75t_L g1580 ( .A(n_1500), .Y(n_1580) );
INVx3_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx3_ASAP7_75t_L g1509 ( .A(n_1501), .Y(n_1509) );
OAI22xp33_ASAP7_75t_L g1503 ( .A1(n_1504), .A2(n_1505), .B1(n_1506), .B2(n_1507), .Y(n_1503) );
BUFx2_ASAP7_75t_SL g1638 ( .A(n_1507), .Y(n_1638) );
AOI21xp5_ASAP7_75t_L g1528 ( .A1(n_1513), .A2(n_1529), .B(n_1531), .Y(n_1528) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1515), .B(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
NOR2xp33_ASAP7_75t_L g1523 ( .A(n_1516), .B(n_1524), .Y(n_1523) );
OAI22xp33_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1522), .B1(n_1525), .B2(n_1526), .Y(n_1519) );
INVxp33_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1564 ( .A(n_1524), .B(n_1565), .Y(n_1564) );
NOR2xp33_ASAP7_75t_L g1591 ( .A(n_1524), .B(n_1592), .Y(n_1591) );
INVx2_ASAP7_75t_L g1615 ( .A(n_1524), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1524), .B(n_1618), .Y(n_1617) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_1524), .B(n_1597), .Y(n_1636) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1525), .Y(n_1552) );
A2O1A1Ixp33_ASAP7_75t_L g1561 ( .A1(n_1525), .A2(n_1562), .B(n_1563), .C(n_1568), .Y(n_1561) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
NOR2xp33_ASAP7_75t_L g1631 ( .A(n_1530), .B(n_1536), .Y(n_1631) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_1532), .A2(n_1541), .B1(n_1573), .B2(n_1574), .C(n_1576), .Y(n_1572) );
CKINVDCx5p33_ASAP7_75t_R g1611 ( .A(n_1532), .Y(n_1611) );
INVxp67_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVxp67_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1541), .Y(n_1538) );
NAND5xp2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1556), .C(n_1561), .D(n_1572), .E(n_1581), .Y(n_1542) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
AOI22xp5_ASAP7_75t_L g1587 ( .A1(n_1552), .A2(n_1588), .B1(n_1590), .B2(n_1591), .Y(n_1587) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1560), .Y(n_1625) );
INVxp67_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1573), .Y(n_1621) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
OAI21xp33_ASAP7_75t_L g1576 ( .A1(n_1577), .A2(n_1578), .B(n_1580), .Y(n_1576) );
NOR2xp33_ASAP7_75t_L g1599 ( .A(n_1577), .B(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
NAND5xp2_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1593), .C(n_1603), .D(n_1612), .E(n_1624), .Y(n_1586) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1589), .Y(n_1610) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1589), .Y(n_1628) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
OR2x2_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1611), .Y(n_1609) );
INVxp67_ASAP7_75t_SL g1613 ( .A(n_1614), .Y(n_1613) );
INVxp67_ASAP7_75t_SL g1616 ( .A(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
O2A1O1Ixp33_ASAP7_75t_L g1624 ( .A1(n_1625), .A2(n_1626), .B(n_1630), .C(n_1632), .Y(n_1624) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
INVxp67_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
HB1xp67_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
NAND3x1_ASAP7_75t_SL g1642 ( .A(n_1643), .B(n_1676), .C(n_1702), .Y(n_1642) );
OAI31xp33_ASAP7_75t_L g1643 ( .A1(n_1644), .A2(n_1653), .A3(n_1667), .B(n_1674), .Y(n_1643) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1647), .B(n_1656), .Y(n_1655) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1647), .Y(n_1659) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx4_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
AND2x4_ASAP7_75t_L g1661 ( .A(n_1651), .B(n_1662), .Y(n_1661) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
CKINVDCx8_ASAP7_75t_R g1657 ( .A(n_1658), .Y(n_1657) );
AOI22xp33_ASAP7_75t_L g1660 ( .A1(n_1661), .A2(n_1664), .B1(n_1665), .B2(n_1666), .Y(n_1660) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
CKINVDCx6p67_ASAP7_75t_R g1668 ( .A(n_1669), .Y(n_1668) );
INVx4_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_SL g1672 ( .A(n_1673), .Y(n_1672) );
INVxp67_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx3_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
AOI22xp33_ASAP7_75t_L g1709 ( .A1(n_1699), .A2(n_1710), .B1(n_1711), .B2(n_1712), .Y(n_1709) );
OAI21xp5_ASAP7_75t_L g1702 ( .A1(n_1703), .A2(n_1718), .B(n_1725), .Y(n_1702) );
NAND3xp33_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1709), .C(n_1715), .Y(n_1703) );
INVxp67_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1708), .Y(n_1717) );
INVx4_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1714), .Y(n_1720) );
AND2x4_ASAP7_75t_L g1722 ( .A(n_1714), .B(n_1723), .Y(n_1722) );
CKINVDCx11_ASAP7_75t_R g1715 ( .A(n_1716), .Y(n_1715) );
INVx5_ASAP7_75t_SL g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
CKINVDCx16_ASAP7_75t_R g1725 ( .A(n_1726), .Y(n_1725) );
INVx2_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
CKINVDCx5p33_ASAP7_75t_R g1733 ( .A(n_1734), .Y(n_1733) );
OAI21xp5_ASAP7_75t_L g1787 ( .A1(n_1735), .A2(n_1788), .B(n_1789), .Y(n_1787) );
INVxp33_ASAP7_75t_SL g1736 ( .A(n_1737), .Y(n_1736) );
INVx1_ASAP7_75t_L g1738 ( .A(n_1739), .Y(n_1738) );
NAND4xp75_ASAP7_75t_L g1739 ( .A(n_1740), .B(n_1758), .C(n_1762), .D(n_1783), .Y(n_1739) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
OAI211xp5_ASAP7_75t_L g1773 ( .A1(n_1748), .A2(n_1774), .B(n_1775), .C(n_1777), .Y(n_1773) );
OAI22xp5_ASAP7_75t_L g1752 ( .A1(n_1753), .A2(n_1754), .B1(n_1755), .B2(n_1756), .Y(n_1752) );
NOR2x1_ASAP7_75t_L g1758 ( .A(n_1759), .B(n_1761), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1768), .B(n_1773), .Y(n_1767) );
BUFx2_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
endmodule