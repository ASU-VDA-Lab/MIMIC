module real_aes_297_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_617;
wire n_552;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g521 ( .A(n_0), .B(n_132), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_1), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_2), .B(n_114), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_3), .B(n_130), .Y(n_149) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_5), .B(n_114), .Y(n_452) );
NAND2xp33_ASAP7_75t_SL g506 ( .A(n_6), .B(n_120), .Y(n_506) );
INVx1_ASAP7_75t_L g499 ( .A(n_7), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_8), .Y(n_747) );
AND2x2_ASAP7_75t_L g450 ( .A(n_9), .B(n_135), .Y(n_450) );
AND2x2_ASAP7_75t_L g151 ( .A(n_10), .B(n_139), .Y(n_151) );
AND2x2_ASAP7_75t_L g160 ( .A(n_11), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_13), .B(n_130), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_14), .Y(n_434) );
AOI221x1_ASAP7_75t_L g502 ( .A1(n_15), .A2(n_123), .B1(n_161), .B2(n_503), .C(n_505), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_16), .B(n_114), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_17), .B(n_114), .Y(n_194) );
INVx1_ASAP7_75t_L g438 ( .A(n_18), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_19), .A2(n_86), .B1(n_114), .B2(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_20), .A2(n_123), .B(n_454), .Y(n_453) );
AOI221xp5_ASAP7_75t_SL g511 ( .A1(n_21), .A2(n_34), .B1(n_114), .B2(n_123), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_22), .B(n_132), .Y(n_455) );
OR2x2_ASAP7_75t_L g137 ( .A(n_23), .B(n_85), .Y(n_137) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_23), .A2(n_85), .B(n_136), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_24), .B(n_130), .Y(n_493) );
INVxp67_ASAP7_75t_L g501 ( .A(n_25), .Y(n_501) );
AND2x2_ASAP7_75t_L g474 ( .A(n_26), .B(n_134), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_27), .A2(n_123), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_28), .A2(n_161), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_29), .B(n_130), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_30), .A2(n_123), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_31), .B(n_130), .Y(n_178) );
AND2x2_ASAP7_75t_L g120 ( .A(n_32), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g124 ( .A(n_32), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g232 ( .A(n_32), .Y(n_232) );
OR2x6_ASAP7_75t_L g436 ( .A(n_33), .B(n_437), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_33), .B(n_434), .C(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_35), .B(n_114), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_36), .A2(n_78), .B1(n_123), .B2(n_230), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_37), .B(n_130), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_38), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_39), .B(n_132), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_40), .A2(n_123), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_41), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g524 ( .A(n_42), .B(n_134), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_43), .B(n_134), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_44), .B(n_114), .Y(n_166) );
INVx1_ASAP7_75t_L g117 ( .A(n_45), .Y(n_117) );
INVx1_ASAP7_75t_L g127 ( .A(n_45), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_46), .B(n_130), .Y(n_158) );
AND2x2_ASAP7_75t_L g185 ( .A(n_47), .B(n_134), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_48), .B(n_114), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_49), .B(n_132), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_50), .B(n_132), .Y(n_177) );
AND2x2_ASAP7_75t_L g465 ( .A(n_51), .B(n_134), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_52), .B(n_114), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_53), .B(n_130), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_54), .B(n_114), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_55), .A2(n_123), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_56), .B(n_132), .Y(n_463) );
AND2x2_ASAP7_75t_SL g494 ( .A(n_57), .B(n_135), .Y(n_494) );
AND2x2_ASAP7_75t_L g200 ( .A(n_58), .B(n_135), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_59), .A2(n_123), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_60), .B(n_130), .Y(n_456) );
AND2x2_ASAP7_75t_SL g484 ( .A(n_61), .B(n_139), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_62), .B(n_132), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_63), .B(n_132), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_64), .A2(n_89), .B1(n_123), .B2(n_230), .Y(n_229) );
AOI221x1_ASAP7_75t_L g102 ( .A1(n_65), .A2(n_103), .B1(n_718), .B2(n_719), .C(n_721), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g718 ( .A(n_65), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_66), .B(n_130), .Y(n_197) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
INVx1_ASAP7_75t_L g125 ( .A(n_67), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_68), .A2(n_720), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_68), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_69), .B(n_132), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_70), .A2(n_123), .B(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_71), .A2(n_123), .B(n_128), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_72), .A2(n_123), .B(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g180 ( .A(n_73), .B(n_135), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_74), .B(n_134), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_75), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_76), .B(n_114), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_77), .A2(n_80), .B1(n_114), .B2(n_224), .Y(n_482) );
INVx1_ASAP7_75t_L g439 ( .A(n_79), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_79), .B(n_438), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_81), .B(n_132), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_82), .B(n_132), .Y(n_514) );
AND2x2_ASAP7_75t_L g138 ( .A(n_83), .B(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_84), .A2(n_123), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_87), .B(n_130), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_88), .A2(n_123), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_90), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_91), .Y(n_725) );
BUFx2_ASAP7_75t_L g199 ( .A(n_92), .Y(n_199) );
INVxp67_ASAP7_75t_L g504 ( .A(n_93), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_94), .B(n_130), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_95), .A2(n_123), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_96), .B(n_114), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_97), .Y(n_749) );
BUFx2_ASAP7_75t_L g729 ( .A(n_98), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_741), .B(n_748), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_730), .Y(n_100) );
AOI21xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_724), .B(n_728), .Y(n_101) );
OAI21x1_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_431), .B(n_440), .Y(n_103) );
AO22x2_ASAP7_75t_L g719 ( .A1(n_104), .A2(n_432), .B1(n_441), .B2(n_720), .Y(n_719) );
INVx4_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_339), .Y(n_105) );
NOR3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_262), .C(n_297), .Y(n_106) );
OAI211xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_162), .B(n_214), .C(n_252), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_141), .Y(n_109) );
AND2x2_ASAP7_75t_L g245 ( .A(n_110), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_110), .B(n_251), .Y(n_285) );
AND2x2_ASAP7_75t_L g310 ( .A(n_110), .B(n_265), .Y(n_310) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g217 ( .A(n_111), .Y(n_217) );
OR2x2_ASAP7_75t_L g248 ( .A(n_111), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g256 ( .A(n_111), .B(n_152), .Y(n_256) );
AND2x2_ASAP7_75t_L g264 ( .A(n_111), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g291 ( .A(n_111), .B(n_292), .Y(n_291) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_111), .B(n_294), .Y(n_302) );
AND2x4_ASAP7_75t_L g319 ( .A(n_111), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g357 ( .A(n_111), .Y(n_357) );
AND2x4_ASAP7_75t_SL g362 ( .A(n_111), .B(n_142), .Y(n_362) );
OR2x6_ASAP7_75t_L g111 ( .A(n_112), .B(n_138), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_122), .B(n_134), .Y(n_112) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_120), .Y(n_114) );
INVx1_ASAP7_75t_L g507 ( .A(n_115), .Y(n_507) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
AND2x6_ASAP7_75t_L g132 ( .A(n_116), .B(n_125), .Y(n_132) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g130 ( .A(n_118), .B(n_127), .Y(n_130) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx5_ASAP7_75t_L g133 ( .A(n_120), .Y(n_133) );
AND2x2_ASAP7_75t_L g126 ( .A(n_121), .B(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_121), .Y(n_227) );
AND2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
BUFx3_ASAP7_75t_L g228 ( .A(n_124), .Y(n_228) );
INVx2_ASAP7_75t_L g234 ( .A(n_125), .Y(n_234) );
AND2x4_ASAP7_75t_L g230 ( .A(n_126), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g226 ( .A(n_127), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_131), .B(n_133), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_132), .B(n_199), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_133), .A2(n_148), .B(n_149), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_133), .A2(n_157), .B(n_158), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_133), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_133), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_133), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_133), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_133), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_133), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_133), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_133), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_133), .A2(n_521), .B(n_522), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_134), .Y(n_144) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_134), .A2(n_223), .B(n_229), .Y(n_222) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_134), .A2(n_511), .B(n_515), .Y(n_510) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x4_ASAP7_75t_L g171 ( .A(n_136), .B(n_137), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_139), .A2(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_SL g480 ( .A(n_139), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_139), .A2(n_489), .B(n_490), .Y(n_488) );
BUFx4f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_141), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_141), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_152), .Y(n_141) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_142), .Y(n_257) );
INVx2_ASAP7_75t_L g293 ( .A(n_142), .Y(n_293) );
INVx1_ASAP7_75t_L g320 ( .A(n_142), .Y(n_320) );
AND2x2_ASAP7_75t_L g419 ( .A(n_142), .B(n_329), .Y(n_419) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_143), .Y(n_251) );
AND2x2_ASAP7_75t_L g265 ( .A(n_143), .B(n_152), .Y(n_265) );
AOI21x1_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_151), .Y(n_143) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_144), .A2(n_459), .B(n_465), .Y(n_458) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_144), .A2(n_468), .B(n_474), .Y(n_467) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_144), .A2(n_468), .B(n_474), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
INVx2_ASAP7_75t_L g294 ( .A(n_152), .Y(n_294) );
INVx2_ASAP7_75t_L g329 ( .A(n_152), .Y(n_329) );
OR2x2_ASAP7_75t_L g414 ( .A(n_152), .B(n_246), .Y(n_414) );
AO21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_160), .Y(n_152) );
INVx4_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
AOI21x1_ASAP7_75t_L g517 ( .A1(n_153), .A2(n_518), .B(n_524), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
INVx3_ASAP7_75t_L g173 ( .A(n_161), .Y(n_173) );
AOI211xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_181), .B(n_201), .C(n_208), .Y(n_162) );
INVx2_ASAP7_75t_SL g303 ( .A(n_163), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_163), .B(n_182), .Y(n_309) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_172), .Y(n_163) );
INVx1_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx1_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx2_ASAP7_75t_L g236 ( .A(n_164), .Y(n_236) );
AND2x2_ASAP7_75t_L g260 ( .A(n_164), .B(n_184), .Y(n_260) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_164), .Y(n_289) );
OR2x2_ASAP7_75t_L g369 ( .A(n_164), .B(n_192), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_171), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_171), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_171), .A2(n_452), .B(n_453), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_171), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_171), .B(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_171), .B(n_504), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_171), .B(n_506), .C(n_507), .Y(n_505) );
AND2x2_ASAP7_75t_L g235 ( .A(n_172), .B(n_236), .Y(n_235) );
NOR2x1_ASAP7_75t_SL g267 ( .A(n_172), .B(n_192), .Y(n_267) );
AO21x1_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_172) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_173), .A2(n_174), .B(n_180), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g281 ( .A(n_182), .B(n_204), .Y(n_281) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_192), .Y(n_182) );
OR2x2_ASAP7_75t_L g213 ( .A(n_183), .B(n_192), .Y(n_213) );
BUFx2_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g288 ( .A(n_183), .B(n_289), .Y(n_288) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_184), .Y(n_240) );
AND2x2_ASAP7_75t_L g266 ( .A(n_184), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g276 ( .A(n_184), .Y(n_276) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_184), .B(n_192), .Y(n_314) );
OR2x2_ASAP7_75t_L g389 ( .A(n_184), .B(n_206), .Y(n_389) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx2_ASAP7_75t_SL g202 ( .A(n_192), .Y(n_202) );
AND2x2_ASAP7_75t_L g261 ( .A(n_192), .B(n_206), .Y(n_261) );
AND2x2_ASAP7_75t_L g332 ( .A(n_192), .B(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g353 ( .A(n_192), .Y(n_353) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_200), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g275 ( .A(n_204), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
BUFx2_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
AND2x2_ASAP7_75t_L g242 ( .A(n_206), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g333 ( .A(n_206), .Y(n_333) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
OR2x2_ASAP7_75t_L g279 ( .A(n_210), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_SL g321 ( .A(n_210), .B(n_322), .Y(n_321) );
AOI322xp5_ASAP7_75t_L g358 ( .A1(n_210), .A2(n_237), .A3(n_359), .B1(n_361), .B2(n_364), .C1(n_366), .C2(n_368), .Y(n_358) );
AND2x2_ASAP7_75t_L g423 ( .A(n_210), .B(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_211), .B(n_237), .Y(n_247) );
AOI322xp5_ASAP7_75t_L g298 ( .A1(n_212), .A2(n_299), .A3(n_303), .B1(n_304), .B2(n_307), .C1(n_309), .C2(n_310), .Y(n_298) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_L g350 ( .A(n_213), .B(n_303), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_213), .A2(n_410), .B1(n_412), .B2(n_415), .Y(n_409) );
OR2x2_ASAP7_75t_L g427 ( .A(n_213), .B(n_376), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_237), .B(n_238), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
AOI221xp5_ASAP7_75t_SL g277 ( .A1(n_216), .A2(n_253), .B1(n_278), .B2(n_281), .C(n_282), .Y(n_277) );
AND2x2_ASAP7_75t_L g304 ( .A(n_216), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_217), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g346 ( .A(n_217), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g375 ( .A(n_218), .Y(n_375) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_235), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_219), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g317 ( .A(n_219), .Y(n_317) );
OR2x2_ASAP7_75t_L g324 ( .A(n_219), .B(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g367 ( .A(n_220), .B(n_329), .Y(n_367) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AND2x4_ASAP7_75t_L g246 ( .A(n_221), .B(n_222), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_224), .A2(n_230), .B1(n_498), .B2(n_500), .Y(n_497) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_228), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NOR2x1p5_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_235), .B(n_296), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_235), .B(n_276), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_235), .Y(n_376) );
INVx1_ASAP7_75t_L g243 ( .A(n_236), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_244), .B1(n_247), .B2(n_248), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_SL g354 ( .A(n_242), .Y(n_354) );
AND2x2_ASAP7_75t_L g411 ( .A(n_243), .B(n_267), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_245), .B(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_SL g283 ( .A(n_245), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_245), .B(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
INVx2_ASAP7_75t_L g301 ( .A(n_246), .Y(n_301) );
AND2x2_ASAP7_75t_L g344 ( .A(n_246), .B(n_328), .Y(n_344) );
INVx1_ASAP7_75t_L g258 ( .A(n_248), .Y(n_258) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI21xp5_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_258), .B(n_259), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g337 ( .A(n_256), .Y(n_337) );
INVx2_ASAP7_75t_L g325 ( .A(n_257), .Y(n_325) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g322 ( .A(n_261), .B(n_276), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_261), .A2(n_359), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_263), .B(n_277), .Y(n_262) );
AOI32xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .A3(n_268), .B1(n_272), .B2(n_275), .Y(n_263) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_264), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_264), .A2(n_353), .B1(n_371), .B2(n_373), .C(n_379), .Y(n_370) );
AND2x2_ASAP7_75t_L g390 ( .A(n_264), .B(n_271), .Y(n_390) );
BUFx2_ASAP7_75t_L g274 ( .A(n_265), .Y(n_274) );
INVx1_ASAP7_75t_L g399 ( .A(n_265), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_265), .Y(n_404) );
INVx1_ASAP7_75t_SL g397 ( .A(n_266), .Y(n_397) );
INVx2_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
AND2x2_ASAP7_75t_L g392 ( .A(n_268), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x2_ASAP7_75t_L g364 ( .A(n_270), .B(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g336 ( .A(n_271), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_271), .B(n_362), .Y(n_384) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g296 ( .A(n_276), .Y(n_296) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g286 ( .A(n_280), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g295 ( .A(n_280), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g400 ( .A(n_281), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_286), .B1(n_290), .B2(n_295), .Y(n_282) );
INVx2_ASAP7_75t_SL g374 ( .A(n_284), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_284), .B(n_413), .Y(n_415) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_286), .A2(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g331 ( .A(n_288), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g359 ( .A(n_291), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g306 ( .A(n_292), .Y(n_306) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g348 ( .A(n_294), .Y(n_348) );
INVx1_ASAP7_75t_L g393 ( .A(n_295), .Y(n_393) );
NAND3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_311), .C(n_334), .Y(n_297) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_L g360 ( .A(n_300), .Y(n_360) );
AND2x2_ASAP7_75t_L g378 ( .A(n_300), .B(n_319), .Y(n_378) );
OR2x2_ASAP7_75t_L g417 ( .A(n_300), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_301), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g313 ( .A(n_303), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g380 ( .A(n_306), .B(n_317), .Y(n_380) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_309), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g421 ( .A(n_309), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B1(n_319), .B2(n_321), .C(n_323), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_312), .A2(n_335), .B(n_338), .Y(n_334) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx3_ASAP7_75t_L g365 ( .A(n_314), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_314), .B(n_408), .Y(n_407) );
INVxp33_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g326 ( .A(n_322), .Y(n_326) );
OAI22xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B1(n_327), .B2(n_330), .Y(n_323) );
INVx2_ASAP7_75t_L g429 ( .A(n_325), .Y(n_429) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g408 ( .A(n_333), .Y(n_408) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_385), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g340 ( .A(n_341), .B(n_358), .C(n_370), .D(n_382), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B(n_349), .C(n_351), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_346), .A2(n_352), .B(n_355), .Y(n_351) );
INVx2_ASAP7_75t_L g430 ( .A(n_347), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_348), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g363 ( .A(n_348), .Y(n_363) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
OR2x2_ASAP7_75t_L g425 ( .A(n_353), .B(n_389), .Y(n_425) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_360), .Y(n_396) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g366 ( .A(n_362), .B(n_367), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_362), .A2(n_392), .B(n_394), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_362), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g420 ( .A(n_362), .Y(n_420) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp33_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND4xp25_ASAP7_75t_L g385 ( .A(n_386), .B(n_391), .C(n_401), .D(n_422), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B1(n_398), .B2(n_400), .Y(n_394) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI211xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_405), .B(n_409), .C(n_416), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_421), .Y(n_416) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_426), .B(n_428), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_SL g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x6_ASAP7_75t_SL g441 ( .A(n_434), .B(n_436), .Y(n_441) );
OR2x2_ASAP7_75t_L g723 ( .A(n_434), .B(n_436), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_434), .B(n_435), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx2_ASAP7_75t_L g720 ( .A(n_442), .Y(n_720) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_640), .Y(n_442) );
NOR3xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_564), .C(n_614), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_544), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_485), .B(n_525), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_475), .Y(n_447) );
INVx1_ASAP7_75t_SL g650 ( .A(n_448), .Y(n_650) );
AOI32xp33_ASAP7_75t_L g681 ( .A1(n_448), .A2(n_663), .A3(n_682), .B1(n_683), .B2(n_684), .Y(n_681) );
AND2x2_ASAP7_75t_L g683 ( .A(n_448), .B(n_540), .Y(n_683) );
AND2x4_ASAP7_75t_SL g448 ( .A(n_449), .B(n_457), .Y(n_448) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_449), .Y(n_476) );
INVx5_ASAP7_75t_L g543 ( .A(n_449), .Y(n_543) );
OR2x2_ASAP7_75t_L g550 ( .A(n_449), .B(n_542), .Y(n_550) );
INVx2_ASAP7_75t_L g555 ( .A(n_449), .Y(n_555) );
AND2x2_ASAP7_75t_L g567 ( .A(n_449), .B(n_458), .Y(n_567) );
AND2x2_ASAP7_75t_L g572 ( .A(n_449), .B(n_466), .Y(n_572) );
OR2x2_ASAP7_75t_L g579 ( .A(n_449), .B(n_478), .Y(n_579) );
AND2x4_ASAP7_75t_L g588 ( .A(n_449), .B(n_467), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_SL g630 ( .A1(n_449), .A2(n_546), .B(n_581), .C(n_619), .Y(n_630) );
OR2x6_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx3_ASAP7_75t_SL g580 ( .A(n_457), .Y(n_580) );
AND2x2_ASAP7_75t_L g626 ( .A(n_457), .B(n_543), .Y(n_626) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_466), .Y(n_457) );
AND2x2_ASAP7_75t_L g477 ( .A(n_458), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g557 ( .A(n_458), .B(n_467), .Y(n_557) );
AND2x2_ASAP7_75t_L g561 ( .A(n_458), .B(n_540), .Y(n_561) );
INVx1_ASAP7_75t_L g587 ( .A(n_458), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_458), .B(n_467), .Y(n_609) );
INVx2_ASAP7_75t_L g613 ( .A(n_458), .Y(n_613) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_458), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_458), .B(n_543), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g624 ( .A(n_467), .B(n_478), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g634 ( .A(n_476), .Y(n_634) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_476), .B(n_551), .Y(n_659) );
AND2x2_ASAP7_75t_L g701 ( .A(n_477), .B(n_543), .Y(n_701) );
AND2x2_ASAP7_75t_L g612 ( .A(n_478), .B(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g675 ( .A(n_478), .Y(n_675) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_479), .Y(n_540) );
AOI21x1_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_484), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_485), .A2(n_566), .B1(n_668), .B2(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_508), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_486), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_486), .B(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .Y(n_486) );
INVx2_ASAP7_75t_L g531 ( .A(n_487), .Y(n_531) );
OR2x2_ASAP7_75t_L g535 ( .A(n_487), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_487), .B(n_548), .Y(n_553) );
AND2x4_ASAP7_75t_SL g563 ( .A(n_487), .B(n_496), .Y(n_563) );
OR2x2_ASAP7_75t_L g570 ( .A(n_487), .B(n_510), .Y(n_570) );
OR2x2_ASAP7_75t_L g582 ( .A(n_487), .B(n_496), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_487), .B(n_510), .Y(n_596) );
INVx1_ASAP7_75t_L g601 ( .A(n_487), .Y(n_601) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_487), .Y(n_619) );
AND2x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_602), .Y(n_682) );
INVx2_ASAP7_75t_L g686 ( .A(n_487), .Y(n_686) );
OR2x2_ASAP7_75t_L g693 ( .A(n_487), .B(n_583), .Y(n_693) );
OR2x2_ASAP7_75t_L g715 ( .A(n_487), .B(n_716), .Y(n_715) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
AND2x2_ASAP7_75t_L g532 ( .A(n_495), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_495), .B(n_516), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_495), .B(n_592), .Y(n_654) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
AND2x4_ASAP7_75t_L g602 ( .A(n_496), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_496), .B(n_547), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_496), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_496), .B(n_536), .Y(n_695) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_502), .Y(n_496) );
AND2x2_ASAP7_75t_L g562 ( .A(n_508), .B(n_563), .Y(n_562) );
AO221x1_ASAP7_75t_L g636 ( .A1(n_508), .A2(n_551), .B1(n_582), .B2(n_637), .C(n_638), .Y(n_636) );
OAI322xp33_ASAP7_75t_L g688 ( .A1(n_508), .A2(n_608), .A3(n_689), .B1(n_691), .B2(n_692), .C1(n_693), .C2(n_694), .Y(n_688) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_516), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx3_ASAP7_75t_L g530 ( .A(n_510), .Y(n_530) );
INVx2_ASAP7_75t_L g536 ( .A(n_510), .Y(n_536) );
AND2x2_ASAP7_75t_L g548 ( .A(n_510), .B(n_516), .Y(n_548) );
INVx1_ASAP7_75t_L g593 ( .A(n_510), .Y(n_593) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_510), .Y(n_649) );
INVx1_ASAP7_75t_L g533 ( .A(n_516), .Y(n_533) );
OR2x2_ASAP7_75t_L g583 ( .A(n_516), .B(n_536), .Y(n_583) );
INVx2_ASAP7_75t_L g603 ( .A(n_516), .Y(n_603) );
INVx1_ASAP7_75t_L g656 ( .A(n_516), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_516), .B(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI21xp33_ASAP7_75t_SL g526 ( .A1(n_527), .A2(n_534), .B(n_537), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_527), .A2(n_566), .B1(n_568), .B2(n_572), .C(n_573), .Y(n_565) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
NOR2x1p5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g652 ( .A(n_531), .Y(n_652) );
INVx1_ASAP7_75t_SL g571 ( .A(n_532), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_532), .A2(n_677), .B(n_679), .Y(n_676) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_533), .Y(n_576) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_536), .Y(n_639) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_539), .A2(n_615), .B(n_620), .C(n_631), .Y(n_614) );
OR2x2_ASAP7_75t_L g704 ( .A(n_539), .B(n_609), .Y(n_704) );
AND2x2_ASAP7_75t_L g706 ( .A(n_539), .B(n_572), .Y(n_706) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g546 ( .A(n_540), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g608 ( .A(n_540), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g646 ( .A(n_540), .B(n_613), .Y(n_646) );
OA33x2_ASAP7_75t_L g653 ( .A1(n_540), .A2(n_570), .A3(n_654), .B1(n_655), .B2(n_657), .B3(n_659), .Y(n_653) );
OR2x2_ASAP7_75t_L g664 ( .A(n_540), .B(n_649), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_540), .B(n_588), .Y(n_678) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g566 ( .A(n_542), .B(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_542), .A2(n_572), .B1(n_616), .B2(n_617), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_543), .B(n_623), .C(n_656), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_549), .A3(n_551), .B1(n_552), .B2(n_554), .C1(n_558), .C2(n_562), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g651 ( .A(n_547), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_548), .A2(n_563), .B(n_607), .C(n_610), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_549), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
NAND4xp25_ASAP7_75t_SL g670 ( .A(n_550), .B(n_579), .C(n_671), .D(n_673), .Y(n_670) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g560 ( .A(n_555), .Y(n_560) );
OR2x2_ASAP7_75t_L g605 ( .A(n_555), .B(n_557), .Y(n_605) );
AND2x2_ASAP7_75t_L g674 ( .A(n_556), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g679 ( .A(n_560), .B(n_674), .Y(n_679) );
BUFx2_ASAP7_75t_L g672 ( .A(n_561), .Y(n_672) );
INVx1_ASAP7_75t_SL g702 ( .A(n_562), .Y(n_702) );
AND2x4_ASAP7_75t_L g638 ( .A(n_563), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g691 ( .A(n_563), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_584), .C(n_606), .Y(n_564) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_SL g628 ( .A(n_570), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g696 ( .A1(n_570), .A2(n_697), .B(n_698), .C(n_707), .Y(n_696) );
OR2x2_ASAP7_75t_L g618 ( .A(n_571), .B(n_619), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .B1(n_580), .B2(n_581), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_575), .B(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_578), .B(n_635), .Y(n_717) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g692 ( .A(n_579), .B(n_580), .Y(n_692) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B1(n_594), .B2(n_598), .C1(n_599), .C2(n_604), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_587), .Y(n_598) );
AND2x2_ASAP7_75t_L g645 ( .A(n_588), .B(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_588), .A2(n_661), .B1(n_666), .B2(n_670), .Y(n_660) );
INVx2_ASAP7_75t_SL g713 ( .A(n_588), .Y(n_713) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g669 ( .A(n_593), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_593), .B(n_656), .Y(n_716) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g629 ( .A(n_597), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_599), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g667 ( .A(n_601), .Y(n_667) );
AND2x2_ASAP7_75t_SL g668 ( .A(n_602), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g710 ( .A(n_602), .B(n_639), .Y(n_710) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g635 ( .A(n_609), .Y(n_635) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g714 ( .A(n_612), .Y(n_714) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_613), .Y(n_658) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_625), .B(n_627), .C(n_630), .Y(n_620) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g665 ( .A(n_627), .Y(n_665) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_680), .C(n_696), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_660), .C(n_676), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B1(n_650), .B2(n_651), .C(n_653), .Y(n_643) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_662), .B(n_665), .Y(n_661) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g689 ( .A(n_675), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g697 ( .A(n_679), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_687), .Y(n_680) );
INVx2_ASAP7_75t_L g703 ( .A(n_682), .Y(n_703) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g694 ( .A(n_685), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_703), .B2(n_704), .C(n_705), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B1(n_715), .B2(n_717), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g734 ( .A(n_720), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_724), .A2(n_731), .B(n_738), .Y(n_730) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
BUFx3_ASAP7_75t_L g737 ( .A(n_727), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_729), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g731 ( .A(n_732), .B(n_735), .Y(n_731) );
CKINVDCx11_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g750 ( .A(n_742), .Y(n_750) );
INVx3_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_SL g743 ( .A(n_744), .B(n_745), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
endmodule