module fake_jpeg_14476_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_419;
wire n_133;
wire n_132;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_50),
.B(n_51),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_8),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_57),
.B(n_90),
.Y(n_110)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_23),
.B(n_8),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_32),
.B(n_17),
.Y(n_115)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_28),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_72),
.Y(n_125)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_8),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_14),
.Y(n_99)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_14),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_95),
.B(n_29),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_99),
.B(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_133),
.B1(n_41),
.B2(n_17),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_61),
.B(n_21),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_113),
.A2(n_10),
.B(n_14),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_115),
.B(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_20),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_73),
.A2(n_37),
.B1(n_27),
.B2(n_34),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_151),
.B1(n_89),
.B2(n_79),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_19),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_130),
.B(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_69),
.B1(n_70),
.B2(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_71),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_13),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_45),
.B(n_41),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_29),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_47),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_45),
.A2(n_37),
.B1(n_27),
.B2(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_32),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_158),
.A2(n_195),
.B1(n_196),
.B2(n_152),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_159),
.B(n_177),
.Y(n_226)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_81),
.B1(n_48),
.B2(n_66),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_192),
.B1(n_135),
.B2(n_147),
.Y(n_203)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_42),
.B1(n_30),
.B2(n_39),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_198),
.B1(n_177),
.B2(n_97),
.Y(n_211)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_39),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_128),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_115),
.B(n_139),
.C(n_142),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_167),
.A2(n_103),
.B(n_101),
.C(n_112),
.Y(n_237)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

BUFx4f_ASAP7_75t_SL g173 ( 
.A(n_136),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_173),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_176),
.Y(n_206)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_97),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_33),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_179),
.B(n_183),
.Y(n_214)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_107),
.B(n_33),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_181),
.B(n_191),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_30),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_186),
.B(n_15),
.Y(n_231)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_102),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_29),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_128),
.C(n_146),
.Y(n_215)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_92),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_53),
.B1(n_54),
.B2(n_68),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_194),
.B(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_123),
.A2(n_63),
.B1(n_83),
.B2(n_76),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_151),
.A2(n_77),
.B1(n_59),
.B2(n_15),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_116),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_199),
.B(n_148),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_159),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_116),
.B(n_125),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_215),
.B(n_234),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_205),
.B(n_189),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_211),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_215),
.B(n_188),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_228),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_122),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_186),
.Y(n_239)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_231),
.A2(n_237),
.B(n_173),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_179),
.B1(n_176),
.B2(n_183),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_239),
.B(n_252),
.Y(n_287)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_165),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_246),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_227),
.B1(n_223),
.B2(n_221),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_154),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_259),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_172),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_248),
.B(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_122),
.B1(n_147),
.B2(n_135),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_258),
.B1(n_264),
.B2(n_188),
.Y(n_277)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_233),
.B1(n_184),
.B2(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_254),
.B(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_204),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_189),
.B1(n_104),
.B2(n_180),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_214),
.B(n_170),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_157),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_262),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_266),
.B(n_267),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_178),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_206),
.B(n_199),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_134),
.B1(n_162),
.B2(n_175),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_265),
.B(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_206),
.A2(n_235),
.B1(n_214),
.B2(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_210),
.B(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_233),
.Y(n_294)
);

CKINVDCx6p67_ASAP7_75t_R g270 ( 
.A(n_241),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_273),
.C(n_278),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_241),
.A2(n_235),
.B1(n_219),
.B2(n_209),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_272),
.A2(n_274),
.B(n_299),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_171),
.C(n_168),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_227),
.B1(n_164),
.B2(n_106),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_277),
.B1(n_285),
.B2(n_301),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_187),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_282),
.B(n_297),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_245),
.A2(n_111),
.B1(n_185),
.B2(n_169),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_248),
.B(n_232),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_286),
.B(n_294),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_156),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_260),
.C(n_261),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_259),
.B(n_173),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_241),
.A2(n_219),
.B1(n_209),
.B2(n_208),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_269),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_267),
.A2(n_207),
.B1(n_229),
.B2(n_212),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_305),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_280),
.A2(n_239),
.B(n_267),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_304),
.A2(n_311),
.B(n_335),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_298),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_309),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_280),
.A2(n_266),
.B(n_256),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_312),
.B(n_271),
.Y(n_350)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_275),
.A2(n_253),
.B1(n_256),
.B2(n_261),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_318),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_294),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_321),
.Y(n_347)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_284),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_277),
.A2(n_254),
.B1(n_264),
.B2(n_238),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_291),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_287),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_249),
.B1(n_240),
.B2(n_243),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_242),
.B1(n_251),
.B2(n_255),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_281),
.A2(n_250),
.B1(n_258),
.B2(n_252),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_329),
.B1(n_330),
.B2(n_333),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_268),
.B(n_265),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g345 ( 
.A1(n_328),
.A2(n_293),
.B(n_286),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_281),
.A2(n_258),
.B1(n_247),
.B2(n_207),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_282),
.A2(n_221),
.B1(n_207),
.B2(n_229),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_296),
.A2(n_229),
.B1(n_198),
.B2(n_208),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_295),
.B1(n_285),
.B2(n_270),
.Y(n_358)
);

OAI22x1_ASAP7_75t_SL g333 ( 
.A1(n_274),
.A2(n_212),
.B1(n_218),
.B2(n_166),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_218),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_334),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_297),
.A2(n_225),
.B1(n_108),
.B2(n_193),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_331),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_364),
.Y(n_372)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_311),
.A2(n_272),
.B(n_293),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_355),
.B(n_357),
.Y(n_377)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_350),
.B(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_305),
.B(n_300),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_351),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_307),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_359),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_273),
.B(n_299),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_331),
.A2(n_307),
.B(n_321),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_358),
.A2(n_361),
.B1(n_333),
.B2(n_327),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_306),
.A2(n_270),
.B1(n_283),
.B2(n_288),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_320),
.B(n_283),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_360),
.B(n_362),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_270),
.B1(n_278),
.B2(n_160),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_225),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_334),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_325),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_324),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_318),
.A2(n_270),
.B(n_225),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_367),
.B(n_319),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_367),
.B(n_302),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_370),
.A2(n_378),
.B(n_397),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_310),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_371),
.B(n_376),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_360),
.B(n_322),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_381),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_310),
.C(n_312),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_375),
.C(n_390),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_346),
.C(n_328),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_302),
.Y(n_378)
);

NOR2x1_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

OA22x2_ASAP7_75t_L g381 ( 
.A1(n_352),
.A2(n_314),
.B1(n_323),
.B2(n_333),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_335),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_389),
.Y(n_398)
);

AND2x4_ASAP7_75t_SL g404 ( 
.A(n_383),
.B(n_394),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_354),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_385),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_339),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_356),
.B(n_316),
.Y(n_386)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_351),
.B(n_329),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_324),
.C(n_315),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_308),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_340),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_309),
.C(n_313),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_365),
.C(n_348),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_342),
.A2(n_319),
.B1(n_303),
.B2(n_330),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_396),
.A2(n_340),
.B(n_332),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_319),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_368),
.A2(n_358),
.B1(n_361),
.B2(n_347),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_399),
.A2(n_392),
.B1(n_403),
.B2(n_417),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_400),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_343),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_408),
.Y(n_434)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_372),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_407),
.Y(n_425)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_395),
.B(n_345),
.CI(n_347),
.CON(n_407),
.SN(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_353),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_339),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_413),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_375),
.B(n_365),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_415),
.B(n_419),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_416),
.A2(n_381),
.B1(n_388),
.B2(n_379),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_364),
.C(n_349),
.Y(n_419)
);

AOI21xp33_ASAP7_75t_L g420 ( 
.A1(n_394),
.A2(n_349),
.B(n_363),
.Y(n_420)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_420),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_363),
.C(n_344),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_423),
.C(n_15),
.Y(n_446)
);

FAx1_ASAP7_75t_SL g422 ( 
.A(n_390),
.B(n_380),
.CI(n_393),
.CON(n_422),
.SN(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_389),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_344),
.C(n_341),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_397),
.A2(n_341),
.B(n_338),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_SL g445 ( 
.A(n_424),
.B(n_10),
.C(n_12),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_412),
.A2(n_370),
.B1(n_378),
.B2(n_397),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_426),
.A2(n_422),
.B1(n_398),
.B2(n_400),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_408),
.B(n_378),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_439),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_380),
.B1(n_382),
.B2(n_370),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_432),
.A2(n_444),
.B1(n_132),
.B2(n_124),
.Y(n_467)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_435),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_414),
.A2(n_369),
.B1(n_381),
.B2(n_336),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_440),
.Y(n_454)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_438),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_419),
.A2(n_381),
.B1(n_338),
.B2(n_336),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_407),
.B(n_421),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_418),
.A2(n_388),
.B1(n_303),
.B2(n_225),
.Y(n_442)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_443),
.B(n_447),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_415),
.A2(n_303),
.B1(n_190),
.B2(n_155),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_445),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_406),
.Y(n_465)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_448),
.B(n_398),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_402),
.C(n_413),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_451),
.B(n_452),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_402),
.C(n_401),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_425),
.B(n_429),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_12),
.Y(n_483)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_455),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_435),
.B(n_441),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_459),
.A2(n_462),
.B(n_430),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_409),
.C(n_406),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_432),
.A2(n_426),
.B1(n_428),
.B2(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_465),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_467),
.B(n_444),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_434),
.C(n_428),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_468),
.B(n_470),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_434),
.C(n_446),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_471),
.B(n_473),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_457),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_472),
.B(n_474),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_440),
.C(n_439),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_481),
.C(n_483),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_442),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_477),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_131),
.B(n_12),
.Y(n_478)
);

AOI21xp33_ASAP7_75t_L g493 ( 
.A1(n_478),
.A2(n_11),
.B(n_10),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_456),
.A2(n_131),
.B1(n_12),
.B2(n_11),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_466),
.C(n_454),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_484),
.B(n_486),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_463),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_492),
.C(n_497),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_466),
.C(n_454),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_463),
.C(n_462),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_2),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_480),
.A2(n_449),
.B(n_458),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_491),
.A2(n_0),
.B(n_2),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_461),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_493),
.B(n_3),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_SL g496 ( 
.A(n_475),
.B(n_464),
.C(n_465),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_0),
.B(n_2),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_131),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_495),
.A2(n_480),
.B(n_474),
.Y(n_498)
);

AOI21x1_ASAP7_75t_SL g513 ( 
.A1(n_498),
.A2(n_503),
.B(n_504),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_11),
.C(n_2),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_499),
.B(n_505),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_484),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_500),
.B(n_494),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_506),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_488),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_507),
.A2(n_489),
.B1(n_485),
.B2(n_496),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_508),
.B(n_499),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_487),
.B(n_492),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_512),
.B(n_514),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_502),
.B(n_490),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_517),
.B(n_518),
.Y(n_519)
);

AOI21xp33_ASAP7_75t_L g517 ( 
.A1(n_513),
.A2(n_501),
.B(n_497),
.Y(n_517)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_509),
.A2(n_3),
.B(n_4),
.Y(n_518)
);

AO21x1_ASAP7_75t_SL g520 ( 
.A1(n_516),
.A2(n_511),
.B(n_5),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_511),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_519),
.B(n_5),
.C(n_6),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_522),
.A2(n_5),
.B(n_6),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_5),
.C(n_6),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_6),
.Y(n_525)
);


endmodule