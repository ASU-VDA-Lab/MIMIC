module fake_jpeg_14947_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_27),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_16),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_34),
.B1(n_19),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_31),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_34),
.B1(n_17),
.B2(n_30),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_19),
.B1(n_34),
.B2(n_17),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_68),
.A2(n_32),
.B1(n_25),
.B2(n_13),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_21),
.B1(n_24),
.B2(n_33),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_127)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_81),
.Y(n_143)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_99),
.Y(n_121)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_27),
.B1(n_29),
.B2(n_23),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_21),
.B1(n_24),
.B2(n_33),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_26),
.B1(n_36),
.B2(n_23),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_67),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_71),
.B(n_69),
.C(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_35),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_51),
.B(n_28),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_111),
.C(n_69),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_21),
.B1(n_24),
.B2(n_33),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_103),
.B1(n_109),
.B2(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_110),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_36),
.B1(n_31),
.B2(n_33),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_24),
.B1(n_15),
.B2(n_14),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_63),
.B1(n_61),
.B2(n_2),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_71),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_22),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_4),
.Y(n_139)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_35),
.B1(n_25),
.B2(n_32),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_35),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_49),
.B(n_32),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_0),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_32),
.B1(n_61),
.B2(n_70),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_25),
.B1(n_32),
.B2(n_2),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_112),
.A2(n_72),
.B1(n_63),
.B2(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_115),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_117),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_98),
.B1(n_108),
.B2(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_104),
.B1(n_101),
.B2(n_105),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_108),
.B1(n_88),
.B2(n_80),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_134),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_69),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_79),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_5),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_5),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_142),
.C(n_85),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_5),
.C(n_6),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_145),
.B(n_174),
.Y(n_193)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_143),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_165),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_SL g211 ( 
.A1(n_147),
.A2(n_153),
.B(n_10),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_88),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_154),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_79),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_171),
.C(n_127),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_117),
.B1(n_122),
.B2(n_138),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_98),
.B1(n_96),
.B2(n_86),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_156),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_100),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_77),
.B(n_97),
.C(n_78),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_159),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_82),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_161),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_83),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_77),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_76),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_78),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_90),
.B(n_7),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_167),
.A2(n_123),
.B(n_140),
.Y(n_182)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_124),
.A2(n_92),
.B1(n_91),
.B2(n_109),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_94),
.C(n_81),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_6),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_94),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_94),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_179),
.A2(n_189),
.B1(n_192),
.B2(n_174),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_184),
.C(n_209),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_185),
.B(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_144),
.B1(n_118),
.B2(n_140),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_144),
.B1(n_126),
.B2(n_133),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_125),
.B(n_126),
.C(n_8),
.D(n_9),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_202),
.B(n_161),
.C(n_151),
.D(n_12),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_133),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_6),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_157),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_7),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_7),
.B(n_8),
.Y(n_197)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_8),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_148),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_148),
.B(n_162),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_211),
.B1(n_190),
.B2(n_209),
.Y(n_238)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_9),
.C(n_10),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_149),
.C(n_145),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_221),
.C(n_224),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_158),
.B(n_176),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_222),
.B(n_223),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_171),
.C(n_175),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_175),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_164),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_228),
.C(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_166),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_169),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_170),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_229),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_173),
.B(n_172),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_240),
.B(n_204),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_235),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_12),
.B(n_182),
.C(n_178),
.Y(n_235)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_185),
.A2(n_191),
.B(n_183),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_192),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_200),
.B1(n_188),
.B2(n_201),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_195),
.C(n_189),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_203),
.A2(n_197),
.B(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_243),
.B1(n_253),
.B2(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_265),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_181),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_200),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_207),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_231),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_188),
.C(n_198),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_263),
.C(n_224),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_230),
.A2(n_198),
.B1(n_239),
.B2(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_261),
.B1(n_223),
.B2(n_220),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_229),
.B1(n_221),
.B2(n_228),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_217),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_213),
.C(n_225),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_238),
.B1(n_215),
.B2(n_219),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_268),
.C(n_270),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_224),
.C(n_218),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_214),
.C(n_240),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_214),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_278),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_222),
.C(n_237),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_285),
.C(n_286),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_237),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_235),
.B(n_237),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_280),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_235),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_245),
.A2(n_220),
.B1(n_223),
.B2(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_261),
.C(n_260),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_256),
.C(n_246),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_243),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_294),
.C(n_295),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_274),
.C(n_286),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_242),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_245),
.B1(n_250),
.B2(n_265),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_271),
.B1(n_266),
.B2(n_273),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_249),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_254),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_303),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_290),
.B1(n_280),
.B2(n_300),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_276),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_315),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_282),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_312),
.C(n_316),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_298),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_270),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_266),
.B1(n_246),
.B2(n_256),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_294),
.B1(n_303),
.B2(n_288),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_257),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_293),
.A2(n_259),
.B(n_241),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_287),
.B(n_259),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_298),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_248),
.Y(n_319)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_321),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_288),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_312),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_329),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_307),
.B(n_317),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_324),
.B(n_327),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_323),
.A2(n_322),
.B(n_318),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_336),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_308),
.C(n_307),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_333),
.A2(n_320),
.B(n_330),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_332),
.B(n_334),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_341),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_345),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_342),
.B(n_335),
.Y(n_347)
);


endmodule