module fake_jpeg_1044_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_18),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_63),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_60),
.B(n_51),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_61),
.B(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_71),
.Y(n_89)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_57),
.B1(n_66),
.B2(n_50),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_64),
.B1(n_49),
.B2(n_51),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_64),
.B1(n_84),
.B2(n_54),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_49),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_65),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_65),
.B(n_59),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_5),
.C(n_6),
.Y(n_117)
);

AO21x1_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_0),
.B(n_1),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_72),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_64),
.B1(n_70),
.B2(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_54),
.B1(n_57),
.B2(n_47),
.Y(n_108)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_108),
.B1(n_112),
.B2(n_116),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_66),
.B1(n_60),
.B2(n_47),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_113),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_61),
.A3(n_57),
.B1(n_52),
.B2(n_3),
.Y(n_110)
);

XOR2x2_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_8),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_61),
.B1(n_52),
.B2(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_118),
.B1(n_8),
.B2(n_9),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_14),
.B(n_15),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_15),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_88),
.B1(n_97),
.B2(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_7),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_139),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_44),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_133),
.C(n_137),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_110),
.B(n_115),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_26),
.C(n_42),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_25),
.C(n_40),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_21),
.CI(n_22),
.CON(n_148),
.SN(n_148)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_14),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_43),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_20),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_16),
.B(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_123),
.C(n_135),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_24),
.B(n_29),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_151),
.B1(n_138),
.B2(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_154),
.B(n_157),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_135),
.C(n_128),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.C(n_160),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_130),
.C(n_37),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_150),
.C(n_156),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_167),
.B1(n_161),
.B2(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_165),
.B(n_143),
.C(n_140),
.D(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_141),
.C(n_149),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_151),
.Y(n_174)
);


endmodule