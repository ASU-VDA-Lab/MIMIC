module real_aes_7788_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_754;
wire n_182;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g125 ( .A(n_0), .Y(n_125) );
INVx1_ASAP7_75t_L g522 ( .A(n_1), .Y(n_522) );
INVx1_ASAP7_75t_L g159 ( .A(n_2), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_3), .A2(n_747), .B1(n_750), .B2(n_751), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_3), .Y(n_751) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_4), .A2(n_21), .B1(n_128), .B2(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_4), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_5), .A2(n_39), .B1(n_184), .B2(n_478), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g203 ( .A1(n_6), .A2(n_175), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_7), .B(n_173), .Y(n_533) );
AND2x6_ASAP7_75t_L g152 ( .A(n_8), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_9), .A2(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_10), .B(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g209 ( .A(n_11), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_12), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_14), .B(n_165), .Y(n_486) );
INVx1_ASAP7_75t_L g263 ( .A(n_15), .Y(n_263) );
INVx1_ASAP7_75t_L g516 ( .A(n_16), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_17), .B(n_140), .Y(n_538) );
AO32x2_ASAP7_75t_L g505 ( .A1(n_18), .A2(n_139), .A3(n_173), .B1(n_480), .B2(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_19), .B(n_184), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_20), .B(n_180), .Y(n_251) );
INVxp67_ASAP7_75t_L g128 ( .A(n_21), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_21), .B(n_140), .Y(n_524) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_22), .A2(n_32), .B1(n_451), .B2(n_452), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_22), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_23), .A2(n_52), .B1(n_184), .B2(n_478), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_24), .B(n_175), .Y(n_220) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_25), .A2(n_80), .B1(n_165), .B2(n_184), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_26), .B(n_184), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_27), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_28), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_30), .B(n_170), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_31), .B(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_32), .Y(n_452) );
INVx1_ASAP7_75t_L g198 ( .A(n_33), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_34), .B(n_170), .Y(n_503) );
INVx2_ASAP7_75t_L g150 ( .A(n_35), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_36), .B(n_184), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_37), .B(n_170), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_38), .A2(n_152), .B(n_155), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g196 ( .A(n_41), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_42), .B(n_163), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_43), .B(n_456), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_44), .A2(n_460), .B1(n_742), .B2(n_743), .C1(n_752), .C2(n_754), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_45), .B(n_184), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_46), .A2(n_90), .B1(n_227), .B2(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_47), .B(n_184), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_48), .B(n_184), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_49), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_50), .B(n_521), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_51), .B(n_175), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_53), .A2(n_64), .B1(n_165), .B2(n_184), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_54), .A2(n_155), .B1(n_165), .B2(n_194), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_55), .A2(n_105), .B1(n_114), .B2(n_759), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_56), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_57), .B(n_184), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_58), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_59), .B(n_184), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_60), .A2(n_183), .B(n_207), .C(n_208), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_61), .Y(n_254) );
INVx1_ASAP7_75t_L g205 ( .A(n_62), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_63), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_63), .Y(n_744) );
INVx1_ASAP7_75t_L g153 ( .A(n_65), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_66), .B(n_184), .Y(n_523) );
INVx1_ASAP7_75t_L g143 ( .A(n_67), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_68), .Y(n_119) );
AO32x2_ASAP7_75t_L g475 ( .A1(n_69), .A2(n_173), .A3(n_232), .B1(n_476), .B2(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g555 ( .A(n_70), .Y(n_555) );
INVx1_ASAP7_75t_L g498 ( .A(n_71), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_72), .A2(n_79), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_72), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_73), .A2(n_180), .B(n_181), .C(n_183), .Y(n_179) );
INVxp67_ASAP7_75t_L g182 ( .A(n_74), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_75), .B(n_165), .Y(n_499) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_77), .Y(n_201) );
INVx1_ASAP7_75t_L g247 ( .A(n_78), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_79), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_81), .A2(n_152), .B(n_155), .C(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_82), .B(n_478), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_83), .B(n_165), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_84), .B(n_160), .Y(n_223) );
INVx2_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_86), .B(n_180), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_87), .B(n_165), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_88), .A2(n_152), .B(n_155), .C(n_158), .Y(n_154) );
INVx2_ASAP7_75t_L g108 ( .A(n_89), .Y(n_108) );
OR2x2_ASAP7_75t_L g122 ( .A(n_89), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g463 ( .A(n_89), .B(n_124), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_91), .A2(n_103), .B1(n_165), .B2(n_166), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_92), .B(n_170), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_93), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_94), .A2(n_152), .B(n_155), .C(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_95), .Y(n_242) );
INVx1_ASAP7_75t_L g178 ( .A(n_96), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_97), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_98), .B(n_160), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_99), .B(n_165), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_100), .B(n_173), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_102), .A2(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_106), .Y(n_760) );
OR2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_112), .Y(n_106) );
OR2x2_ASAP7_75t_L g466 ( .A(n_108), .B(n_124), .Y(n_466) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_108), .B(n_123), .Y(n_756) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g124 ( .A(n_113), .B(n_125), .Y(n_124) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_458), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g758 ( .A(n_118), .Y(n_758) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_126), .B(n_455), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_122), .Y(n_457) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_131), .B2(n_454), .Y(n_126) );
INVx1_ASAP7_75t_L g454 ( .A(n_127), .Y(n_454) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_449), .B1(n_450), .B2(n_453), .Y(n_131) );
INVx2_ASAP7_75t_L g453 ( .A(n_132), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_132), .A2(n_461), .B1(n_468), .B2(n_753), .Y(n_752) );
OR4x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_338), .C(n_398), .D(n_425), .Y(n_132) );
NAND4xp25_ASAP7_75t_SL g133 ( .A(n_134), .B(n_286), .C(n_317), .D(n_334), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_211), .B(n_213), .C(n_266), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_189), .Y(n_135) );
INVx1_ASAP7_75t_L g328 ( .A(n_136), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_136), .A2(n_369), .B1(n_417), .B2(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_171), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_137), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g279 ( .A(n_137), .B(n_191), .Y(n_279) );
AND2x2_ASAP7_75t_L g321 ( .A(n_137), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_137), .B(n_212), .Y(n_333) );
INVx1_ASAP7_75t_L g373 ( .A(n_137), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_137), .B(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g301 ( .A(n_138), .B(n_191), .Y(n_301) );
INVx3_ASAP7_75t_L g305 ( .A(n_138), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_138), .B(n_363), .Y(n_362) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_167), .Y(n_138) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_139), .A2(n_192), .B(n_200), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_139), .B(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g228 ( .A(n_139), .Y(n_228) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_141), .B(n_142), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_154), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_147), .A2(n_185), .B1(n_193), .B2(n_199), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_147), .A2(n_247), .B(n_248), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AND2x4_ASAP7_75t_L g175 ( .A(n_148), .B(n_152), .Y(n_175) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g521 ( .A(n_149), .Y(n_521) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx3_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
INVx4_ASAP7_75t_SL g185 ( .A(n_152), .Y(n_185) );
BUFx3_ASAP7_75t_L g480 ( .A(n_152), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_152), .A2(n_484), .B(n_488), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_152), .A2(n_497), .B(n_500), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_152), .A2(n_515), .B(n_519), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_152), .A2(n_527), .B(n_530), .Y(n_526) );
INVx5_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
BUFx3_ASAP7_75t_L g227 ( .A(n_156), .Y(n_227) );
INVx1_ASAP7_75t_L g478 ( .A(n_156), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .C(n_164), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_SL g497 ( .A1(n_160), .A2(n_183), .B(n_498), .C(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g508 ( .A(n_160), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_160), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_160), .A2(n_552), .B(n_553), .Y(n_551) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_161), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_161), .B(n_209), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g476 ( .A1(n_161), .A2(n_163), .B1(n_477), .B2(n_479), .Y(n_476) );
INVx2_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
INVx4_ASAP7_75t_L g238 ( .A(n_163), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_163), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_163), .A2(n_508), .B1(n_541), .B2(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_164), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_169), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_169), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g232 ( .A(n_170), .Y(n_232) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_170), .A2(n_256), .B(n_265), .Y(n_255) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_170), .A2(n_483), .B(n_491), .Y(n_482) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_170), .A2(n_496), .B(n_503), .Y(n_495) );
AND2x2_ASAP7_75t_L g392 ( .A(n_171), .B(n_202), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_171), .B(n_305), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_171), .B(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g212 ( .A(n_172), .B(n_191), .Y(n_212) );
INVx1_ASAP7_75t_L g274 ( .A(n_172), .Y(n_274) );
BUFx2_ASAP7_75t_L g278 ( .A(n_172), .Y(n_278) );
AND2x2_ASAP7_75t_L g322 ( .A(n_172), .B(n_190), .Y(n_322) );
OR2x2_ASAP7_75t_L g361 ( .A(n_172), .B(n_190), .Y(n_361) );
AND2x2_ASAP7_75t_L g386 ( .A(n_172), .B(n_202), .Y(n_386) );
AND2x2_ASAP7_75t_L g445 ( .A(n_172), .B(n_275), .Y(n_445) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_186), .Y(n_172) );
INVx4_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_173), .A2(n_526), .B(n_533), .Y(n_525) );
BUFx2_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_185), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_177), .A2(n_185), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_177), .A2(n_185), .B(n_259), .C(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g487 ( .A(n_180), .Y(n_487) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_187), .A2(n_203), .B(n_210), .Y(n_202) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_SL g229 ( .A(n_188), .B(n_230), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_188), .B(n_480), .C(n_540), .Y(n_539) );
AO21x1_ASAP7_75t_L g586 ( .A1(n_188), .A2(n_540), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g420 ( .A(n_189), .Y(n_420) );
OR2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_202), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_190), .B(n_202), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_190), .B(n_305), .Y(n_316) );
BUFx2_ASAP7_75t_L g327 ( .A(n_190), .Y(n_327) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g349 ( .A(n_191), .B(n_202), .Y(n_349) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_191), .Y(n_404) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
INVx2_ASAP7_75t_L g197 ( .A(n_195), .Y(n_197) );
INVx4_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_202), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_SL g275 ( .A(n_202), .Y(n_275) );
BUFx2_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
INVx2_ASAP7_75t_L g319 ( .A(n_202), .Y(n_319) );
AND2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_305), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_207), .A2(n_489), .B(n_490), .Y(n_488) );
O2A1O1Ixp5_ASAP7_75t_L g554 ( .A1(n_207), .A2(n_520), .B(n_555), .C(n_556), .Y(n_554) );
AOI321xp33_ASAP7_75t_L g400 ( .A1(n_211), .A2(n_401), .A3(n_402), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_212), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_212), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g394 ( .A(n_212), .B(n_373), .Y(n_394) );
AND2x2_ASAP7_75t_L g427 ( .A(n_212), .B(n_319), .Y(n_427) );
INVx1_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_243), .Y(n_214) );
OR2x2_ASAP7_75t_L g329 ( .A(n_215), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_231), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g281 ( .A(n_218), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_218), .B(n_245), .Y(n_291) );
AND2x2_ASAP7_75t_L g296 ( .A(n_218), .B(n_271), .Y(n_296) );
INVx1_ASAP7_75t_L g313 ( .A(n_218), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_218), .B(n_294), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_218), .B(n_270), .Y(n_337) );
OR2x2_ASAP7_75t_L g369 ( .A(n_218), .B(n_358), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_218), .B(n_282), .Y(n_408) );
AND2x2_ASAP7_75t_L g442 ( .A(n_218), .B(n_268), .Y(n_442) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B(n_228), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_225), .A2(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx1_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_228), .A2(n_514), .B(n_524), .Y(n_513) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_228), .A2(n_550), .B(n_557), .Y(n_549) );
INVx1_ASAP7_75t_L g269 ( .A(n_231), .Y(n_269) );
INVx2_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
AND2x2_ASAP7_75t_L g324 ( .A(n_231), .B(n_295), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_231), .B(n_271), .Y(n_346) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_241), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_239), .Y(n_235) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g430 ( .A(n_244), .B(n_281), .Y(n_430) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_255), .Y(n_244) );
INVx2_ASAP7_75t_L g271 ( .A(n_245), .Y(n_271) );
AND2x2_ASAP7_75t_L g424 ( .A(n_245), .B(n_284), .Y(n_424) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B(n_253), .Y(n_245) );
AND2x2_ASAP7_75t_L g270 ( .A(n_255), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
INVx1_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_261), .B(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_261), .A2(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g518 ( .A(n_261), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_272), .B1(n_276), .B2(n_280), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_267), .A2(n_385), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g331 ( .A(n_271), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_271), .B(n_284), .Y(n_358) );
INVx1_ASAP7_75t_L g374 ( .A(n_271), .Y(n_374) );
AND2x2_ASAP7_75t_L g315 ( .A(n_273), .B(n_316), .Y(n_315) );
INVx3_ASAP7_75t_SL g354 ( .A(n_273), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_273), .B(n_279), .Y(n_431) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g440 ( .A(n_276), .Y(n_440) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_277), .B(n_373), .Y(n_415) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx3_ASAP7_75t_SL g320 ( .A(n_279), .Y(n_320) );
NAND2x1_ASAP7_75t_SL g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g341 ( .A(n_281), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g348 ( .A(n_281), .B(n_285), .Y(n_348) );
AND2x2_ASAP7_75t_L g353 ( .A(n_281), .B(n_294), .Y(n_353) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_281), .Y(n_402) );
OAI311xp33_ASAP7_75t_L g425 ( .A1(n_282), .A2(n_426), .A3(n_428), .B1(n_429), .C1(n_439), .Y(n_425) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g438 ( .A(n_283), .B(n_311), .Y(n_438) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g294 ( .A(n_284), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g342 ( .A(n_284), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g397 ( .A(n_284), .Y(n_397) );
INVx1_ASAP7_75t_L g290 ( .A(n_285), .Y(n_290) );
INVx1_ASAP7_75t_L g310 ( .A(n_285), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_285), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g343 ( .A(n_285), .Y(n_343) );
AOI221xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_289), .B1(n_297), .B2(n_302), .C(n_307), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_292), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx4_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
AND2x2_ASAP7_75t_L g405 ( .A(n_291), .B(n_324), .Y(n_405) );
AND2x2_ASAP7_75t_L g412 ( .A(n_291), .B(n_294), .Y(n_412) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_294), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_299), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g448 ( .A(n_301), .B(n_392), .Y(n_448) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g433 ( .A(n_305), .B(n_361), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_306), .A2(n_399), .B(n_400), .C(n_413), .Y(n_398) );
AOI21xp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_312), .B(n_314), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g377 ( .A(n_311), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_312), .A2(n_407), .B1(n_408), .B2(n_409), .C(n_410), .Y(n_406) );
AND2x2_ASAP7_75t_L g383 ( .A(n_313), .B(n_324), .Y(n_383) );
AND2x2_ASAP7_75t_L g436 ( .A(n_313), .B(n_331), .Y(n_436) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_316), .B(n_354), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_323), .C(n_325), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g364 ( .A(n_319), .B(n_322), .Y(n_364) );
OR2x2_ASAP7_75t_L g407 ( .A(n_319), .B(n_361), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_320), .B(n_386), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_320), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g351 ( .A(n_321), .Y(n_351) );
INVx1_ASAP7_75t_L g417 ( .A(n_324), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_332), .B2(n_333), .Y(n_325) );
INVx1_ASAP7_75t_L g340 ( .A(n_326), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_327), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_328), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g389 ( .A(n_330), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_331), .B(n_417), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_332), .A2(n_391), .B1(n_393), .B2(n_395), .Y(n_390) );
INVx1_ASAP7_75t_L g399 ( .A(n_335), .Y(n_399) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g441 ( .A(n_336), .B(n_436), .Y(n_441) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_337), .A2(n_371), .B1(n_374), .B2(n_375), .C1(n_378), .C2(n_379), .Y(n_370) );
NAND4xp25_ASAP7_75t_SL g338 ( .A(n_339), .B(n_359), .C(n_370), .D(n_382), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_344), .B2(n_349), .C(n_350), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_342), .B(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_344), .A2(n_414), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_413) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_348), .B(n_357), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_349), .A2(n_411), .B(n_412), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_354), .B2(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_365), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_373), .B(n_392), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_373), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_377), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g409 ( .A(n_381), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_387), .B2(n_389), .C(n_390), .Y(n_382) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI222xp33_ASAP7_75t_L g429 ( .A1(n_392), .A2(n_430), .B1(n_431), .B2(n_432), .C1(n_434), .C2(n_437), .Y(n_429) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_396), .B(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g428 ( .A(n_402), .Y(n_428) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp33_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_442), .B2(n_443), .C(n_446), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_453), .A2(n_461), .B1(n_464), .B2(n_467), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_455), .B(n_459), .C(n_757), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g753 ( .A(n_465), .Y(n_753) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND3x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_662), .C(n_710), .Y(n_469) );
NOR4xp25_ASAP7_75t_L g470 ( .A(n_471), .B(n_590), .C(n_635), .D(n_649), .Y(n_470) );
OAI311xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_510), .A3(n_534), .B1(n_543), .C1(n_558), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
OAI21xp33_ASAP7_75t_L g543 ( .A1(n_473), .A2(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g651 ( .A(n_473), .B(n_578), .Y(n_651) );
AND2x2_ASAP7_75t_L g708 ( .A(n_473), .B(n_594), .Y(n_708) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g601 ( .A(n_474), .B(n_504), .Y(n_601) );
AND2x2_ASAP7_75t_L g658 ( .A(n_474), .B(n_606), .Y(n_658) );
INVx1_ASAP7_75t_L g699 ( .A(n_474), .Y(n_699) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_475), .Y(n_567) );
AND2x2_ASAP7_75t_L g608 ( .A(n_475), .B(n_504), .Y(n_608) );
AND2x2_ASAP7_75t_L g612 ( .A(n_475), .B(n_505), .Y(n_612) );
INVx1_ASAP7_75t_L g624 ( .A(n_475), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_480), .A2(n_551), .B(n_554), .Y(n_550) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
AND2x2_ASAP7_75t_L g545 ( .A(n_482), .B(n_504), .Y(n_545) );
INVx2_ASAP7_75t_L g579 ( .A(n_482), .Y(n_579) );
AND2x2_ASAP7_75t_L g594 ( .A(n_482), .B(n_505), .Y(n_594) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_482), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_482), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g614 ( .A(n_482), .B(n_577), .Y(n_614) );
INVx1_ASAP7_75t_L g626 ( .A(n_482), .Y(n_626) );
INVx1_ASAP7_75t_L g667 ( .A(n_482), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_482), .B(n_567), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_487), .Y(n_484) );
NOR2xp67_ASAP7_75t_L g492 ( .A(n_493), .B(n_504), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g544 ( .A(n_494), .B(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_494), .Y(n_572) );
AND2x2_ASAP7_75t_SL g625 ( .A(n_494), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g629 ( .A(n_494), .B(n_504), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_494), .B(n_624), .Y(n_687) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g577 ( .A(n_495), .Y(n_577) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_495), .Y(n_593) );
OR2x2_ASAP7_75t_L g666 ( .A(n_495), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g573 ( .A(n_505), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_505), .B(n_579), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_508), .A2(n_520), .B(n_522), .C(n_523), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_508), .A2(n_531), .B(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_510), .B(n_561), .Y(n_724) );
INVx1_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g694 ( .A(n_511), .B(n_536), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_525), .Y(n_511) );
AND2x2_ASAP7_75t_L g570 ( .A(n_512), .B(n_561), .Y(n_570) );
INVx2_ASAP7_75t_L g582 ( .A(n_512), .Y(n_582) );
AND2x2_ASAP7_75t_L g616 ( .A(n_512), .B(n_564), .Y(n_616) );
AND2x2_ASAP7_75t_L g683 ( .A(n_512), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_513), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g563 ( .A(n_513), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g603 ( .A(n_513), .B(n_525), .Y(n_603) );
AND2x2_ASAP7_75t_L g620 ( .A(n_513), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g546 ( .A(n_525), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g564 ( .A(n_525), .Y(n_564) );
AND2x2_ASAP7_75t_L g569 ( .A(n_525), .B(n_549), .Y(n_569) );
AND2x2_ASAP7_75t_L g642 ( .A(n_525), .B(n_621), .Y(n_642) );
AND2x2_ASAP7_75t_L g707 ( .A(n_525), .B(n_697), .Y(n_707) );
OAI311xp33_ASAP7_75t_L g590 ( .A1(n_534), .A2(n_591), .A3(n_595), .B1(n_597), .C1(n_617), .Y(n_590) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g602 ( .A(n_535), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g661 ( .A(n_535), .B(n_569), .Y(n_661) );
AND2x2_ASAP7_75t_L g735 ( .A(n_535), .B(n_616), .Y(n_735) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_536), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g670 ( .A(n_536), .Y(n_670) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_537), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g690 ( .A(n_537), .B(n_564), .Y(n_690) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g587 ( .A(n_538), .Y(n_587) );
AND2x2_ASAP7_75t_L g565 ( .A(n_545), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g618 ( .A(n_545), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g698 ( .A(n_545), .B(n_699), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_546), .A2(n_578), .B1(n_598), .B2(n_602), .C(n_604), .Y(n_597) );
INVx1_ASAP7_75t_L g722 ( .A(n_547), .Y(n_722) );
OR2x2_ASAP7_75t_L g688 ( .A(n_548), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g583 ( .A(n_549), .B(n_564), .Y(n_583) );
OR2x2_ASAP7_75t_L g585 ( .A(n_549), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
INVx2_ASAP7_75t_L g621 ( .A(n_549), .Y(n_621) );
AND2x2_ASAP7_75t_L g648 ( .A(n_549), .B(n_586), .Y(n_648) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_549), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_565), .B1(n_568), .B2(n_571), .C(n_574), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
AND2x2_ASAP7_75t_L g659 ( .A(n_561), .B(n_569), .Y(n_659) );
AND2x2_ASAP7_75t_L g709 ( .A(n_561), .B(n_563), .Y(n_709) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g596 ( .A(n_563), .B(n_567), .Y(n_596) );
AND2x2_ASAP7_75t_L g675 ( .A(n_563), .B(n_648), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_564), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g634 ( .A(n_564), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g644 ( .A1(n_565), .A2(n_645), .B(n_647), .Y(n_644) );
OR2x2_ASAP7_75t_L g588 ( .A(n_566), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g654 ( .A(n_566), .B(n_614), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_566), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g631 ( .A(n_567), .B(n_600), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_567), .B(n_714), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_568), .B(n_594), .Y(n_704) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g627 ( .A(n_569), .B(n_582), .Y(n_627) );
INVx1_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_580), .B1(n_584), .B2(n_588), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g606 ( .A(n_577), .Y(n_606) );
INVx1_ASAP7_75t_L g619 ( .A(n_577), .Y(n_619) );
INVx1_ASAP7_75t_L g589 ( .A(n_578), .Y(n_589) );
AND2x2_ASAP7_75t_L g660 ( .A(n_578), .B(n_606), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_578), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
OR2x2_ASAP7_75t_L g584 ( .A(n_581), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_581), .B(n_697), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g728 ( .A(n_581), .B(n_729), .Y(n_728) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g731 ( .A(n_583), .B(n_683), .Y(n_731) );
INVx1_ASAP7_75t_SL g697 ( .A(n_585), .Y(n_697) );
AND2x2_ASAP7_75t_L g637 ( .A(n_586), .B(n_621), .Y(n_637) );
INVx1_ASAP7_75t_L g684 ( .A(n_586), .Y(n_684) );
OAI222xp33_ASAP7_75t_L g725 ( .A1(n_591), .A2(n_681), .B1(n_726), .B2(n_727), .C1(n_730), .C2(n_732), .Y(n_725) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g646 ( .A(n_593), .Y(n_646) );
AND2x2_ASAP7_75t_L g657 ( .A(n_594), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_594), .B(n_699), .Y(n_726) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_596), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g701 ( .A(n_598), .Y(n_701) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g639 ( .A(n_601), .Y(n_639) );
AND2x2_ASAP7_75t_L g718 ( .A(n_601), .B(n_679), .Y(n_718) );
AND2x2_ASAP7_75t_L g741 ( .A(n_601), .B(n_625), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_603), .B(n_637), .Y(n_636) );
OAI32xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .A3(n_609), .B1(n_611), .B2(n_615), .Y(n_604) );
BUFx2_ASAP7_75t_L g679 ( .A(n_606), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_607), .B(n_625), .Y(n_706) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g713 ( .A(n_608), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g702 ( .A(n_609), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g673 ( .A(n_612), .B(n_646), .Y(n_673) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OAI221xp5_ASAP7_75t_SL g635 ( .A1(n_614), .A2(n_636), .B1(n_638), .B2(n_640), .C(n_644), .Y(n_635) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g647 ( .A(n_616), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g653 ( .A(n_616), .B(n_637), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_622), .B2(n_627), .C(n_628), .Y(n_617) );
INVx1_ASAP7_75t_L g736 ( .A(n_618), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_619), .B(n_713), .Y(n_712) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_620), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_625), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g691 ( .A(n_625), .Y(n_691) );
BUFx3_ASAP7_75t_L g714 ( .A(n_626), .Y(n_714) );
INVx1_ASAP7_75t_SL g655 ( .A(n_627), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_627), .B(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_630), .B(n_632), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_629), .A2(n_730), .B1(n_734), .B2(n_736), .C(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g676 ( .A(n_634), .B(n_637), .Y(n_676) );
INVx1_ASAP7_75t_L g740 ( .A(n_634), .Y(n_740) );
INVx2_ASAP7_75t_L g729 ( .A(n_637), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_637), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g682 ( .A(n_642), .B(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_652), .B1(n_654), .B2(n_655), .C(n_656), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_658), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_719) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_661), .A2(n_738), .B(n_741), .Y(n_737) );
NOR4xp25_ASAP7_75t_SL g662 ( .A(n_663), .B(n_671), .C(n_680), .D(n_700), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_677), .B2(n_678), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g716 ( .A(n_676), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B1(n_688), .B2(n_691), .C(n_692), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g703 ( .A(n_683), .Y(n_703) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_695), .B(n_698), .Y(n_692) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_704), .C(n_705), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_705) );
CKINVDCx14_ASAP7_75t_R g715 ( .A(n_709), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_725), .C(n_733), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B1(n_716), .B2(n_717), .C(n_719), .Y(n_711) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g750 ( .A(n_747), .Y(n_750) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx3_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
endmodule