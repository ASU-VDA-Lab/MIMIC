module fake_netlist_5_76_n_1949 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1949);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1949;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_191),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_39),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_87),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_37),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_73),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_50),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_31),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_83),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_108),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_25),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_103),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_149),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_93),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_65),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_115),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_181),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_124),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_3),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_88),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_195),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_155),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_138),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_94),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_39),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_150),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_131),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_156),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_0),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_119),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_30),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_67),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_172),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_46),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_86),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_122),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_13),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_78),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_178),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_146),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_110),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_49),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_152),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_68),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_82),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_62),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_90),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_25),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_153),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_70),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_187),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_72),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_170),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_6),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_30),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_81),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_157),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_48),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_40),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_43),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_16),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_133),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_106),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_111),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_80),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_189),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_143),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_60),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_184),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_89),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_44),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_154),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_116),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_75),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_185),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_117),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_5),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_140),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_35),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_137),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_59),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_139),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_100),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_57),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_23),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_28),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_99),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_190),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_56),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_69),
.Y(n_324)
);

BUFx2_ASAP7_75t_SL g325 ( 
.A(n_34),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_102),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_38),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_3),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_41),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_120),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_76),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_162),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_42),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_186),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_92),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_85),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_144),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_53),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_31),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_33),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_193),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_77),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_126),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_35),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_28),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_97),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_98),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_17),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_42),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_129),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_96),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_12),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_52),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_183),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_79),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_180),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_56),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_66),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_7),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_91),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_60),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_6),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_71),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_20),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_47),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_159),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_4),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_16),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_161),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_4),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_9),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_27),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_173),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_171),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_36),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_168),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_128),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_52),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_7),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_125),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_182),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_57),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_8),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_34),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_55),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_132),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_53),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_2),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_269),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_269),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_269),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_269),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_225),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_234),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_236),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_225),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_272),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_272),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_301),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_237),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_251),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_301),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_304),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_304),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_204),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_204),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_239),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_229),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_206),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_241),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_210),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_336),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_317),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_366),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_294),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_213),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_240),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_362),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_244),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_366),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_214),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_226),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_207),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_291),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_245),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_324),
.Y(n_435)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_206),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_255),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_250),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_258),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_266),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_267),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_251),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_263),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_247),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_331),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_249),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_285),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_290),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_216),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_291),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_295),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_253),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_310),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_257),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_338),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_259),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_260),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_209),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_339),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_291),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_209),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_359),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_262),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_264),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_270),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_363),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_271),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_273),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_275),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_277),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_319),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_246),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_319),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_282),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_337),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_287),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_340),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_340),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_198),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_288),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_354),
.Y(n_487)
);

INVxp33_ASAP7_75t_SL g488 ( 
.A(n_232),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_232),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_354),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_296),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_201),
.Y(n_492)
);

BUFx12f_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_398),
.B(n_375),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_403),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_392),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_414),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_375),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_200),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_413),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_393),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_196),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_425),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_394),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_481),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_395),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_318),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_449),
.B(n_230),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_395),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_449),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_396),
.A2(n_220),
.B(n_216),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_396),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_429),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_427),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_417),
.A2(n_278),
.B1(n_286),
.B2(n_345),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_404),
.B(n_263),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g531 ( 
.A(n_424),
.B(n_220),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_442),
.B(n_263),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_196),
.Y(n_535)
);

XNOR2x2_ASAP7_75t_R g536 ( 
.A(n_450),
.B(n_420),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_444),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_415),
.B(n_197),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_R g540 ( 
.A(n_436),
.B(n_197),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_421),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_399),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_399),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_421),
.B(n_199),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_422),
.Y(n_547)
);

BUFx8_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_400),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_458),
.B(n_256),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_400),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_423),
.A2(n_435),
.B1(n_426),
.B2(n_445),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_401),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_434),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_454),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_422),
.B(n_256),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_428),
.B(n_203),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_457),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_446),
.B(n_361),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_428),
.B(n_478),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_401),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_402),
.B(n_230),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_437),
.B(n_447),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_402),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_405),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_552),
.A2(n_323),
.B1(n_364),
.B2(n_361),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_531),
.B(n_452),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_494),
.B(n_456),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_495),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_498),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_500),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_498),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_507),
.A2(n_519),
.B1(n_557),
.B2(n_506),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_509),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_531),
.B(n_464),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_531),
.B(n_465),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_509),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_552),
.A2(n_372),
.B1(n_373),
.B2(n_364),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_510),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_497),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_502),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_521),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_539),
.B(n_474),
.C(n_473),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_521),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_552),
.B(n_475),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_496),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_540),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_493),
.B(n_325),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_548),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_493),
.B(n_208),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_507),
.B(n_433),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_510),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_510),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_497),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_493),
.B(n_477),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_512),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_497),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_559),
.B(n_221),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_557),
.B(n_482),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_512),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_496),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_496),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_496),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_508),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_530),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_548),
.Y(n_621)
);

NOR2x1_ASAP7_75t_L g622 ( 
.A(n_501),
.B(n_539),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_503),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_497),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

AOI21x1_ASAP7_75t_L g626 ( 
.A1(n_524),
.A2(n_233),
.B(n_224),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_516),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_568),
.B(n_491),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_501),
.B(n_488),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_568),
.B(n_238),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_515),
.B(n_528),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_547),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_548),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_505),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_497),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_503),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_535),
.B(n_463),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_503),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_569),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_524),
.A2(n_254),
.B(n_235),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_516),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_504),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_535),
.B(n_468),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_497),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_559),
.B(n_477),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_516),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_544),
.B(n_480),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_562),
.B(n_541),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_554),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_504),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_499),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_562),
.B(n_541),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_554),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_529),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_499),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_554),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

AND3x2_ASAP7_75t_L g660 ( 
.A(n_511),
.B(n_462),
.C(n_460),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_499),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_530),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_554),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_554),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_499),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_554),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_534),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_534),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_567),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_567),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_499),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_548),
.B(n_438),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_519),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_559),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_538),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_562),
.B(n_541),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_544),
.B(n_486),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_504),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_511),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_561),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_547),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_499),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_517),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_533),
.Y(n_688)
);

NOR2x1p5_ASAP7_75t_L g689 ( 
.A(n_566),
.B(n_372),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_563),
.B(n_405),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_567),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_560),
.B(n_419),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_517),
.Y(n_693)
);

INVxp33_ASAP7_75t_L g694 ( 
.A(n_533),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_560),
.B(n_568),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_567),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_546),
.B(n_448),
.C(n_243),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_517),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_499),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_568),
.B(n_279),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_568),
.B(n_280),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_568),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_506),
.A2(n_365),
.B1(n_349),
.B2(n_230),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_564),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_518),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_546),
.B(n_248),
.C(n_242),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_543),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_L g709 ( 
.A(n_513),
.B(n_230),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_518),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_518),
.Y(n_711)
);

AO21x2_ASAP7_75t_L g712 ( 
.A1(n_513),
.A2(n_274),
.B(n_265),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_566),
.A2(n_299),
.B1(n_312),
.B2(n_314),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_565),
.B(n_261),
.C(n_252),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_563),
.B(n_199),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_563),
.Y(n_716)
);

AND3x2_ASAP7_75t_L g717 ( 
.A(n_543),
.B(n_293),
.C(n_283),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_518),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_545),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_522),
.Y(n_720)
);

AND2x6_ASAP7_75t_L g721 ( 
.A(n_563),
.B(n_230),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_545),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_523),
.B(n_297),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_712),
.A2(n_649),
.B1(n_677),
.B2(n_654),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_620),
.B(n_349),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_597),
.B(n_526),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_597),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_575),
.B(n_523),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_620),
.B(n_349),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_662),
.B(n_349),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_703),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_573),
.A2(n_526),
.B1(n_527),
.B2(n_549),
.C(n_532),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_662),
.B(n_365),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_703),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_649),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_SL g736 ( 
.A(n_598),
.B(n_373),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_581),
.B(n_529),
.C(n_570),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_654),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_667),
.B(n_365),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_716),
.B(n_523),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_632),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_582),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_595),
.B(n_586),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_681),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_638),
.A2(n_357),
.B1(n_322),
.B2(n_321),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_716),
.B(n_523),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_582),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_667),
.B(n_365),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_677),
.B(n_545),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_668),
.B(n_337),
.Y(n_750)
);

NAND2x1_ASAP7_75t_L g751 ( 
.A(n_720),
.B(n_524),
.Y(n_751)
);

INVxp33_ASAP7_75t_L g752 ( 
.A(n_692),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_690),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_573),
.A2(n_588),
.B(n_644),
.C(n_690),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_632),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_576),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_668),
.B(n_337),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_576),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_588),
.A2(n_527),
.B(n_532),
.C(n_556),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_622),
.B(n_337),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_574),
.B(n_202),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_585),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_583),
.B(n_202),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_622),
.B(n_337),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_719),
.B(n_522),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_689),
.A2(n_316),
.B1(n_298),
.B2(n_300),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_585),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_598),
.B(n_537),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_675),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_577),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_577),
.B(n_545),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_673),
.B(n_537),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_719),
.B(n_522),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_SL g774 ( 
.A(n_689),
.B(n_374),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_605),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_681),
.B(n_688),
.Y(n_776)
);

O2A1O1Ixp5_ASAP7_75t_L g777 ( 
.A1(n_626),
.A2(n_320),
.B(n_379),
.C(n_376),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_587),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_578),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_587),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_589),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_712),
.A2(n_524),
.B1(n_342),
.B2(n_330),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_675),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_688),
.B(n_549),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_722),
.B(n_522),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_578),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_694),
.B(n_551),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_593),
.B(n_205),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_580),
.B(n_572),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_602),
.B(n_205),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_589),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_580),
.B(n_572),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_683),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_584),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_674),
.B(n_536),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_584),
.B(n_591),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_683),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_611),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_602),
.B(n_551),
.Y(n_799)
);

OAI221xp5_ASAP7_75t_L g800 ( 
.A1(n_697),
.A2(n_556),
.B1(n_553),
.B2(n_555),
.C(n_570),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_707),
.A2(n_307),
.B1(n_311),
.B2(n_313),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_591),
.B(n_572),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_592),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_605),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_592),
.B(n_572),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_722),
.B(n_522),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_594),
.B(n_522),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_648),
.B(n_553),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_594),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_706),
.B(n_522),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_674),
.B(n_479),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_712),
.B(n_306),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_704),
.A2(n_309),
.B1(n_308),
.B2(n_346),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_629),
.B(n_555),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_678),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_L g816 ( 
.A(n_656),
.B(n_714),
.C(n_713),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_706),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_635),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_723),
.B(n_360),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_710),
.B(n_520),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_674),
.B(n_211),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_721),
.B(n_630),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_590),
.B(n_525),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_603),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_715),
.B(n_276),
.C(n_268),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_682),
.B(n_479),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_710),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_711),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_590),
.B(n_525),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_695),
.B(n_211),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_709),
.A2(n_315),
.B1(n_326),
.B2(n_332),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_590),
.B(n_525),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_579),
.B(n_483),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_608),
.B(n_613),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_718),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_603),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_604),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_718),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_720),
.B(n_605),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_579),
.B(n_483),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_717),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_720),
.B(n_520),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_605),
.B(n_520),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_721),
.A2(n_386),
.B1(n_381),
.B2(n_374),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_608),
.B(n_542),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_604),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_605),
.B(n_520),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_708),
.B(n_484),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_596),
.B(n_212),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_607),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_579),
.B(n_484),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_613),
.B(n_542),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_596),
.B(n_212),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_613),
.B(n_550),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_607),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_660),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_609),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_600),
.B(n_487),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_609),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_615),
.A2(n_459),
.B(n_440),
.C(n_441),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_624),
.B(n_550),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_624),
.B(n_550),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_615),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_624),
.B(n_645),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_616),
.B(n_618),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_665),
.B(n_334),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_606),
.B(n_441),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_616),
.B(n_618),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_665),
.B(n_335),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_650),
.B(n_487),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_623),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_674),
.B(n_490),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_623),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_665),
.B(n_341),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_645),
.B(n_558),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_606),
.B(n_451),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_619),
.B(n_490),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_721),
.A2(n_386),
.B1(n_384),
.B2(n_377),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_665),
.B(n_343),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_612),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_645),
.B(n_558),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_633),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_600),
.B(n_348),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_708),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_665),
.B(n_352),
.Y(n_885)
);

INVx8_ASAP7_75t_L g886 ( 
.A(n_674),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_721),
.B(n_353),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_621),
.B(n_215),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_721),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_652),
.B(n_558),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_724),
.B(n_619),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_SL g892 ( 
.A(n_737),
.B(n_754),
.C(n_816),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_776),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_808),
.B(n_619),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_744),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_787),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_751),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_770),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_818),
.Y(n_900)
);

NOR2x1p5_ASAP7_75t_L g901 ( 
.A(n_848),
.B(n_621),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_809),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_743),
.A2(n_631),
.B1(n_628),
.B2(n_610),
.Y(n_903)
);

INVxp67_ASAP7_75t_SL g904 ( 
.A(n_741),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_R g905 ( 
.A(n_736),
.B(n_676),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_826),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_743),
.A2(n_721),
.B1(n_637),
.B2(n_686),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_814),
.B(n_637),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_809),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_772),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_795),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_741),
.B(n_640),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_752),
.B(n_672),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_799),
.B(n_631),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_817),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_857),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_724),
.B(n_652),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_815),
.B(n_599),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_735),
.B(n_652),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_795),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_728),
.B(n_639),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_738),
.B(n_639),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_857),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_784),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_884),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_880),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_753),
.A2(n_610),
.B1(n_601),
.B2(n_700),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_867),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_804),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_863),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_754),
.A2(n_643),
.B(n_659),
.C(n_679),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_833),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_768),
.B(n_749),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_756),
.B(n_758),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_779),
.B(n_786),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_795),
.B(n_606),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_794),
.B(n_643),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_L g938 ( 
.A(n_788),
.B(n_634),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_803),
.B(n_651),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_871),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_SL g941 ( 
.A(n_774),
.B(n_656),
.C(n_381),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_873),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_726),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_882),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_727),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_726),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_SL g947 ( 
.A1(n_732),
.A2(n_705),
.B1(n_610),
.B2(n_601),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_880),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_769),
.B(n_657),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_790),
.B(n_599),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_840),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_759),
.A2(n_471),
.B(n_455),
.C(n_453),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_804),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_796),
.B(n_651),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_769),
.B(n_657),
.Y(n_955)
);

NOR2x2_ASAP7_75t_L g956 ( 
.A(n_811),
.B(n_599),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_827),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_755),
.B(n_659),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_755),
.B(n_679),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_828),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_775),
.A2(n_661),
.B(n_636),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_761),
.A2(n_721),
.B1(n_686),
.B2(n_693),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_793),
.B(n_693),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_769),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_793),
.B(n_698),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_769),
.B(n_657),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_761),
.A2(n_698),
.B1(n_627),
.B2(n_617),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_825),
.B(n_384),
.C(n_377),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_804),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_804),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_727),
.Y(n_971)
);

NOR2x1p5_ASAP7_75t_L g972 ( 
.A(n_867),
.B(n_634),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_783),
.B(n_606),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_797),
.B(n_889),
.Y(n_974)
);

NOR2xp67_ASAP7_75t_L g975 ( 
.A(n_788),
.B(n_705),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_759),
.B(n_685),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_763),
.A2(n_627),
.B1(n_612),
.B2(n_614),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_763),
.B(n_599),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_783),
.B(n_646),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_849),
.B(n_685),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_835),
.Y(n_981)
);

AND2x2_ASAP7_75t_SL g982 ( 
.A(n_844),
.B(n_701),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_851),
.B(n_601),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_849),
.B(n_685),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_856),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_782),
.A2(n_601),
.B1(n_610),
.B2(n_646),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_853),
.B(n_699),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_797),
.B(n_699),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_797),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_876),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_797),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_877),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_750),
.A2(n_610),
.B1(n_601),
.B2(n_646),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_782),
.A2(n_646),
.B1(n_699),
.B2(n_641),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_745),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_853),
.B(n_636),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_838),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_813),
.A2(n_626),
.B1(n_641),
.B2(n_636),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_889),
.B(n_640),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_865),
.B(n_661),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_742),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_747),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_886),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_762),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_750),
.A2(n_661),
.B1(n_671),
.B2(n_691),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_876),
.B(n_359),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_771),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_858),
.B(n_359),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_841),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_767),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_789),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_812),
.A2(n_729),
.B(n_730),
.C(n_725),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_811),
.B(n_650),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_886),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_865),
.B(n_671),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_778),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_844),
.A2(n_625),
.B1(n_642),
.B2(n_647),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_SL g1019 ( 
.A1(n_878),
.A2(n_389),
.B1(n_328),
.B2(n_329),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_889),
.B(n_640),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_811),
.B(n_653),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_888),
.B(n_281),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_872),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_800),
.B(n_284),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_798),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_868),
.B(n_642),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_R g1027 ( 
.A(n_821),
.B(n_215),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_889),
.B(n_640),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_819),
.B(n_289),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_872),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_792),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_766),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_872),
.B(n_653),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_868),
.B(n_647),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_757),
.A2(n_874),
.B1(n_879),
.B2(n_869),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_802),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_830),
.B(n_655),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_740),
.B(n_655),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_870),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_780),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_870),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_883),
.B(n_459),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_805),
.B(n_658),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_807),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_870),
.Y(n_1045)
);

AND2x4_ASAP7_75t_SL g1046 ( 
.A(n_878),
.B(n_466),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_801),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_725),
.B(n_729),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_831),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_843),
.B(n_640),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_733),
.B(n_467),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_731),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_733),
.B(n_658),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_870),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_781),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_760),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_791),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_739),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_866),
.A2(n_670),
.B1(n_696),
.B2(n_687),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_824),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_836),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_870),
.Y(n_1062)
);

AND2x4_ASAP7_75t_SL g1063 ( 
.A(n_734),
.B(n_467),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_777),
.A2(n_666),
.B(n_687),
.Y(n_1064)
);

AOI22x1_ASAP7_75t_L g1065 ( 
.A1(n_837),
.A2(n_859),
.B1(n_846),
.B2(n_850),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_866),
.A2(n_879),
.B1(n_874),
.B2(n_885),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_855),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_839),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_739),
.B(n_663),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_746),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_810),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_760),
.B(n_640),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_810),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_SL g1074 ( 
.A(n_860),
.B(n_344),
.C(n_333),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_823),
.Y(n_1075)
);

AO21x2_ASAP7_75t_L g1076 ( 
.A1(n_892),
.A2(n_764),
.B(n_885),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_917),
.A2(n_764),
.B(n_820),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_SL g1078 ( 
.A(n_986),
.B(n_217),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_945),
.B(n_973),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_899),
.Y(n_1080)
);

OR2x6_ASAP7_75t_SL g1081 ( 
.A(n_995),
.B(n_292),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_895),
.B(n_748),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_899),
.Y(n_1083)
);

AOI33xp33_ASAP7_75t_L g1084 ( 
.A1(n_906),
.A2(n_476),
.A3(n_472),
.B1(n_471),
.B2(n_470),
.B3(n_469),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_902),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1007),
.B(n_829),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1024),
.A2(n_822),
.B(n_869),
.C(n_813),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1046),
.A2(n_847),
.B1(n_843),
.B2(n_860),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_932),
.B(n_218),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1000),
.A2(n_1016),
.B(n_996),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_924),
.B(n_469),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_902),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_951),
.B(n_219),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_897),
.B(n_910),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_908),
.B(n_832),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_961),
.A2(n_847),
.B(n_839),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_909),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1029),
.B(n_934),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_1014),
.B(n_842),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1012),
.A2(n_834),
.B(n_864),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_893),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_935),
.B(n_845),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_917),
.A2(n_842),
.B(n_820),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1011),
.B(n_852),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_915),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_992),
.B(n_914),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_930),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_940),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1037),
.A2(n_887),
.B(n_862),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_942),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1024),
.A2(n_890),
.B(n_881),
.C(n_875),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_964),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_916),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_950),
.B(n_219),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1031),
.B(n_854),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_891),
.A2(n_861),
.B(n_806),
.C(n_785),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1036),
.B(n_765),
.Y(n_1117)
);

OAI22xp33_ASAP7_75t_SL g1118 ( 
.A1(n_891),
.A2(n_978),
.B1(n_1022),
.B2(n_950),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_916),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_964),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_933),
.A2(n_806),
.B(n_785),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_R g1122 ( 
.A(n_1047),
.B(n_222),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1070),
.B(n_765),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_933),
.A2(n_702),
.B(n_773),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_923),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_978),
.A2(n_356),
.B1(n_773),
.B2(n_388),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1046),
.A2(n_222),
.B1(n_358),
.B2(n_368),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1056),
.A2(n_982),
.B1(n_907),
.B2(n_1032),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_944),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_964),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_983),
.A2(n_663),
.B(n_684),
.C(n_680),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_896),
.B(n_470),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_964),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_900),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_980),
.A2(n_684),
.B(n_680),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_984),
.A2(n_702),
.B(n_670),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_926),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1008),
.B(n_476),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_943),
.Y(n_1139)
);

BUFx12f_ASAP7_75t_L g1140 ( 
.A(n_985),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_945),
.B(n_407),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1044),
.B(n_664),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_983),
.B(n_327),
.C(n_347),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1022),
.A2(n_669),
.B(n_666),
.C(n_664),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_969),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_952),
.A2(n_1025),
.B(n_913),
.C(n_918),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_987),
.A2(n_669),
.B(n_378),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_952),
.A2(n_412),
.B(n_409),
.C(n_408),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_928),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1075),
.B(n_571),
.Y(n_1150)
);

CKINVDCx16_ASAP7_75t_R g1151 ( 
.A(n_905),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_913),
.A2(n_412),
.B(n_409),
.C(n_408),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_982),
.A2(n_350),
.B1(n_351),
.B2(n_383),
.Y(n_1153)
);

AO32x1_ASAP7_75t_L g1154 ( 
.A1(n_994),
.A2(n_407),
.A3(n_571),
.B1(n_9),
.B2(n_11),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_894),
.B(n_368),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_918),
.A2(n_571),
.B(n_8),
.C(n_11),
.Y(n_1156)
);

AOI22x1_ASAP7_75t_L g1157 ( 
.A1(n_1042),
.A2(n_358),
.B1(n_383),
.B2(n_382),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_926),
.Y(n_1158)
);

NOR2xp67_ASAP7_75t_L g1159 ( 
.A(n_938),
.B(n_223),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_925),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_975),
.B(n_223),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_969),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1026),
.A2(n_1034),
.B(n_921),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1075),
.B(n_382),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_948),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_954),
.B(n_378),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_976),
.A2(n_134),
.B(n_64),
.C(n_74),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1032),
.A2(n_371),
.B1(n_231),
.B2(n_228),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_969),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_973),
.B(n_141),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_998),
.A2(n_227),
.B(n_371),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_919),
.A2(n_922),
.B(n_1058),
.C(n_946),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1049),
.A2(n_231),
.B1(n_228),
.B2(n_227),
.Y(n_1173)
);

AOI222xp33_ASAP7_75t_L g1174 ( 
.A1(n_1019),
.A2(n_2),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_18),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_981),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_920),
.B(n_1003),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_973),
.B(n_194),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_974),
.A2(n_123),
.B(n_188),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_971),
.B(n_947),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_919),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_903),
.A2(n_569),
.B1(n_167),
.B2(n_163),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_997),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_SL g1183 ( 
.A(n_1027),
.B(n_19),
.C(n_21),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_R g1184 ( 
.A(n_1003),
.B(n_145),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_SL g1185 ( 
.A1(n_936),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_990),
.Y(n_1186)
);

AO21x1_ASAP7_75t_L g1187 ( 
.A1(n_1066),
.A2(n_22),
.B(n_24),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_968),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1072),
.A2(n_113),
.B(n_136),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1051),
.B(n_26),
.Y(n_1190)
);

NOR2x1_ASAP7_75t_L g1191 ( 
.A(n_1015),
.B(n_130),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_931),
.A2(n_32),
.B(n_33),
.C(n_36),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_1006),
.B(n_32),
.C(n_37),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_997),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1072),
.A2(n_114),
.B(n_109),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_SL g1196 ( 
.A(n_1027),
.B(n_38),
.C(n_40),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_957),
.A2(n_45),
.B(n_47),
.C(n_50),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1048),
.A2(n_45),
.B(n_51),
.C(n_54),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1071),
.B(n_569),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_979),
.B(n_107),
.Y(n_1200)
);

XOR2xp5_ASAP7_75t_L g1201 ( 
.A(n_927),
.B(n_104),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_937),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1009),
.B(n_51),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_939),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1048),
.A2(n_54),
.B(n_61),
.C(n_63),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1015),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1030),
.B(n_61),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_962),
.A2(n_569),
.B1(n_993),
.B2(n_1035),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_904),
.B(n_1063),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_960),
.B(n_569),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1043),
.A2(n_569),
.B(n_949),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1073),
.B(n_1068),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1023),
.B(n_1068),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_905),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_989),
.B(n_991),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1018),
.A2(n_1068),
.B1(n_977),
.B2(n_967),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_955),
.A2(n_988),
.B(n_966),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_936),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_901),
.B(n_941),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_989),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_955),
.A2(n_898),
.B(n_965),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1001),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1023),
.B(n_1052),
.Y(n_1223)
);

OA22x2_ASAP7_75t_L g1224 ( 
.A1(n_936),
.A2(n_1013),
.B1(n_1021),
.B2(n_1033),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1001),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1098),
.A2(n_1021),
.B(n_1013),
.Y(n_1226)
);

NAND3x1_ASAP7_75t_L g1227 ( 
.A(n_1219),
.B(n_911),
.C(n_956),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1202),
.B(n_1038),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_1087),
.A2(n_959),
.B(n_958),
.C(n_963),
.Y(n_1229)
);

AO32x2_ASAP7_75t_L g1230 ( 
.A1(n_1128),
.A2(n_970),
.A3(n_1074),
.B1(n_956),
.B2(n_1014),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1111),
.A2(n_1064),
.B(n_1059),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1204),
.B(n_1055),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1105),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1187),
.A2(n_1041),
.A3(n_1069),
.B(n_1053),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1160),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1132),
.Y(n_1236)
);

INVx3_ASAP7_75t_R g1237 ( 
.A(n_1214),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1096),
.A2(n_1065),
.B(n_898),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1163),
.A2(n_970),
.B(n_898),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_L g1240 ( 
.A(n_1140),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1107),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1101),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1128),
.A2(n_1033),
.B1(n_1021),
.B2(n_1013),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1134),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1086),
.B(n_1067),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1086),
.B(n_1040),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1108),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1095),
.B(n_1040),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_1186),
.B(n_911),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1110),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1138),
.B(n_972),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1176),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1145),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1109),
.A2(n_1038),
.B(n_1050),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1174),
.B(n_1033),
.C(n_1054),
.Y(n_1255)
);

NOR3xp33_ASAP7_75t_L g1256 ( 
.A(n_1143),
.B(n_1060),
.C(n_1039),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1091),
.B(n_1017),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1103),
.A2(n_1038),
.B(n_1050),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1224),
.B(n_1045),
.Y(n_1259)
);

AOI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1135),
.A2(n_1004),
.B(n_1061),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1129),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1121),
.A2(n_1060),
.B(n_1055),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1102),
.A2(n_912),
.B(n_1005),
.Y(n_1263)
);

AO21x1_ASAP7_75t_L g1264 ( 
.A1(n_1118),
.A2(n_1017),
.B(n_1057),
.Y(n_1264)
);

AOI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1078),
.A2(n_1004),
.B(n_1010),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1173),
.B(n_1002),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1149),
.B(n_1164),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1077),
.A2(n_1057),
.B(n_1002),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_SL g1269 ( 
.A1(n_1212),
.A2(n_1192),
.B(n_1146),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1106),
.B(n_1010),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1145),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1162),
.Y(n_1272)
);

AO22x2_ASAP7_75t_L g1273 ( 
.A1(n_1208),
.A2(n_1062),
.B1(n_1039),
.B2(n_953),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1206),
.Y(n_1274)
);

AOI21xp33_ASAP7_75t_L g1275 ( 
.A1(n_1078),
.A2(n_1062),
.B(n_1054),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1216),
.A2(n_912),
.B(n_1020),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1131),
.A2(n_999),
.B(n_1028),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1206),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1194),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1136),
.A2(n_929),
.B(n_953),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1097),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1077),
.A2(n_1124),
.B(n_1211),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1139),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1104),
.B(n_929),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1116),
.A2(n_929),
.B(n_953),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1216),
.A2(n_1045),
.B(n_1054),
.Y(n_1287)
);

NOR2x1_ASAP7_75t_R g1288 ( 
.A(n_1206),
.B(n_1045),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1079),
.B(n_1045),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1174),
.A2(n_1054),
.B(n_1201),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1198),
.A2(n_1196),
.B(n_1183),
.C(n_1188),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1156),
.A2(n_1168),
.B(n_1173),
.C(n_1193),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1115),
.B(n_1082),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1112),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1224),
.B(n_1170),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1208),
.A2(n_1088),
.B(n_1147),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1162),
.A2(n_1088),
.B(n_1076),
.Y(n_1297)
);

AOI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_1212),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1172),
.A2(n_1181),
.B(n_1171),
.C(n_1114),
.Y(n_1299)
);

NOR2x1_ASAP7_75t_SL g1300 ( 
.A(n_1162),
.B(n_1076),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1170),
.A2(n_1177),
.B1(n_1200),
.B2(n_1179),
.Y(n_1301)
);

AO21x1_ASAP7_75t_L g1302 ( 
.A1(n_1180),
.A2(n_1144),
.B(n_1197),
.Y(n_1302)
);

O2A1O1Ixp5_ASAP7_75t_L g1303 ( 
.A1(n_1161),
.A2(n_1153),
.B(n_1166),
.C(n_1190),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1166),
.B(n_1123),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_1117),
.Y(n_1305)
);

OAI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1122),
.A2(n_1168),
.B(n_1127),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1083),
.B(n_1092),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1207),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1085),
.B(n_1080),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1199),
.A2(n_1178),
.B(n_1164),
.Y(n_1310)
);

INVx3_ASAP7_75t_SL g1311 ( 
.A(n_1151),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1220),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1222),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1094),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1225),
.B(n_1119),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1162),
.A2(n_1099),
.B(n_1209),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1113),
.A2(n_1165),
.B(n_1158),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1079),
.Y(n_1318)
);

O2A1O1Ixp5_ASAP7_75t_L g1319 ( 
.A1(n_1089),
.A2(n_1093),
.B(n_1155),
.C(n_1223),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1081),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1125),
.A2(n_1137),
.B(n_1199),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1189),
.A2(n_1195),
.B(n_1169),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1177),
.B(n_1213),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1203),
.A2(n_1152),
.B(n_1218),
.C(n_1167),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1215),
.A2(n_1154),
.B(n_1210),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1126),
.A2(n_1148),
.B(n_1159),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1084),
.B(n_1130),
.Y(n_1327)
);

OAI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1141),
.A2(n_1157),
.B(n_1184),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1141),
.A2(n_1191),
.B1(n_1130),
.B2(n_1133),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1112),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1120),
.A2(n_1014),
.B(n_1216),
.Y(n_1331)
);

NOR4xp25_ASAP7_75t_L g1332 ( 
.A(n_1120),
.B(n_892),
.C(n_1188),
.D(n_1183),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1128),
.A2(n_1098),
.B1(n_1046),
.B2(n_724),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1160),
.Y(n_1334)
);

AND2x6_ASAP7_75t_SL g1335 ( 
.A(n_1219),
.B(n_795),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1105),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1216),
.A2(n_1014),
.B(n_1208),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1098),
.B(n_895),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1105),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1118),
.A2(n_743),
.B(n_1098),
.C(n_892),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1176),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1087),
.A2(n_1111),
.B(n_892),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1128),
.A2(n_1098),
.B1(n_1046),
.B2(n_724),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1087),
.A2(n_1111),
.B(n_892),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1174),
.A2(n_648),
.B(n_581),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1175),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1135),
.A2(n_1100),
.B(n_1109),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1187),
.A2(n_1208),
.A3(n_1090),
.B(n_952),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1146),
.A2(n_743),
.B(n_978),
.C(n_950),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1098),
.B(n_895),
.Y(n_1350)
);

NAND2xp33_ASAP7_75t_R g1351 ( 
.A(n_1122),
.B(n_598),
.Y(n_1351)
);

O2A1O1Ixp5_ASAP7_75t_L g1352 ( 
.A1(n_1098),
.A2(n_978),
.B(n_950),
.C(n_788),
.Y(n_1352)
);

AO21x2_ASAP7_75t_L g1353 ( 
.A1(n_1090),
.A2(n_1131),
.B(n_1135),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1160),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1175),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1087),
.A2(n_1111),
.B(n_892),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1098),
.B(n_1202),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1128),
.A2(n_1098),
.B1(n_1046),
.B2(n_724),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1096),
.A2(n_1221),
.B(n_1217),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1105),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1096),
.A2(n_1221),
.B(n_1217),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1096),
.A2(n_1221),
.B(n_1217),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1098),
.B(n_895),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1345),
.A2(n_1349),
.B(n_1292),
.C(n_1306),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1340),
.A2(n_1344),
.B(n_1342),
.C(n_1356),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1273),
.Y(n_1366)
);

BUFx2_ASAP7_75t_SL g1367 ( 
.A(n_1235),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1257),
.B(n_1270),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1359),
.A2(n_1362),
.B(n_1361),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1272),
.Y(n_1370)
);

NAND2x1_ASAP7_75t_L g1371 ( 
.A(n_1331),
.B(n_1253),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1347),
.A2(n_1262),
.B(n_1283),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1322),
.A2(n_1297),
.B(n_1226),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1281),
.A2(n_1258),
.B(n_1286),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1272),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1311),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1354),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1352),
.A2(n_1303),
.B(n_1299),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1317),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1295),
.B(n_1289),
.Y(n_1380)
);

BUFx8_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1321),
.A2(n_1310),
.B(n_1231),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1338),
.A2(n_1363),
.B(n_1350),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_SL g1384 ( 
.A(n_1240),
.B(n_1252),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1342),
.A2(n_1356),
.B(n_1344),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1304),
.A2(n_1293),
.B(n_1310),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1304),
.A2(n_1293),
.B(n_1291),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1319),
.A2(n_1326),
.B(n_1357),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1233),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1295),
.B(n_1259),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1357),
.B(n_1236),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1278),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1296),
.A2(n_1268),
.B(n_1276),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1269),
.A2(n_1324),
.B(n_1264),
.Y(n_1394)
);

CKINVDCx16_ASAP7_75t_R g1395 ( 
.A(n_1351),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1280),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1302),
.A2(n_1300),
.A3(n_1325),
.B(n_1333),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_SL g1398 ( 
.A(n_1240),
.B(n_1341),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1301),
.A2(n_1290),
.B1(n_1323),
.B2(n_1236),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1272),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1267),
.B(n_1323),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1263),
.A2(n_1337),
.B(n_1229),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1305),
.A2(n_1298),
.B(n_1287),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1320),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1244),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1237),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1272),
.B(n_1253),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1241),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1279),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1247),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1271),
.B(n_1329),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1335),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1334),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1346),
.Y(n_1414)
);

AOI21xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1251),
.A2(n_1308),
.B(n_1301),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1326),
.A2(n_1343),
.B(n_1333),
.Y(n_1416)
);

CKINVDCx6p67_ASAP7_75t_R g1417 ( 
.A(n_1312),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1268),
.A2(n_1287),
.B(n_1316),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1318),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1314),
.B(n_1232),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1343),
.A2(n_1358),
.B(n_1328),
.C(n_1332),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1232),
.B(n_1228),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1255),
.A2(n_1295),
.B1(n_1358),
.B2(n_1259),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1266),
.A2(n_1256),
.B1(n_1327),
.B2(n_1243),
.Y(n_1425)
);

NOR3xp33_ASAP7_75t_L g1426 ( 
.A(n_1243),
.B(n_1275),
.C(n_1327),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1250),
.Y(n_1427)
);

O2A1O1Ixp5_ASAP7_75t_L g1428 ( 
.A1(n_1275),
.A2(n_1265),
.B(n_1248),
.C(n_1285),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1289),
.B(n_1284),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1273),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1248),
.A2(n_1285),
.B(n_1246),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1271),
.B(n_1282),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1294),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1261),
.B(n_1360),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1307),
.A2(n_1309),
.B(n_1315),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1227),
.A2(n_1313),
.B(n_1355),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1336),
.A2(n_1339),
.B(n_1353),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1259),
.B(n_1274),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1353),
.A2(n_1348),
.B(n_1273),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1348),
.A2(n_1277),
.B(n_1249),
.Y(n_1440)
);

BUFx2_ASAP7_75t_R g1441 ( 
.A(n_1330),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1294),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1294),
.B(n_1348),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1288),
.B(n_1230),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1234),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1230),
.A2(n_1234),
.B(n_1277),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1234),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1233),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1233),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1295),
.B(n_1289),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1272),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1233),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1233),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1238),
.A2(n_1260),
.B(n_1239),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1295),
.B(n_1289),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1345),
.A2(n_1349),
.B(n_1292),
.C(n_1306),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1295),
.B(n_1259),
.Y(n_1457)
);

AO32x2_ASAP7_75t_L g1458 ( 
.A1(n_1333),
.A2(n_1343),
.A3(n_1358),
.B1(n_1185),
.B2(n_1128),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1352),
.A2(n_1349),
.B(n_1345),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1349),
.A2(n_1205),
.B(n_1198),
.C(n_1299),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1345),
.A2(n_1340),
.B(n_1356),
.C(n_1344),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1252),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1311),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1317),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1279),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1272),
.B(n_1162),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1317),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1257),
.B(n_895),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1233),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1233),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1317),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1238),
.A2(n_1239),
.B(n_1254),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1236),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1231),
.A2(n_1296),
.B(n_1342),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1317),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1233),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1317),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1317),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1352),
.A2(n_1349),
.B(n_1345),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1272),
.B(n_1162),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1317),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1257),
.B(n_895),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1345),
.A2(n_1349),
.B(n_1292),
.C(n_1306),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1238),
.A2(n_1239),
.B(n_1254),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1272),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1233),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1233),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1345),
.A2(n_1340),
.B(n_1356),
.C(n_1344),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1233),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1235),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1233),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1306),
.A2(n_1174),
.B1(n_892),
.B2(n_737),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1272),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_SL g1494 ( 
.A1(n_1349),
.A2(n_1205),
.B(n_1198),
.C(n_1299),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1345),
.A2(n_598),
.B1(n_1301),
.B2(n_1357),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1238),
.A2(n_1260),
.B(n_1239),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1317),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1306),
.A2(n_1174),
.B1(n_892),
.B2(n_737),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1233),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1233),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1357),
.B(n_1304),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1231),
.A2(n_1296),
.B(n_1342),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1345),
.A2(n_1340),
.B(n_1356),
.C(n_1344),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1257),
.B(n_895),
.Y(n_1504)
);

INVxp33_ASAP7_75t_L g1505 ( 
.A(n_1468),
.Y(n_1505)
);

NOR2xp67_ASAP7_75t_L g1506 ( 
.A(n_1391),
.B(n_1462),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1380),
.B(n_1450),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1365),
.A2(n_1402),
.B(n_1460),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1365),
.A2(n_1494),
.B(n_1460),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1380),
.B(n_1450),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1409),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1368),
.B(n_1482),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1492),
.A2(n_1498),
.B1(n_1503),
.B2(n_1461),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1504),
.B(n_1429),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1364),
.A2(n_1456),
.B(n_1483),
.C(n_1461),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1401),
.B(n_1473),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1400),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1380),
.B(n_1450),
.Y(n_1518)
);

NOR2xp67_ASAP7_75t_L g1519 ( 
.A(n_1462),
.B(n_1413),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1459),
.B(n_1479),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1455),
.B(n_1399),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1503),
.A2(n_1488),
.B(n_1421),
.C(n_1498),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1488),
.A2(n_1480),
.B(n_1466),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1501),
.B(n_1387),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1492),
.A2(n_1395),
.B1(n_1495),
.B2(n_1425),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1420),
.B(n_1422),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1381),
.Y(n_1527)
);

AOI21x1_ASAP7_75t_SL g1528 ( 
.A1(n_1443),
.A2(n_1430),
.B(n_1366),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1388),
.A2(n_1415),
.B(n_1416),
.C(n_1383),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1466),
.A2(n_1480),
.B(n_1385),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1446),
.A2(n_1454),
.B(n_1496),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1437),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1390),
.B(n_1457),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1425),
.A2(n_1390),
.B1(n_1457),
.B2(n_1406),
.Y(n_1534)
);

O2A1O1Ixp5_ASAP7_75t_L g1535 ( 
.A1(n_1424),
.A2(n_1445),
.B(n_1386),
.C(n_1436),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1437),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1390),
.B(n_1457),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1406),
.A2(n_1417),
.B1(n_1419),
.B2(n_1412),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1392),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_R g1540 ( 
.A(n_1384),
.B(n_1398),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1454),
.A2(n_1496),
.B(n_1439),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1400),
.A2(n_1485),
.B(n_1451),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1377),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_SL g1544 ( 
.A1(n_1443),
.A2(n_1366),
.B(n_1430),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1394),
.A2(n_1426),
.B(n_1502),
.C(n_1474),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1426),
.A2(n_1434),
.B1(n_1428),
.B2(n_1412),
.C(n_1500),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1438),
.B(n_1409),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1423),
.B(n_1434),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1419),
.A2(n_1441),
.B1(n_1411),
.B2(n_1444),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1396),
.B(n_1389),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1414),
.B(n_1408),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1393),
.A2(n_1458),
.B(n_1371),
.C(n_1418),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1410),
.B(n_1427),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1411),
.A2(n_1444),
.B1(n_1438),
.B2(n_1490),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1448),
.B(n_1449),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1376),
.Y(n_1557)
);

O2A1O1Ixp5_ASAP7_75t_L g1558 ( 
.A1(n_1379),
.A2(n_1478),
.B(n_1497),
.C(n_1464),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1469),
.B(n_1499),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1405),
.A2(n_1367),
.B1(n_1432),
.B2(n_1463),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1447),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1465),
.B(n_1487),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1432),
.A2(n_1463),
.B1(n_1376),
.B2(n_1470),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1476),
.A2(n_1486),
.B1(n_1489),
.B2(n_1491),
.Y(n_1564)
);

O2A1O1Ixp5_ASAP7_75t_L g1565 ( 
.A1(n_1379),
.A2(n_1497),
.B(n_1464),
.C(n_1467),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1403),
.A2(n_1382),
.B(n_1373),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1404),
.A2(n_1407),
.B1(n_1485),
.B2(n_1400),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1458),
.B(n_1442),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1404),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1431),
.B(n_1435),
.Y(n_1570)
);

AOI21x1_ASAP7_75t_SL g1571 ( 
.A1(n_1440),
.A2(n_1397),
.B(n_1447),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1381),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1407),
.A2(n_1485),
.B1(n_1400),
.B2(n_1493),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1381),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1431),
.B(n_1397),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1431),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1372),
.A2(n_1484),
.B(n_1472),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1433),
.B(n_1397),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1433),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1433),
.Y(n_1580)
);

O2A1O1Ixp5_ASAP7_75t_L g1581 ( 
.A1(n_1471),
.A2(n_1475),
.B(n_1481),
.C(n_1477),
.Y(n_1581)
);

O2A1O1Ixp5_ASAP7_75t_L g1582 ( 
.A1(n_1478),
.A2(n_1451),
.B(n_1370),
.C(n_1375),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1374),
.A2(n_1369),
.B(n_1485),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1374),
.A2(n_1345),
.B1(n_1498),
.B2(n_1492),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1401),
.B(n_1391),
.Y(n_1585)
);

O2A1O1Ixp5_ASAP7_75t_L g1586 ( 
.A1(n_1378),
.A2(n_1342),
.B(n_1356),
.C(n_1344),
.Y(n_1586)
);

O2A1O1Ixp5_ASAP7_75t_L g1587 ( 
.A1(n_1378),
.A2(n_1342),
.B(n_1356),
.C(n_1344),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1365),
.A2(n_1288),
.B(n_1349),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1368),
.B(n_1468),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1462),
.Y(n_1590)
);

AND2x2_ASAP7_75t_SL g1591 ( 
.A(n_1385),
.B(n_1078),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1501),
.B(n_1387),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1364),
.A2(n_1345),
.B(n_1483),
.C(n_1456),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1437),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1368),
.B(n_1468),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1401),
.B(n_1391),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1492),
.A2(n_1345),
.B1(n_1498),
.B2(n_1290),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1501),
.B(n_1387),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1368),
.B(n_1468),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1409),
.Y(n_1600)
);

BUFx8_ASAP7_75t_SL g1601 ( 
.A(n_1376),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1461),
.A2(n_1345),
.B(n_1292),
.C(n_1349),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1492),
.A2(n_1345),
.B1(n_1498),
.B2(n_1290),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1501),
.B(n_1387),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1492),
.A2(n_1345),
.B1(n_1498),
.B2(n_1290),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1461),
.A2(n_1345),
.B(n_1292),
.C(n_1349),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1437),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1368),
.B(n_1468),
.Y(n_1608)
);

O2A1O1Ixp5_ASAP7_75t_L g1609 ( 
.A1(n_1378),
.A2(n_1342),
.B(n_1356),
.C(n_1344),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1492),
.A2(n_1345),
.B1(n_1498),
.B2(n_1290),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1409),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1492),
.A2(n_1345),
.B1(n_1498),
.B2(n_1290),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1378),
.A2(n_1446),
.B(n_1454),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1512),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1561),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1576),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1533),
.B(n_1537),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1593),
.A2(n_1515),
.B(n_1602),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1555),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1533),
.B(n_1537),
.Y(n_1620)
);

AOI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1508),
.A2(n_1509),
.B(n_1513),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1552),
.A2(n_1535),
.B(n_1586),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1601),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1571),
.A2(n_1565),
.B(n_1558),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1507),
.B(n_1510),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1591),
.B(n_1568),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1575),
.B(n_1570),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1507),
.B(n_1510),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1520),
.B(n_1561),
.Y(n_1630)
);

AO21x2_ASAP7_75t_L g1631 ( 
.A1(n_1532),
.A2(n_1607),
.B(n_1536),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1511),
.Y(n_1632)
);

OR2x2_ASAP7_75t_SL g1633 ( 
.A(n_1524),
.B(n_1592),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1518),
.B(n_1539),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1564),
.Y(n_1635)
);

AO21x2_ASAP7_75t_L g1636 ( 
.A1(n_1532),
.A2(n_1594),
.B(n_1607),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1571),
.A2(n_1565),
.B(n_1581),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1530),
.B(n_1523),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1550),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1559),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1583),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1562),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1516),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1553),
.Y(n_1644)
);

AO21x2_ASAP7_75t_L g1645 ( 
.A1(n_1545),
.A2(n_1522),
.B(n_1584),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1515),
.B(n_1593),
.C(n_1522),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1562),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1556),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1551),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1586),
.A2(n_1587),
.B(n_1609),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1588),
.A2(n_1606),
.B(n_1529),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1583),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1583),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1505),
.Y(n_1654)
);

OR2x6_ASAP7_75t_L g1655 ( 
.A(n_1554),
.B(n_1542),
.Y(n_1655)
);

BUFx4f_ASAP7_75t_SL g1656 ( 
.A(n_1557),
.Y(n_1656)
);

AOI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1525),
.A2(n_1597),
.B(n_1612),
.Y(n_1657)
);

INVx6_ASAP7_75t_L g1658 ( 
.A(n_1579),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1585),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1613),
.B(n_1596),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1535),
.A2(n_1587),
.B(n_1609),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1566),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1582),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1582),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1598),
.A2(n_1604),
.B(n_1605),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1603),
.A2(n_1610),
.B(n_1534),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1505),
.B(n_1514),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1531),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1549),
.B(n_1567),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1541),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1631),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1654),
.B(n_1531),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1531),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1660),
.B(n_1628),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1668),
.B(n_1627),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1641),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1668),
.B(n_1541),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1616),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1641),
.B(n_1547),
.Y(n_1679)
);

OAI222xp33_ASAP7_75t_L g1680 ( 
.A1(n_1657),
.A2(n_1521),
.B1(n_1563),
.B2(n_1548),
.C1(n_1560),
.C2(n_1526),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1665),
.B(n_1546),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1624),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1631),
.Y(n_1683)
);

AO21x2_ASAP7_75t_L g1684 ( 
.A1(n_1650),
.A2(n_1528),
.B(n_1544),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1665),
.B(n_1577),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1616),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1660),
.B(n_1543),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1665),
.B(n_1506),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1670),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1628),
.B(n_1644),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1664),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1636),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1663),
.B(n_1595),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1653),
.B(n_1608),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_SL g1695 ( 
.A(n_1638),
.B(n_1573),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1599),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_SL g1697 ( 
.A(n_1618),
.B(n_1540),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1517),
.Y(n_1698)
);

AND2x4_ASAP7_75t_SL g1699 ( 
.A(n_1638),
.B(n_1517),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1662),
.B(n_1589),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1687),
.B(n_1659),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1681),
.A2(n_1646),
.B1(n_1666),
.B2(n_1697),
.C(n_1680),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1678),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1666),
.C(n_1664),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1697),
.A2(n_1651),
.B1(n_1645),
.B2(n_1669),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1681),
.A2(n_1651),
.B(n_1645),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1678),
.Y(n_1707)
);

OAI31xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1675),
.A2(n_1651),
.A3(n_1620),
.B(n_1617),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1688),
.A2(n_1614),
.B(n_1648),
.C(n_1619),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1687),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1698),
.B(n_1638),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1680),
.A2(n_1645),
.B1(n_1635),
.B2(n_1643),
.C(n_1640),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1689),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1688),
.A2(n_1669),
.B1(n_1655),
.B2(n_1638),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_SL g1716 ( 
.A1(n_1695),
.A2(n_1669),
.B1(n_1657),
.B2(n_1622),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1675),
.B(n_1625),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1688),
.A2(n_1644),
.B1(n_1667),
.B2(n_1649),
.C(n_1634),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1687),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1675),
.B(n_1615),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1698),
.B(n_1615),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1691),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1693),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1691),
.A2(n_1669),
.B1(n_1655),
.B2(n_1538),
.C(n_1642),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1691),
.B(n_1661),
.C(n_1622),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1698),
.Y(n_1726)
);

OAI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1693),
.A2(n_1655),
.B1(n_1621),
.B2(n_1622),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1690),
.A2(n_1667),
.B1(n_1649),
.B2(n_1634),
.C(n_1639),
.Y(n_1728)
);

AOI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1691),
.A2(n_1630),
.B(n_1655),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1699),
.A2(n_1621),
.B(n_1620),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1630),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1694),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_SL g1733 ( 
.A(n_1685),
.B(n_1623),
.C(n_1569),
.Y(n_1733)
);

AOI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1700),
.A2(n_1647),
.B1(n_1629),
.B2(n_1626),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1703),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1722),
.B(n_1700),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1703),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1726),
.B(n_1672),
.Y(n_1738)
);

NOR2x1p5_ASAP7_75t_L g1739 ( 
.A(n_1704),
.B(n_1574),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1707),
.Y(n_1740)
);

AO21x2_ASAP7_75t_L g1741 ( 
.A1(n_1706),
.A2(n_1692),
.B(n_1671),
.Y(n_1741)
);

NOR2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1708),
.B(n_1623),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1710),
.B(n_1700),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1707),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1725),
.A2(n_1637),
.B(n_1676),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1714),
.Y(n_1746)
);

BUFx12f_ASAP7_75t_L g1747 ( 
.A(n_1711),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1719),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1712),
.B(n_1632),
.Y(n_1749)
);

NAND3x1_ASAP7_75t_L g1750 ( 
.A(n_1702),
.B(n_1677),
.C(n_1695),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1732),
.B(n_1672),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1732),
.B(n_1672),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1723),
.Y(n_1753)
);

OA21x2_ASAP7_75t_L g1754 ( 
.A1(n_1730),
.A2(n_1683),
.B(n_1671),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1718),
.B(n_1690),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1727),
.A2(n_1540),
.B(n_1519),
.C(n_1682),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1731),
.B(n_1673),
.Y(n_1757)
);

AOI32xp33_ASAP7_75t_L g1758 ( 
.A1(n_1749),
.A2(n_1705),
.A3(n_1716),
.B1(n_1709),
.B2(n_1724),
.Y(n_1758)
);

INVxp67_ASAP7_75t_SL g1759 ( 
.A(n_1750),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1755),
.B(n_1728),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1735),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_L g1762 ( 
.A(n_1739),
.B(n_1719),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1735),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1747),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1748),
.Y(n_1765)
);

BUFx3_ASAP7_75t_L g1766 ( 
.A(n_1747),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1735),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1755),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1747),
.B(n_1656),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1742),
.B(n_1731),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1737),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1756),
.B(n_1733),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1748),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1739),
.B(n_1742),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_SL g1775 ( 
.A(n_1756),
.B(n_1715),
.C(n_1734),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1749),
.B(n_1694),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1742),
.B(n_1721),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1753),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1743),
.B(n_1674),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1757),
.B(n_1721),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1739),
.B(n_1694),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1751),
.B(n_1711),
.Y(n_1782)
);

INVxp67_ASAP7_75t_SL g1783 ( 
.A(n_1750),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1743),
.B(n_1694),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1736),
.B(n_1674),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1750),
.A2(n_1729),
.B(n_1701),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1757),
.B(n_1721),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1737),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1747),
.A2(n_1661),
.B1(n_1684),
.B2(n_1679),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1746),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1751),
.B(n_1695),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1736),
.B(n_1674),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1746),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1740),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1740),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1746),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1757),
.B(n_1720),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1751),
.B(n_1717),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1751),
.B(n_1717),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1752),
.B(n_1713),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1674),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1761),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1768),
.B(n_1590),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1765),
.B(n_1773),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1761),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1763),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1760),
.B(n_1696),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1778),
.B(n_1633),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1762),
.B(n_1738),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1763),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1764),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1802),
.B(n_1633),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1758),
.B(n_1696),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1767),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1767),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1791),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1771),
.Y(n_1818)
);

NAND2x1_ASAP7_75t_L g1819 ( 
.A(n_1777),
.B(n_1754),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1771),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1758),
.B(n_1696),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1770),
.B(n_1754),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1784),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1766),
.B(n_1696),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1774),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1802),
.B(n_1740),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1776),
.B(n_1744),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1764),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1759),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1770),
.B(n_1754),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1784),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1789),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1795),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1774),
.B(n_1754),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1795),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1777),
.B(n_1754),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1796),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1796),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1791),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1810),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1805),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1825),
.B(n_1772),
.Y(n_1843)
);

BUFx3_ASAP7_75t_L g1844 ( 
.A(n_1825),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1829),
.B(n_1783),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1804),
.B(n_1766),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1810),
.B(n_1764),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1804),
.Y(n_1848)
);

NAND2x1p5_ASAP7_75t_L g1849 ( 
.A(n_1835),
.B(n_1769),
.Y(n_1849)
);

OAI21x1_ASAP7_75t_L g1850 ( 
.A1(n_1819),
.A2(n_1750),
.B(n_1794),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1815),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1810),
.B(n_1782),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1813),
.B(n_1786),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1839),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1812),
.B(n_1782),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1803),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1813),
.B(n_1786),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1808),
.B(n_1793),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1812),
.B(n_1799),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1809),
.Y(n_1860)
);

AO21x1_ASAP7_75t_SL g1861 ( 
.A1(n_1809),
.A2(n_1781),
.B(n_1787),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1828),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1806),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1828),
.B(n_1782),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1807),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1826),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1835),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1843),
.A2(n_1814),
.B(n_1821),
.C(n_1819),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1866),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1866),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1849),
.B(n_1792),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1849),
.A2(n_1790),
.B1(n_1824),
.B2(n_1792),
.Y(n_1872)
);

INVx1_ASAP7_75t_SL g1873 ( 
.A(n_1855),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1860),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1852),
.B(n_1837),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1842),
.B(n_1799),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1852),
.B(n_1837),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1845),
.A2(n_1775),
.B1(n_1830),
.B2(n_1822),
.C(n_1834),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1844),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1866),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1850),
.A2(n_1754),
.B(n_1822),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1851),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1849),
.A2(n_1792),
.B1(n_1754),
.B2(n_1800),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1848),
.A2(n_1830),
.B(n_1572),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1862),
.B(n_1800),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1851),
.Y(n_1886)
);

OAI31xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1850),
.A2(n_1867),
.A3(n_1861),
.B(n_1847),
.Y(n_1887)
);

INVxp67_ASAP7_75t_L g1888 ( 
.A(n_1844),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1879),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1873),
.B(n_1844),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1870),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1874),
.B(n_1862),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1870),
.Y(n_1893)
);

NAND2xp33_ASAP7_75t_R g1894 ( 
.A(n_1887),
.B(n_1854),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1875),
.B(n_1847),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1869),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1888),
.B(n_1841),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1875),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1880),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1877),
.B(n_1855),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1889),
.A2(n_1878),
.B(n_1868),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1892),
.A2(n_1886),
.B1(n_1882),
.B2(n_1872),
.C(n_1854),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1890),
.A2(n_1871),
.B(n_1881),
.C(n_1883),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1898),
.A2(n_1876),
.B1(n_1871),
.B2(n_1885),
.C(n_1867),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1897),
.A2(n_1846),
.B(n_1884),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1891),
.B(n_1841),
.Y(n_1906)
);

OAI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1894),
.A2(n_1898),
.B1(n_1859),
.B2(n_1895),
.C(n_1841),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1900),
.B(n_1864),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1894),
.B(n_1861),
.C(n_1864),
.Y(n_1909)
);

OAI21xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1900),
.A2(n_1877),
.B(n_1857),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1896),
.B(n_1853),
.Y(n_1911)
);

NAND3xp33_ASAP7_75t_L g1912 ( 
.A(n_1899),
.B(n_1863),
.C(n_1856),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1906),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1909),
.A2(n_1908),
.B1(n_1901),
.B2(n_1910),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1911),
.Y(n_1915)
);

NOR2x1_ASAP7_75t_L g1916 ( 
.A(n_1907),
.B(n_1893),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1912),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1903),
.A2(n_1865),
.B1(n_1863),
.B2(n_1856),
.C(n_1840),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1913),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1914),
.B(n_1904),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1915),
.B(n_1905),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1916),
.B(n_1902),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1917),
.B(n_1865),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1918),
.B(n_1853),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1914),
.B(n_1857),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1921),
.B(n_1858),
.Y(n_1926)
);

AO22x1_ASAP7_75t_L g1927 ( 
.A1(n_1922),
.A2(n_1817),
.B1(n_1840),
.B2(n_1838),
.Y(n_1927)
);

AOI332xp33_ASAP7_75t_L g1928 ( 
.A1(n_1919),
.A2(n_1817),
.A3(n_1836),
.B1(n_1833),
.B2(n_1832),
.B3(n_1831),
.C1(n_1818),
.C2(n_1816),
.Y(n_1928)
);

AOI222xp33_ASAP7_75t_L g1929 ( 
.A1(n_1920),
.A2(n_1823),
.B1(n_1820),
.B2(n_1811),
.C1(n_1794),
.C2(n_1797),
.Y(n_1929)
);

AND3x1_ASAP7_75t_L g1930 ( 
.A(n_1923),
.B(n_1527),
.C(n_1797),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1925),
.B(n_1924),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_L g1932 ( 
.A1(n_1931),
.A2(n_1858),
.B1(n_1827),
.B2(n_1741),
.C(n_1826),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1930),
.B(n_1926),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1929),
.A2(n_1658),
.B1(n_1827),
.B2(n_1741),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1927),
.B(n_1600),
.Y(n_1935)
);

AOI32xp33_ASAP7_75t_L g1936 ( 
.A1(n_1935),
.A2(n_1933),
.A3(n_1932),
.B1(n_1928),
.B2(n_1934),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1936),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1937),
.B(n_1801),
.Y(n_1938)
);

XNOR2x1_ASAP7_75t_L g1939 ( 
.A(n_1937),
.B(n_1580),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1938),
.A2(n_1801),
.B1(n_1658),
.B2(n_1741),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1939),
.Y(n_1941)
);

OAI22x1_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1801),
.B1(n_1746),
.B2(n_1798),
.Y(n_1942)
);

BUFx2_ASAP7_75t_L g1943 ( 
.A(n_1940),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1943),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1944),
.A2(n_1942),
.B(n_1611),
.Y(n_1945)
);

AOI31xp67_ASAP7_75t_SL g1946 ( 
.A1(n_1945),
.A2(n_1658),
.A3(n_1785),
.B(n_1744),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1946),
.A2(n_1658),
.B1(n_1788),
.B2(n_1780),
.Y(n_1947)
);

OAI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1947),
.A2(n_1793),
.B1(n_1779),
.B2(n_1611),
.Y(n_1948)
);

AOI211xp5_ASAP7_75t_L g1949 ( 
.A1(n_1948),
.A2(n_1600),
.B(n_1745),
.C(n_1632),
.Y(n_1949)
);


endmodule