module fake_jpeg_10188_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_32),
.Y(n_60)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_18),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_34),
.B1(n_29),
.B2(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_18),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_21),
.B1(n_24),
.B2(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_60),
.Y(n_95)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_19),
.B1(n_17),
.B2(n_26),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_29),
.B1(n_34),
.B2(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_81),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_92),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_90),
.B1(n_48),
.B2(n_17),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_38),
.B1(n_40),
.B2(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_88),
.B1(n_64),
.B2(n_51),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AOI22x1_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_20),
.B1(n_26),
.B2(n_23),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_114),
.B1(n_122),
.B2(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_101),
.B(n_115),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_110),
.C(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_94),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_65),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_30),
.B(n_20),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_55),
.C(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_55),
.C(n_45),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_117),
.Y(n_129)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_51),
.B1(n_54),
.B2(n_71),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_42),
.B1(n_17),
.B2(n_27),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_86),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_90),
.B1(n_98),
.B2(n_62),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_133),
.B1(n_135),
.B2(n_148),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_26),
.C(n_20),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_147),
.C(n_103),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_143),
.B1(n_150),
.B2(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_79),
.B1(n_76),
.B2(n_63),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_93),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_58),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_144),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_152),
.B(n_22),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_114),
.B1(n_116),
.B2(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_32),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_154),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_74),
.C(n_39),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_63),
.B1(n_81),
.B2(n_27),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_87),
.B1(n_39),
.B2(n_41),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_0),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_77),
.B1(n_41),
.B2(n_39),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_106),
.B1(n_119),
.B2(n_41),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_32),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_159),
.B1(n_139),
.B2(n_138),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_154),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_158),
.Y(n_188)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_105),
.B1(n_106),
.B2(n_104),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_151),
.B1(n_145),
.B2(n_135),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_165),
.B(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_168),
.Y(n_192)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_36),
.B(n_25),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_172),
.C(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_177),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_153),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_99),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_173),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_140),
.B(n_32),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_16),
.C(n_13),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_0),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_182),
.B(n_31),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_41),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_128),
.B1(n_129),
.B2(n_152),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_28),
.B(n_25),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_133),
.B(n_39),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_129),
.C(n_128),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_145),
.A3(n_152),
.B1(n_149),
.B2(n_22),
.Y(n_187)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_191),
.A2(n_193),
.B1(n_203),
.B2(n_206),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_194),
.B(n_195),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_213),
.B(n_216),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_182),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_208),
.C(n_211),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_155),
.B1(n_21),
.B2(n_31),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_36),
.B(n_28),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_204),
.A2(n_1),
.B(n_2),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_36),
.B1(n_25),
.B2(n_24),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_169),
.B1(n_167),
.B2(n_163),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_23),
.C(n_30),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_227),
.B1(n_199),
.B2(n_204),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_186),
.B1(n_165),
.B2(n_166),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_174),
.B1(n_178),
.B2(n_177),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_174),
.B1(n_184),
.B2(n_1),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_226),
.A2(n_207),
.B(n_202),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_30),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_233),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_201),
.C(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_238),
.C(n_242),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_30),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_243),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_30),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_212),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_208),
.C(n_198),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_30),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_239),
.B1(n_220),
.B2(n_232),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_216),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_257),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_202),
.B(n_210),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_222),
.B1(n_190),
.B2(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_210),
.C(n_190),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_254),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_264),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_238),
.B1(n_221),
.B2(n_219),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_257),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_245),
.C(n_261),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_247),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_258),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_247),
.B1(n_249),
.B2(n_244),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_244),
.B1(n_251),
.B2(n_259),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_245),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_236),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_290),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_293),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_264),
.CI(n_265),
.CON(n_290),
.SN(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_234),
.C(n_248),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_297),
.C(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_296),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_243),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_251),
.C(n_189),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_226),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_292),
.A2(n_276),
.B1(n_274),
.B2(n_278),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_266),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_230),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_11),
.C(n_12),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_267),
.B1(n_6),
.B2(n_7),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_288),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_5),
.B(n_8),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_9),
.B(n_10),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_314),
.B(n_316),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_286),
.B(n_10),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_310),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_286),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_9),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_11),
.Y(n_322)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_309),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_325),
.B(n_327),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_306),
.Y(n_328)
);

AOI21x1_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_306),
.B(n_318),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_326),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_313),
.B(n_302),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_315),
.B(n_300),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_334),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_332),
.B(n_13),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_12),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_12),
.B(n_16),
.Y(n_339)
);


endmodule