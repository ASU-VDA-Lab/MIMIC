module fake_jpeg_3592_n_555 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_555);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_555;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_52),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_54),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_61),
.Y(n_127)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_64),
.B(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_30),
.B(n_0),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_96),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_67),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_29),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_1),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_77),
.B(n_80),
.Y(n_151)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_2),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_40),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_85),
.Y(n_156)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

CKINVDCx9p33_ASAP7_75t_R g90 ( 
.A(n_21),
.Y(n_90)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_31),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_16),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_95),
.Y(n_119)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx4f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_99),
.Y(n_131)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_100),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_102),
.B(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_43),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_28),
.B1(n_36),
.B2(n_33),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_106),
.A2(n_117),
.B1(n_143),
.B2(n_147),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_24),
.B1(n_47),
.B2(n_46),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_107),
.A2(n_109),
.B1(n_124),
.B2(n_136),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_28),
.B1(n_37),
.B2(n_32),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_108),
.A2(n_134),
.B1(n_165),
.B2(n_92),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_50),
.B1(n_25),
.B2(n_24),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_56),
.B(n_43),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_114),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_36),
.B1(n_42),
.B2(n_27),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_50),
.B1(n_24),
.B2(n_25),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_138),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_32),
.B1(n_49),
.B2(n_37),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_75),
.A2(n_50),
.B1(n_25),
.B2(n_46),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_47),
.C(n_46),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_91),
.A2(n_42),
.B1(n_33),
.B2(n_47),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_68),
.A2(n_49),
.B1(n_29),
.B2(n_43),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_83),
.A2(n_48),
.B1(n_19),
.B2(n_4),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_150),
.B1(n_57),
.B2(n_87),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_19),
.B1(n_3),
.B2(n_5),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_67),
.B1(n_54),
.B2(n_86),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_154),
.A2(n_15),
.B1(n_144),
.B2(n_148),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_2),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_3),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_62),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_159),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_66),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_52),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_168),
.A2(n_178),
.B1(n_227),
.B2(n_228),
.Y(n_280)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_169),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_171),
.B(n_176),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_70),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_172),
.B(n_181),
.Y(n_236)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_173),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_175),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_101),
.B1(n_97),
.B2(n_69),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_177),
.A2(n_192),
.B1(n_195),
.B2(n_204),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_88),
.B1(n_81),
.B2(n_100),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_6),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_179),
.Y(n_259)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_7),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_133),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_190),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_7),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_185),
.B(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_7),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_187),
.Y(n_263)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_119),
.B(n_8),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_191),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_127),
.B(n_10),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_193),
.B(n_203),
.Y(n_250)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_114),
.A2(n_92),
.B1(n_96),
.B2(n_19),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_10),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_11),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_199),
.B(n_201),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_129),
.B(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_206),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_11),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_12),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_202),
.B(n_205),
.C(n_209),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_123),
.B(n_12),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_16),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_12),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_113),
.B(n_13),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_113),
.B(n_14),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_15),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_217),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_132),
.B(n_15),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_221),
.Y(n_242)
);

BUFx2_ASAP7_75t_SL g215 ( 
.A(n_145),
.Y(n_215)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_122),
.B(n_15),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_219),
.A2(n_180),
.B1(n_184),
.B2(n_201),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_132),
.B(n_164),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_116),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_105),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_138),
.A2(n_159),
.B1(n_165),
.B2(n_121),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_126),
.A2(n_131),
.B1(n_109),
.B2(n_136),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_146),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_218),
.B(n_170),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_234),
.A2(n_274),
.B(n_190),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_197),
.A2(n_170),
.B1(n_220),
.B2(n_168),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_255),
.B1(n_273),
.B2(n_276),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_243),
.B(n_258),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_135),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_176),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_203),
.B(n_220),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_252),
.A2(n_262),
.B(n_202),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_197),
.A2(n_126),
.B1(n_135),
.B2(n_152),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_187),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_170),
.A2(n_145),
.B(n_146),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_150),
.B1(n_152),
.B2(n_141),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_265),
.A2(n_279),
.B1(n_188),
.B2(n_207),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_171),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_267),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_186),
.A2(n_130),
.B(n_115),
.C(n_163),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_269),
.A2(n_223),
.B(n_205),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_196),
.A2(n_130),
.B1(n_141),
.B2(n_140),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_196),
.A2(n_118),
.B(n_111),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_198),
.A2(n_110),
.B1(n_112),
.B2(n_125),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_224),
.A2(n_110),
.B1(n_112),
.B2(n_125),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_177),
.B1(n_195),
.B2(n_208),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_192),
.A2(n_115),
.B1(n_161),
.B2(n_105),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_286),
.B(n_296),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_290),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_199),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_307),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_293),
.A2(n_301),
.B1(n_314),
.B2(n_318),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_182),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_294),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_232),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_238),
.B(n_193),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_297),
.B(n_319),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_242),
.B(n_243),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_310),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_299),
.A2(n_317),
.B(n_320),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_234),
.A2(n_244),
.B1(n_265),
.B2(n_235),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_190),
.B1(n_179),
.B2(n_214),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_303),
.A2(n_313),
.B1(n_231),
.B2(n_230),
.Y(n_337)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_179),
.C(n_199),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_329),
.C(n_231),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_251),
.B(n_210),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_210),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_311),
.B(n_312),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_281),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_244),
.A2(n_209),
.B1(n_201),
.B2(n_205),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_279),
.A2(n_271),
.B1(n_246),
.B2(n_247),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_274),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_326),
.B(n_330),
.Y(n_347)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_245),
.B(n_194),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_209),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_247),
.B(n_202),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_189),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_324),
.B(n_332),
.Y(n_338)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_270),
.A2(n_173),
.B(n_222),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_246),
.A2(n_191),
.B1(n_207),
.B2(n_183),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_327),
.A2(n_328),
.B1(n_276),
.B2(n_277),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_230),
.A2(n_191),
.B1(n_208),
.B2(n_226),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_216),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_269),
.A2(n_213),
.B(n_225),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_118),
.B(n_175),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_283),
.B(n_169),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_259),
.B(n_187),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_239),
.Y(n_333)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

INVx11_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_337),
.A2(n_364),
.B1(n_299),
.B2(n_332),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_323),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_231),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_345),
.C(n_362),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_253),
.C(n_266),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_288),
.A2(n_255),
.B1(n_273),
.B2(n_256),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_346),
.A2(n_348),
.B1(n_361),
.B2(n_370),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_295),
.A2(n_301),
.B1(n_302),
.B2(n_304),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_354),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_298),
.B(n_250),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_352),
.B(n_300),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_289),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_292),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_289),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_331),
.Y(n_356)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_288),
.A2(n_256),
.B1(n_258),
.B2(n_266),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_233),
.C(n_240),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_233),
.C(n_240),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_372),
.C(n_153),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_313),
.A2(n_263),
.B1(n_212),
.B2(n_153),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_295),
.A2(n_254),
.B(n_268),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_368),
.A2(n_326),
.B(n_254),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_303),
.A2(n_263),
.B1(n_212),
.B2(n_264),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_290),
.B(n_241),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_285),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_309),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_361),
.A2(n_314),
.B1(n_330),
.B2(n_317),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_379),
.A2(n_384),
.B1(n_385),
.B2(n_392),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_340),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_380),
.B(n_393),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

FAx1_ASAP7_75t_SL g382 ( 
.A(n_352),
.B(n_306),
.CI(n_315),
.CON(n_382),
.SN(n_382)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_382),
.B(n_400),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_383),
.A2(n_386),
.B(n_409),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_315),
.B1(n_293),
.B2(n_324),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_369),
.A2(n_308),
.B(n_316),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_411),
.C(n_415),
.Y(n_433)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_367),
.A2(n_287),
.B1(n_310),
.B2(n_322),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_390),
.A2(n_391),
.B1(n_414),
.B2(n_370),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_349),
.A2(n_325),
.B1(n_305),
.B2(n_291),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_346),
.A2(n_329),
.B1(n_327),
.B2(n_307),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_L g393 ( 
.A1(n_369),
.A2(n_334),
.B(n_284),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_335),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_398),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_309),
.B1(n_285),
.B2(n_263),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_396),
.A2(n_405),
.B1(n_354),
.B2(n_355),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_397),
.B(n_403),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_351),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_284),
.Y(n_400)
);

BUFx12f_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_407),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_402),
.B(n_345),
.Y(n_431)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_347),
.A2(n_264),
.B1(n_241),
.B2(n_161),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_358),
.B(n_174),
.Y(n_406)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_339),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g409 ( 
.A(n_358),
.B(n_268),
.CI(n_169),
.CON(n_409),
.SN(n_409)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_175),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_411),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_350),
.A2(n_174),
.B1(n_348),
.B2(n_366),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_343),
.B(n_174),
.C(n_341),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_417),
.A2(n_428),
.B1(n_444),
.B2(n_401),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_371),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_422),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_371),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_375),
.B(n_377),
.Y(n_426)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_414),
.A2(n_337),
.B1(n_350),
.B2(n_338),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_386),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_439),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_431),
.B(n_438),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_385),
.A2(n_376),
.B1(n_374),
.B2(n_368),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_437),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_372),
.C(n_362),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_440),
.C(n_441),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_384),
.A2(n_376),
.B1(n_374),
.B2(n_373),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_399),
.B(n_338),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_403),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_373),
.C(n_344),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_396),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_446),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_391),
.A2(n_408),
.B1(n_390),
.B2(n_410),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_410),
.A2(n_344),
.B1(n_355),
.B2(n_378),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_405),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_413),
.C(n_387),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_460),
.C(n_466),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_416),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_471),
.Y(n_481)
);

XNOR2x2_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_382),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_451),
.B(n_342),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_428),
.A2(n_410),
.B1(n_392),
.B2(n_383),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_453),
.A2(n_458),
.B1(n_463),
.B2(n_434),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_454),
.A2(n_443),
.B1(n_417),
.B2(n_442),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_397),
.B(n_395),
.Y(n_455)
);

AOI21x1_ASAP7_75t_SL g496 ( 
.A1(n_455),
.A2(n_467),
.B(n_465),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_433),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_469),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_444),
.A2(n_387),
.B1(n_395),
.B2(n_382),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_402),
.C(n_404),
.Y(n_460)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_SL g466 ( 
.A(n_432),
.B(n_409),
.C(n_401),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_419),
.B(n_409),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_474),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_425),
.B(n_401),
.Y(n_468)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_420),
.B(n_364),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_357),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_359),
.Y(n_472)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_357),
.C(n_359),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_445),
.C(n_441),
.Y(n_480)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_418),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_476),
.A2(n_461),
.B1(n_454),
.B2(n_465),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_468),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_489),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_485),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_437),
.Y(n_484)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_457),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_494),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_486),
.A2(n_487),
.B1(n_452),
.B2(n_493),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_453),
.A2(n_442),
.B1(n_446),
.B2(n_421),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_431),
.C(n_430),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_430),
.C(n_423),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_491),
.C(n_492),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_423),
.C(n_427),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_424),
.C(n_365),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_455),
.A2(n_365),
.B(n_342),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_495),
.A2(n_496),
.B(n_454),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_459),
.Y(n_499)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_514),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_512),
.Y(n_519)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_503),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_473),
.C(n_460),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_508),
.C(n_492),
.Y(n_520)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_505),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_461),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_506),
.B(n_510),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_507),
.A2(n_496),
.B(n_487),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_452),
.C(n_469),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_476),
.A2(n_458),
.B1(n_466),
.B2(n_464),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_482),
.A2(n_470),
.B(n_451),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_511),
.A2(n_488),
.B(n_495),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_489),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_517),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_516),
.A2(n_526),
.B(n_520),
.Y(n_537)
);

FAx1_ASAP7_75t_SL g517 ( 
.A(n_511),
.B(n_508),
.CI(n_475),
.CON(n_517),
.SN(n_517)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_523),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_486),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_521),
.B(n_522),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_483),
.C(n_494),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_483),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_502),
.B(n_484),
.C(n_512),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_527),
.B(n_509),
.Y(n_530)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_530),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_497),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_534),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_525),
.A2(n_513),
.B(n_504),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_519),
.C(n_522),
.Y(n_544)
);

NOR2xp67_ASAP7_75t_R g534 ( 
.A(n_524),
.B(n_500),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_527),
.A2(n_501),
.B1(n_510),
.B2(n_507),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_535),
.B(n_518),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_537),
.Y(n_543)
);

AOI211xp5_ASAP7_75t_L g538 ( 
.A1(n_516),
.A2(n_515),
.B(n_528),
.C(n_517),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_526),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_R g546 ( 
.A(n_539),
.B(n_532),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_529),
.C(n_518),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_536),
.Y(n_545)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_545),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_546),
.B(n_547),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_543),
.B(n_530),
.Y(n_548)
);

AO21x1_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_539),
.B(n_548),
.Y(n_551)
);

AO21x1_ASAP7_75t_L g553 ( 
.A1(n_551),
.A2(n_552),
.B(n_540),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_549),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_553),
.B(n_541),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_517),
.B(n_523),
.Y(n_555)
);


endmodule