module real_jpeg_17638_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_487;
wire n_93;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_536),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_0),
.B(n_537),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_1),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

AOI22x1_ASAP7_75t_SL g287 ( 
.A1(n_1),
.A2(n_123),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_1),
.A2(n_123),
.B1(n_233),
.B2(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_1),
.A2(n_123),
.B1(n_368),
.B2(n_493),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_2),
.A2(n_313),
.B1(n_317),
.B2(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_2),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_2),
.A2(n_318),
.B1(n_426),
.B2(n_429),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_2),
.A2(n_318),
.B1(n_485),
.B2(n_487),
.Y(n_484)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_89),
.B1(n_90),
.B2(n_94),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_4),
.A2(n_89),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_4),
.A2(n_89),
.B1(n_236),
.B2(n_239),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_4),
.A2(n_89),
.B1(n_377),
.B2(n_380),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_6),
.A2(n_274),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

OAI22x1_ASAP7_75t_SL g453 ( 
.A1(n_6),
.A2(n_274),
.B1(n_454),
.B2(n_456),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_6),
.A2(n_274),
.B1(n_526),
.B2(n_529),
.Y(n_525)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_7),
.Y(n_537)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_8),
.A2(n_103),
.B1(n_199),
.B2(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_8),
.A2(n_103),
.B1(n_385),
.B2(n_389),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_8),
.A2(n_103),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_9),
.Y(n_117)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_9),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_9),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_10),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_10),
.A2(n_132),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_10),
.A2(n_132),
.B1(n_240),
.B2(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_10),
.A2(n_132),
.B1(n_368),
.B2(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_11),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_11),
.Y(n_442)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_12),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_12),
.Y(n_360)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_13),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_13),
.B(n_87),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_47),
.B1(n_225),
.B2(n_230),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_248),
.A3(n_253),
.B1(n_254),
.B2(n_257),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_13),
.B(n_298),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g347 ( 
.A1(n_13),
.A2(n_226),
.A3(n_348),
.B1(n_352),
.B2(n_355),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_13),
.A2(n_47),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_14),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_15),
.A2(n_341),
.B1(n_344),
.B2(n_346),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_15),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_15),
.A2(n_31),
.B1(n_346),
.B2(n_440),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_15),
.A2(n_346),
.B1(n_512),
.B2(n_515),
.Y(n_511)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g351 ( 
.A(n_17),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_17),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_17),
.Y(n_369)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_17),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_503),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_468),
.B(n_500),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_400),
.B(n_465),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_326),
.B(n_399),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_279),
.B(n_325),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_192),
.B(n_278),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_145),
.B(n_191),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_96),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_29),
.B(n_96),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_53),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_30),
.A2(n_53),
.B1(n_54),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_30),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.A3(n_41),
.B1(n_46),
.B2(n_49),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_39),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_47),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_47),
.A2(n_108),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_47),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_47),
.B(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_87),
.B2(n_88),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_59),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_60),
.A2(n_87),
.B1(n_88),
.B2(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_60),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_60),
.B(n_394),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_64),
.Y(n_398)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_71),
.Y(n_253)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_73),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_73),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_73),
.B(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_73),
.A2(n_196),
.B1(n_438),
.B2(n_439),
.Y(n_437)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_81),
.B2(n_83),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_75),
.Y(n_182)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_81),
.Y(n_345)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_82),
.Y(n_276)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_87),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_87),
.B(n_425),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_126),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_97),
.B(n_127),
.C(n_136),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_108),
.B(n_113),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_106),
.Y(n_343)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_107),
.Y(n_273)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_108),
.A2(n_149),
.B1(n_172),
.B2(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_108),
.B(n_270),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_108),
.A2(n_118),
.B(n_475),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_114),
.B(n_319),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_118),
.Y(n_267)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_130),
.Y(n_289)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AO22x2_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_137),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_137),
.B(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_137),
.A2(n_414),
.B1(n_510),
.B2(n_511),
.Y(n_509)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_139),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_166),
.B(n_190),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_164),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_158),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_158),
.A2(n_312),
.B1(n_336),
.B2(n_340),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_158),
.A2(n_268),
.B(n_340),
.Y(n_422)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_163),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_183),
.B(n_189),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_182),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_187),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_277),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_193),
.B(n_277),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_246),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_208),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_195),
.B(n_208),
.C(n_246),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_196),
.A2(n_287),
.B(n_393),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_196),
.A2(n_393),
.B(n_439),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_202),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_203),
.Y(n_428)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_224),
.B1(n_235),
.B2(n_245),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_209),
.A2(n_235),
.B1(n_245),
.B2(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_209),
.A2(n_245),
.B1(n_321),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_209),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_209),
.A2(n_417),
.B(n_452),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_209),
.A2(n_245),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_214),
.B1(n_217),
.B2(n_220),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_214),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_215),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_216),
.Y(n_388)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_222),
.Y(n_459)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_222),
.Y(n_514)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_228),
.Y(n_354)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_228),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_238),
.Y(n_323)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_245),
.B(n_417),
.Y(n_416)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_266),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_266),
.Y(n_283)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_263),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_262),
.Y(n_391)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_262),
.Y(n_455)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_280),
.B(n_281),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_293),
.B1(n_294),
.B2(n_324),
.Y(n_281)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_284),
.C(n_293),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_286),
.B(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_320),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_306),
.B2(n_307),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_320),
.C(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_298),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_298),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_298),
.B(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_298),
.B(n_525),
.Y(n_524)
);

AO22x2_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_302),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_305),
.Y(n_365)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_312),
.B(n_319),
.Y(n_307)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx6_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_328),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_361),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_333),
.B2(n_334),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_331),
.B(n_333),
.C(n_361),
.Y(n_462)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_347),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_335),
.B(n_347),
.Y(n_419)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_351),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_360),
.A2(n_365),
.B1(n_366),
.B2(n_368),
.Y(n_364)
);

XOR2x2_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_382),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_383),
.C(n_392),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_370),
.B1(n_376),
.B2(n_381),
.Y(n_362)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

OAI22x1_ASAP7_75t_SL g447 ( 
.A1(n_363),
.A2(n_381),
.B1(n_410),
.B2(n_448),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_363),
.A2(n_448),
.B(n_491),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_363),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx8_ASAP7_75t_L g495 ( 
.A(n_374),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_375),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_376),
.Y(n_407)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_378),
.Y(n_450)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_379),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_380),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

INVx3_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_461),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_432),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_403),
.B(n_432),
.C(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_420),
.C(n_421),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_404),
.B(n_464),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_419),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_413),
.C(n_419),
.Y(n_433)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B(n_416),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_421),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_423),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_431),
.Y(n_423)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_443),
.C(n_460),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_443),
.B1(n_444),
.B2(n_460),
.Y(n_434)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_436),
.B(n_437),
.Y(n_496)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_447),
.C(n_451),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_459),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_463),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_470),
.B(n_471),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_472),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_480),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_473),
.B(n_480),
.C(n_497),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_473)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_474),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_474),
.A2(n_479),
.B1(n_522),
.B2(n_530),
.Y(n_521)
);

NOR2x1_ASAP7_75t_R g531 ( 
.A(n_474),
.B(n_478),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2x1_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_496),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_490),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_490),
.C(n_496),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_492),
.Y(n_523)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g503 ( 
.A(n_504),
.B(n_535),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_534),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_534),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_520),
.B1(n_532),
.B2(n_533),
.Y(n_507)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

OAI21xp33_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_517),
.B(n_519),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_517),
.Y(n_519)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_520),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_531),
.Y(n_520)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_522),
.Y(n_530)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);


endmodule