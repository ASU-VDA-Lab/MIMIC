module fake_ariane_1717_n_2171 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2171);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2171;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_145),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_127),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_47),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_152),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_120),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_53),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_0),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_64),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_74),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_209),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_199),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_87),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_51),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_34),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_75),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_158),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_71),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_16),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_72),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_59),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_143),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_84),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_94),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_128),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_69),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_69),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_86),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_150),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_29),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_27),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_151),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_35),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_51),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_35),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_213),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_82),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_200),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_8),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_173),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_6),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_121),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_107),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_206),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_18),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_103),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_101),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_201),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_46),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_210),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_142),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_27),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_58),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_31),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_222),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_122),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_168),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_115),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_38),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_137),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_112),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_98),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_6),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_39),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_12),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_116),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_89),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_141),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_17),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_133),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_74),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_68),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_108),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_34),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_149),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_109),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_154),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_114),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_92),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_78),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_29),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_186),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_205),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_54),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_25),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_148),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_134),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_104),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_11),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_48),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_130),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_138),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_118),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_110),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_221),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_41),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_36),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_50),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_119),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_90),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_91),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_140),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_188),
.Y(n_355)
);

BUFx8_ASAP7_75t_SL g356 ( 
.A(n_40),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_102),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_38),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_44),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_159),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_117),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_124),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_1),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_180),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_53),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_48),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_163),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_106),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_67),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_24),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_166),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_49),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_167),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_214),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_105),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_223),
.Y(n_376)
);

BUFx8_ASAP7_75t_SL g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_85),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_40),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_192),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_125),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_129),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_100),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_23),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_81),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_79),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_62),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_181),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_57),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_66),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_160),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_26),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_24),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_170),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_136),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_37),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_97),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_126),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_55),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_196),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_220),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_30),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_219),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_83),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_66),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_64),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_75),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_203),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_135),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_3),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_39),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_16),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_70),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_123),
.Y(n_414)
);

BUFx2_ASAP7_75t_SL g415 ( 
.A(n_211),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_59),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_54),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_187),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_155),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_43),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_215),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_20),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_174),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_71),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_161),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_9),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_46),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_2),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_172),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_157),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_12),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_146),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_164),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_132),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_32),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_93),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_13),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_56),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_50),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_73),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_197),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_67),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_10),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_72),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_399),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_251),
.B(n_1),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_264),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_251),
.B(n_2),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_356),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_271),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_236),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_246),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_264),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_279),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_236),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_272),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_334),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_334),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_262),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_279),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_229),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_229),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_235),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_262),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_262),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_266),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_262),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_235),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_273),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_389),
.B(n_3),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_333),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_273),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_275),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_333),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_307),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_275),
.B(n_4),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_285),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_230),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_267),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_239),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_287),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_239),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_255),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_329),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_255),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_256),
.Y(n_487)
);

INVxp33_ASAP7_75t_SL g488 ( 
.A(n_327),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_256),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_307),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_265),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_265),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_386),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_419),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_307),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_268),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_268),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_307),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_430),
.B(n_4),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_269),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_315),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_269),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_260),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_276),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_332),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_389),
.B(n_5),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_402),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_416),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_276),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_428),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_233),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_289),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_289),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_243),
.B(n_10),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_332),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_237),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_377),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_285),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_361),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_332),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_293),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_332),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_240),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_260),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_293),
.Y(n_525)
);

BUFx2_ASAP7_75t_SL g526 ( 
.A(n_290),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_301),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_301),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_303),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_242),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_303),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_281),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_247),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_281),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_309),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_291),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_249),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_288),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_309),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_288),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_292),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_252),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_314),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_292),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_253),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_257),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_291),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_312),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_312),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_314),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_320),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_320),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_R g553 ( 
.A(n_226),
.B(n_77),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_272),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_336),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_243),
.B(n_11),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_272),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_336),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_350),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_228),
.B(n_182),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_350),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_406),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_406),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_258),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_518),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_517),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_501),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_507),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_462),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_463),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_453),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_463),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_508),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_526),
.B(n_306),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_464),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_460),
.B(n_231),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_467),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_488),
.B(n_346),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_469),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_480),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_526),
.B(n_306),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_510),
.Y(n_585)
);

AND2x6_ASAP7_75t_L g586 ( 
.A(n_470),
.B(n_346),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_447),
.B(n_313),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_470),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_454),
.B(n_313),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_482),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_455),
.B(n_406),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_473),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_461),
.B(n_431),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_474),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_481),
.B(n_431),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_539),
.B(n_431),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_452),
.B(n_227),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_474),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_478),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_485),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_478),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_493),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_494),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_503),
.B(n_410),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_449),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_511),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_538),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_540),
.B(n_346),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_540),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_541),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_519),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_541),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_445),
.B(n_259),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_503),
.B(n_460),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_530),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_465),
.B(n_466),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_544),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_544),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_483),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_484),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_486),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_458),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_487),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_543),
.B(n_410),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_489),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_491),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_533),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_514),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_492),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_451),
.B(n_358),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_496),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_524),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_500),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_502),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_488),
.B(n_305),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_532),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_533),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_509),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_458),
.A2(n_396),
.B1(n_411),
.B2(n_323),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_512),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_513),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_537),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_521),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_537),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_525),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_545),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_527),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_528),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_465),
.B(n_466),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_534),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_456),
.B(n_358),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_468),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_628),
.B(n_514),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_566),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_618),
.B(n_468),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_566),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_600),
.B(n_446),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_620),
.B(n_476),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_639),
.B(n_476),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_566),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_595),
.B(n_490),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_654),
.B(n_490),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_632),
.B(n_495),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_570),
.B(n_495),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_570),
.B(n_498),
.Y(n_671)
);

NAND3x1_ASAP7_75t_L g672 ( 
.A(n_598),
.B(n_448),
.C(n_499),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_595),
.B(n_498),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_628),
.B(n_497),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_595),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_570),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_570),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_574),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_566),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_566),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_593),
.B(n_319),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_574),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_570),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_595),
.B(n_505),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_619),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_628),
.B(n_555),
.Y(n_687)
);

AO21x2_ASAP7_75t_L g688 ( 
.A1(n_576),
.A2(n_506),
.B(n_471),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_632),
.B(n_505),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_577),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_570),
.B(n_515),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_631),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_590),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_632),
.B(n_515),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_590),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_566),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_632),
.B(n_520),
.Y(n_697)
);

AO21x2_ASAP7_75t_L g698 ( 
.A1(n_584),
.A2(n_326),
.B(n_319),
.Y(n_698)
);

BUFx4f_ASAP7_75t_L g699 ( 
.A(n_590),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_577),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_626),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_581),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_567),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_598),
.A2(n_459),
.B1(n_522),
.B2(n_520),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_590),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_590),
.B(n_522),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_597),
.Y(n_707)
);

OAI21xp33_ASAP7_75t_SL g708 ( 
.A1(n_581),
.A2(n_477),
.B(n_556),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_599),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_597),
.B(n_459),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_593),
.B(n_326),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_599),
.A2(n_546),
.B1(n_564),
.B2(n_545),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_597),
.B(n_601),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_590),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_578),
.B(n_641),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_614),
.B(n_340),
.Y(n_716)
);

INVxp67_ASAP7_75t_SL g717 ( 
.A(n_597),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_614),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_614),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_614),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_647),
.B(n_564),
.C(n_546),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_614),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_588),
.B(n_516),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_582),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_614),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_586),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_601),
.B(n_602),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_591),
.B(n_523),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_626),
.B(n_457),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_587),
.B(n_557),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_602),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_601),
.B(n_340),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_601),
.B(n_542),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_610),
.B(n_450),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_604),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_604),
.B(n_536),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_628),
.A2(n_363),
.B1(n_365),
.B2(n_359),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_613),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_609),
.B(n_547),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_649),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_586),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_586),
.A2(n_363),
.B1(n_365),
.B2(n_359),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_624),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_609),
.B(n_531),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_624),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_611),
.B(n_548),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_586),
.A2(n_372),
.B1(n_387),
.B2(n_370),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_613),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_611),
.B(n_343),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_636),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_651),
.A2(n_277),
.B1(n_282),
.B2(n_274),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_616),
.B(n_535),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_589),
.B(n_472),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_616),
.B(n_343),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_612),
.A2(n_347),
.B(n_345),
.Y(n_757)
);

BUFx4f_ASAP7_75t_L g758 ( 
.A(n_643),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_586),
.A2(n_372),
.B1(n_387),
.B2(n_370),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_655),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_621),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_622),
.B(n_550),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_622),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_640),
.B(n_475),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_643),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_643),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_596),
.B(n_345),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_596),
.B(n_551),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_565),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_634),
.B(n_549),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_565),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_634),
.B(n_552),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_656),
.B(n_294),
.C(n_284),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_630),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_656),
.B(n_558),
.Y(n_775)
);

AND3x4_ASAP7_75t_L g776 ( 
.A(n_624),
.B(n_562),
.C(n_554),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_586),
.A2(n_417),
.B1(n_420),
.B2(n_393),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_637),
.B(n_559),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_637),
.B(n_561),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_637),
.B(n_617),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_607),
.B(n_393),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_630),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_SL g783 ( 
.A(n_644),
.B(n_563),
.Y(n_783)
);

BUFx10_ASAP7_75t_L g784 ( 
.A(n_615),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_645),
.B(n_646),
.Y(n_785)
);

AND2x2_ASAP7_75t_SL g786 ( 
.A(n_573),
.B(n_238),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_572),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_586),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_573),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_645),
.B(n_432),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_643),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_594),
.A2(n_417),
.B1(n_420),
.B2(n_443),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_645),
.B(n_347),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_607),
.B(n_443),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_594),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_643),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_607),
.B(n_298),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_607),
.B(n_355),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_643),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_633),
.Y(n_800)
);

INVx4_ASAP7_75t_SL g801 ( 
.A(n_623),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_579),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_645),
.A2(n_366),
.B1(n_444),
.B2(n_442),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_633),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_623),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_608),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_568),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_646),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_633),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_646),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_650),
.B(n_355),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_665),
.B(n_650),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_658),
.B(n_650),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_769),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_710),
.A2(n_650),
.B(n_625),
.C(n_629),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_730),
.B(n_583),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_769),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_658),
.B(n_625),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_664),
.B(n_657),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_627),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_810),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_738),
.A2(n_644),
.B1(n_653),
.B2(n_652),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_709),
.B(n_627),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_764),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_668),
.B(n_629),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_696),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_810),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_661),
.B(n_724),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_661),
.B(n_724),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_SL g831 ( 
.A(n_668),
.B(n_635),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_770),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_744),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_729),
.B(n_635),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_771),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_729),
.B(n_657),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_669),
.B(n_638),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_682),
.A2(n_648),
.B1(n_638),
.B2(n_612),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_727),
.B(n_642),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_682),
.A2(n_648),
.B1(n_652),
.B2(n_653),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_SL g842 ( 
.A1(n_783),
.A2(n_606),
.B1(n_605),
.B2(n_603),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_669),
.B(n_642),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_678),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_810),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_735),
.B(n_592),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_679),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_689),
.B(n_642),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_708),
.A2(n_653),
.B(n_652),
.C(n_373),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_689),
.B(n_360),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_694),
.B(n_360),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_694),
.B(n_367),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_701),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_738),
.A2(n_381),
.B1(n_394),
.B2(n_367),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_727),
.B(n_338),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_742),
.B(n_371),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_683),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_780),
.B(n_569),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_772),
.B(n_575),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_810),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_690),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_697),
.B(n_371),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_697),
.B(n_373),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_700),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_768),
.B(n_778),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_682),
.A2(n_376),
.B1(n_380),
.B2(n_381),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_667),
.B(n_299),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_673),
.B(n_300),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_738),
.A2(n_394),
.B1(n_421),
.B2(n_376),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_702),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_742),
.B(n_380),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_768),
.B(n_385),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_685),
.A2(n_672),
.B1(n_707),
.B2(n_675),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_772),
.B(n_585),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_788),
.B(n_385),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_778),
.B(n_421),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_731),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_718),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_779),
.B(n_433),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_754),
.B(n_302),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_807),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_674),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_725),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_779),
.B(n_433),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_682),
.B(n_308),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_712),
.B(n_553),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_674),
.B(n_316),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_704),
.B(n_560),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_737),
.B(n_322),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_740),
.B(n_325),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_682),
.B(n_330),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_711),
.B(n_337),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_732),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_811),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_788),
.B(n_290),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_739),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_747),
.B(n_341),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_715),
.B(n_342),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_736),
.Y(n_899)
);

NAND2x1_ASAP7_75t_L g900 ( 
.A(n_808),
.B(n_809),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_674),
.B(n_687),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_756),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_761),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_808),
.B(n_310),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_711),
.B(n_348),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_739),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_715),
.B(n_349),
.Y(n_907)
);

INVxp67_ASAP7_75t_SL g908 ( 
.A(n_744),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_711),
.B(n_369),
.Y(n_909)
);

NOR2x2_ASAP7_75t_L g910 ( 
.A(n_686),
.B(n_379),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_711),
.B(n_384),
.Y(n_911)
);

O2A1O1Ixp5_ASAP7_75t_L g912 ( 
.A1(n_733),
.A2(n_441),
.B(n_244),
.C(n_248),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_722),
.B(n_310),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_711),
.B(n_390),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_734),
.B(n_392),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_763),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_809),
.B(n_404),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_787),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_663),
.A2(n_404),
.B1(n_415),
.B2(n_441),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_749),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_767),
.B(n_405),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_746),
.B(n_407),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_767),
.B(n_412),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_767),
.A2(n_415),
.B1(n_232),
.B2(n_368),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_687),
.Y(n_925)
);

O2A1O1Ixp5_ASAP7_75t_L g926 ( 
.A1(n_733),
.A2(n_238),
.B(n_244),
.C(n_248),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_802),
.B(n_261),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_767),
.B(n_413),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_767),
.B(n_422),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_805),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_717),
.A2(n_261),
.B(n_280),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_749),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_785),
.B(n_424),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_663),
.A2(n_382),
.B1(n_324),
.B2(n_280),
.Y(n_934)
);

INVx8_ASAP7_75t_L g935 ( 
.A(n_772),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_728),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_751),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_792),
.A2(n_382),
.B1(n_324),
.B2(n_438),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_785),
.B(n_426),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_792),
.A2(n_440),
.B1(n_439),
.B2(n_437),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_786),
.B(n_427),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_746),
.B(n_317),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_713),
.A2(n_354),
.B(n_241),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_775),
.B(n_435),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_786),
.A2(n_317),
.B1(n_374),
.B2(n_429),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_789),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_745),
.B(n_234),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_743),
.A2(n_317),
.B1(n_374),
.B2(n_425),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_775),
.B(n_245),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_745),
.B(n_250),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_741),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_760),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_686),
.B(n_14),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_721),
.B(n_374),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_703),
.B(n_15),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_670),
.A2(n_436),
.B1(n_434),
.B2(n_423),
.Y(n_956)
);

OAI221xp5_ASAP7_75t_L g957 ( 
.A1(n_659),
.A2(n_418),
.B1(n_414),
.B2(n_409),
.C(n_408),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_670),
.A2(n_403),
.B1(n_401),
.B2(n_400),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_798),
.B(n_317),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_741),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_753),
.B(n_254),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_795),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_721),
.B(n_374),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_774),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_753),
.B(n_263),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_800),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_659),
.B(n_15),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_773),
.B(n_17),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_804),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_782),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_686),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_692),
.B(n_19),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_721),
.B(n_723),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_762),
.B(n_270),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_752),
.B(n_19),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_811),
.B(n_20),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_804),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_692),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_762),
.B(n_278),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_L g980 ( 
.A(n_829),
.B(n_691),
.C(n_671),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_830),
.B(n_671),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_865),
.A2(n_706),
.B(n_691),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_843),
.A2(n_706),
.B(n_699),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_819),
.B(n_775),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_848),
.A2(n_699),
.B(n_758),
.Y(n_985)
);

AO22x1_ASAP7_75t_L g986 ( 
.A1(n_846),
.A2(n_776),
.B1(n_874),
.B2(n_859),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_819),
.B(n_798),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_825),
.B(n_692),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_880),
.B(n_784),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_814),
.A2(n_758),
.B(n_693),
.Y(n_990)
);

AOI21x1_ASAP7_75t_L g991 ( 
.A1(n_973),
.A2(n_799),
.B(n_796),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_834),
.A2(n_803),
.B(n_812),
.C(n_793),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_821),
.B(n_798),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_821),
.B(n_790),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_900),
.A2(n_917),
.B(n_904),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_930),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_827),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_820),
.A2(n_743),
.B1(n_759),
.B2(n_748),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_904),
.A2(n_693),
.B(n_677),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_836),
.B(n_797),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_896),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_827),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_906),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_920),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_915),
.B(n_826),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_917),
.A2(n_677),
.B(n_684),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_915),
.B(n_781),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_859),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_932),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_826),
.B(n_781),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_813),
.A2(n_705),
.B(n_714),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_850),
.A2(n_748),
.B1(n_759),
.B2(n_777),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_840),
.A2(n_676),
.B(n_684),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_851),
.A2(n_755),
.B(n_750),
.C(n_716),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_813),
.B(n_781),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_877),
.B(n_688),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_827),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_849),
.A2(n_714),
.B(n_719),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_919),
.A2(n_688),
.B1(n_794),
.B2(n_777),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_874),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_852),
.A2(n_755),
.B(n_750),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_827),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_881),
.B(n_784),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_894),
.B(n_721),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_824),
.B(n_698),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_840),
.A2(n_676),
.B(n_705),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_954),
.A2(n_662),
.B(n_666),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_824),
.B(n_698),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_973),
.A2(n_719),
.B(n_799),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_844),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_936),
.A2(n_796),
.B(n_720),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_867),
.B(n_801),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_822),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_882),
.B(n_695),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_954),
.A2(n_662),
.B(n_666),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_867),
.B(n_801),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_862),
.A2(n_726),
.B1(n_720),
.B2(n_695),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_858),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_838),
.A2(n_726),
.B(n_680),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_968),
.A2(n_716),
.B(n_681),
.C(n_660),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_960),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_855),
.A2(n_660),
.B(n_680),
.Y(n_1043)
);

NAND2x1p5_ASAP7_75t_L g1044 ( 
.A(n_925),
.B(n_765),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_847),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_966),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_894),
.B(n_723),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_855),
.A2(n_681),
.B(n_723),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_857),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_832),
.B(n_784),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_868),
.B(n_801),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_868),
.B(n_757),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_889),
.B(n_757),
.Y(n_1053)
);

NOR2x1_ASAP7_75t_L g1054 ( 
.A(n_955),
.B(n_776),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_863),
.A2(n_723),
.B1(n_765),
.B2(n_766),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_968),
.A2(n_766),
.B(n_765),
.C(n_791),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_927),
.B(n_765),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_895),
.A2(n_791),
.B(n_766),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_895),
.A2(n_791),
.B(n_766),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_873),
.A2(n_791),
.B(n_696),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_889),
.B(n_696),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_816),
.A2(n_696),
.B(n_283),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_831),
.A2(n_286),
.B(n_398),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_890),
.B(n_806),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_969),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_842),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_890),
.B(n_806),
.Y(n_1067)
);

OAI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_897),
.A2(n_351),
.B(n_397),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_897),
.B(n_806),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_856),
.A2(n_875),
.B(n_871),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_977),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_934),
.B(n_295),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_886),
.B(n_395),
.C(n_391),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_828),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_919),
.A2(n_317),
.B(n_383),
.C(n_378),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_963),
.A2(n_374),
.B(n_375),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_872),
.A2(n_388),
.B1(n_364),
.B2(n_362),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_975),
.A2(n_374),
.B1(n_357),
.B2(n_353),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_858),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_934),
.B(n_297),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_935),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_947),
.B(n_304),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_950),
.B(n_311),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_888),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_894),
.B(n_374),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_856),
.A2(n_335),
.B(n_352),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_871),
.A2(n_344),
.B(n_339),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_861),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_887),
.B(n_21),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_933),
.A2(n_22),
.B(n_26),
.C(n_28),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_961),
.B(n_318),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_875),
.A2(n_331),
.B(n_328),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_815),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_853),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_L g1095 ( 
.A1(n_963),
.A2(n_374),
.B(n_321),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_965),
.B(n_30),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_817),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_935),
.A2(n_374),
.B1(n_32),
.B2(n_33),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_841),
.A2(n_96),
.B(n_218),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_935),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_864),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_967),
.B(n_31),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_941),
.B(n_33),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_974),
.B(n_870),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_943),
.A2(n_99),
.B(n_216),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_937),
.B(n_36),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_939),
.A2(n_95),
.B(n_212),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_918),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_944),
.B(n_37),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_878),
.B(n_883),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_833),
.A2(n_111),
.B(n_207),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_818),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_908),
.A2(n_88),
.B(n_202),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_893),
.B(n_41),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_899),
.A2(n_902),
.B(n_903),
.C(n_916),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_951),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_922),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_931),
.A2(n_113),
.B(n_198),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_976),
.A2(n_42),
.B(n_45),
.C(n_47),
.Y(n_1119)
);

CKINVDCx11_ASAP7_75t_R g1120 ( 
.A(n_927),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_845),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_835),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_922),
.B(n_52),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_945),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_971),
.B(n_57),
.Y(n_1125)
);

NOR2x1p5_ASAP7_75t_SL g1126 ( 
.A(n_894),
.B(n_153),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_854),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_860),
.A2(n_162),
.B(n_194),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_952),
.B(n_60),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_959),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_979),
.A2(n_169),
.B(n_193),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_837),
.A2(n_139),
.B(n_191),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_959),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_946),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_978),
.B(n_131),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_898),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_962),
.A2(n_80),
.B(n_190),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_894),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_949),
.A2(n_224),
.B(n_185),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_876),
.A2(n_184),
.B(n_183),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_839),
.A2(n_912),
.B(n_926),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_854),
.A2(n_61),
.B(n_63),
.C(n_65),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_927),
.B(n_63),
.Y(n_1143)
);

OAI321xp33_ASAP7_75t_L g1144 ( 
.A1(n_940),
.A2(n_869),
.A3(n_938),
.B1(n_948),
.B2(n_866),
.C(n_945),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_964),
.A2(n_171),
.B(n_175),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_953),
.B(n_972),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_938),
.B(n_68),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_879),
.B(n_70),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_970),
.B(n_73),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_884),
.A2(n_76),
.B(n_976),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_894),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_959),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_885),
.A2(n_914),
.B(n_929),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_957),
.A2(n_907),
.B(n_905),
.C(n_911),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_869),
.B(n_76),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_959),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_891),
.A2(n_921),
.B(n_892),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_909),
.A2(n_928),
.B(n_923),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_823),
.B(n_940),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_823),
.B(n_898),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_924),
.A2(n_913),
.B(n_942),
.Y(n_1161)
);

AO21x1_ASAP7_75t_L g1162 ( 
.A1(n_942),
.A2(n_956),
.B(n_958),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_959),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_948),
.Y(n_1164)
);

AND3x1_ASAP7_75t_L g1165 ( 
.A(n_910),
.B(n_846),
.C(n_783),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1100),
.B(n_1081),
.Y(n_1166)
);

AOI222xp33_ASAP7_75t_L g1167 ( 
.A1(n_1159),
.A2(n_986),
.B1(n_1144),
.B2(n_1160),
.C1(n_984),
.C2(n_998),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_984),
.B(n_1097),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1001),
.B(n_1006),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1081),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1001),
.B(n_994),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_991),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_SL g1173 ( 
.A1(n_1150),
.A2(n_1022),
.B(n_1105),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1052),
.A2(n_1053),
.B(n_1153),
.Y(n_1174)
);

AOI21xp33_ASAP7_75t_L g1175 ( 
.A1(n_1103),
.A2(n_1008),
.B(n_987),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_993),
.B(n_1011),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_981),
.B(n_1064),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1102),
.A2(n_988),
.B1(n_989),
.B2(n_1024),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1157),
.A2(n_1158),
.B(n_1029),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_981),
.B(n_1067),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1030),
.A2(n_1019),
.B(n_1060),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1069),
.B(n_999),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1043),
.A2(n_1085),
.B(n_1076),
.Y(n_1183)
);

O2A1O1Ixp5_ASAP7_75t_L g1184 ( 
.A1(n_1123),
.A2(n_982),
.B(n_1085),
.C(n_1099),
.Y(n_1184)
);

OA22x2_ASAP7_75t_L g1185 ( 
.A1(n_1127),
.A2(n_1009),
.B1(n_1021),
.B2(n_1066),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_999),
.B(n_1104),
.Y(n_1186)
);

O2A1O1Ixp5_ASAP7_75t_L g1187 ( 
.A1(n_1162),
.A2(n_1055),
.B(n_1061),
.C(n_1096),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_980),
.A2(n_992),
.B(n_983),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_SL g1189 ( 
.A1(n_1138),
.A2(n_1016),
.B(n_1033),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1106),
.A2(n_1155),
.B1(n_1102),
.B2(n_1147),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_L g1191 ( 
.A(n_1103),
.B(n_1117),
.C(n_1078),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1070),
.A2(n_1015),
.B(n_1012),
.Y(n_1192)
);

OAI21xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1148),
.A2(n_1110),
.B(n_1149),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1010),
.Y(n_1194)
);

OAI22x1_ASAP7_75t_L g1195 ( 
.A1(n_1054),
.A2(n_1109),
.B1(n_1143),
.B2(n_1125),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1071),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1095),
.A2(n_1048),
.B(n_1032),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_985),
.A2(n_1025),
.B(n_1047),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1025),
.A2(n_1047),
.B(n_990),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1041),
.A2(n_1056),
.A3(n_1026),
.B(n_1075),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1081),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1071),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1081),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1013),
.A2(n_1078),
.B1(n_1164),
.B2(n_1124),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1041),
.A2(n_1040),
.B(n_1115),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1058),
.A2(n_1059),
.B(n_1118),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1108),
.B(n_1094),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1027),
.A2(n_1151),
.B(n_995),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1014),
.A2(n_1000),
.B(n_1007),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1137),
.A2(n_1145),
.B(n_1141),
.Y(n_1210)
);

O2A1O1Ixp5_ASAP7_75t_L g1211 ( 
.A1(n_1056),
.A2(n_1062),
.B(n_1037),
.C(n_1051),
.Y(n_1211)
);

OAI22x1_ASAP7_75t_L g1212 ( 
.A1(n_1109),
.A2(n_1125),
.B1(n_1098),
.B2(n_1039),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1164),
.A2(n_1017),
.B1(n_1020),
.B2(n_1146),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1108),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1031),
.B(n_1045),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1023),
.B(n_1154),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1049),
.B(n_1088),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1042),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1002),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1101),
.B(n_1017),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1038),
.A2(n_1114),
.B(n_1075),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1091),
.Y(n_1222)
);

NAND3xp33_ASAP7_75t_SL g1223 ( 
.A(n_1142),
.B(n_1068),
.C(n_1050),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1089),
.B(n_1134),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1138),
.A2(n_1107),
.B(n_1161),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1149),
.A2(n_1093),
.B(n_1122),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1131),
.A2(n_1111),
.B(n_1113),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1136),
.B(n_1100),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1050),
.B(n_1112),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1079),
.B(n_1165),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1142),
.A2(n_1084),
.B(n_1090),
.C(n_1073),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_1035),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1132),
.A2(n_1140),
.B(n_1003),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_997),
.A2(n_1003),
.B(n_1018),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1035),
.B(n_1146),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_L g1236 ( 
.A1(n_1139),
.A2(n_997),
.B(n_1018),
.C(n_1121),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1156),
.A2(n_1163),
.B(n_1128),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1005),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1023),
.A2(n_1073),
.B(n_1080),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1146),
.B(n_1116),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1034),
.A2(n_1121),
.B(n_1074),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1106),
.B(n_1120),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1120),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1023),
.A2(n_1072),
.B(n_1063),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1034),
.A2(n_1074),
.B(n_1044),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1044),
.A2(n_1046),
.B(n_1065),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1023),
.B(n_1163),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1086),
.A2(n_1087),
.B(n_1092),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1126),
.A2(n_1077),
.B(n_1129),
.Y(n_1250)
);

AND2x2_ASAP7_75t_SL g1251 ( 
.A(n_1130),
.B(n_1133),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1152),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1152),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1130),
.A2(n_1133),
.B1(n_1152),
.B2(n_1119),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1119),
.A2(n_1135),
.B(n_1133),
.Y(n_1255)
);

CKINVDCx6p67_ASAP7_75t_R g1256 ( 
.A(n_1130),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_R g1257 ( 
.A(n_1130),
.B(n_1133),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1152),
.A2(n_830),
.B1(n_829),
.B2(n_984),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1135),
.B(n_984),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_993),
.A2(n_987),
.B(n_994),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_984),
.A2(n_1006),
.B(n_829),
.C(n_830),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_984),
.B(n_829),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_993),
.A2(n_987),
.B(n_994),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1081),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1006),
.A2(n_830),
.B(n_829),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1022),
.A2(n_1041),
.A3(n_1056),
.B(n_1150),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1006),
.A2(n_830),
.B(n_829),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1160),
.B(n_770),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_996),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1160),
.B(n_770),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_991),
.A2(n_1036),
.B(n_1028),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_984),
.B(n_829),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_984),
.B(n_829),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_986),
.B(n_935),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1006),
.A2(n_1052),
.B(n_830),
.Y(n_1275)
);

NAND2x1_ASAP7_75t_L g1276 ( 
.A(n_997),
.B(n_1003),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_996),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_984),
.A2(n_830),
.B1(n_829),
.B2(n_1006),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1022),
.A2(n_1041),
.A3(n_1056),
.B(n_1150),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1006),
.B(n_984),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1160),
.B(n_770),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_984),
.B(n_829),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_984),
.B(n_829),
.Y(n_1283)
);

OA22x2_ASAP7_75t_L g1284 ( 
.A1(n_1159),
.A2(n_776),
.B1(n_1160),
.B2(n_874),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_984),
.B(n_829),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_984),
.B(n_829),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_993),
.A2(n_987),
.B(n_994),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1094),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_984),
.B(n_829),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_984),
.B(n_829),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1160),
.B(n_770),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_984),
.B(n_829),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1042),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1004),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_993),
.A2(n_987),
.B(n_994),
.Y(n_1295)
);

AO21x1_ASAP7_75t_L g1296 ( 
.A1(n_1006),
.A2(n_1052),
.B(n_830),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_L g1297 ( 
.A1(n_1105),
.A2(n_1006),
.B(n_1150),
.C(n_1022),
.Y(n_1297)
);

AOI21x1_ASAP7_75t_SL g1298 ( 
.A1(n_1096),
.A2(n_1006),
.B(n_1123),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_984),
.B(n_829),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_984),
.B(n_829),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1004),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_984),
.B(n_829),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1006),
.A2(n_830),
.B(n_829),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1120),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1100),
.B(n_1081),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1006),
.A2(n_830),
.B(n_829),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1006),
.A2(n_829),
.B(n_830),
.C(n_658),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_984),
.A2(n_1006),
.B(n_829),
.C(n_830),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_984),
.B(n_829),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_984),
.B(n_829),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_991),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_991),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_991),
.Y(n_1313)
);

NAND2x1_ASAP7_75t_L g1314 ( 
.A(n_997),
.B(n_1003),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_984),
.B(n_829),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_984),
.B(n_829),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_984),
.B(n_829),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1006),
.A2(n_830),
.B(n_829),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_991),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1006),
.B(n_984),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_984),
.B(n_829),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_993),
.A2(n_987),
.B(n_994),
.Y(n_1322)
);

AOI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1006),
.A2(n_830),
.B(n_829),
.Y(n_1323)
);

OAI22x1_ASAP7_75t_L g1324 ( 
.A1(n_1160),
.A2(n_776),
.B1(n_1159),
.B2(n_1127),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1166),
.B(n_1305),
.Y(n_1325)
);

AO21x1_ASAP7_75t_L g1326 ( 
.A1(n_1190),
.A2(n_1278),
.B(n_1175),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1270),
.B(n_1281),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1291),
.B(n_1214),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1274),
.B(n_1240),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1288),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1251),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1170),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1334)
);

CKINVDCx11_ASAP7_75t_R g1335 ( 
.A(n_1293),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1219),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1166),
.B(n_1305),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1315),
.B(n_1272),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1293),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1304),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1207),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1259),
.B(n_1258),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1315),
.B(n_1273),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1269),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1218),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1277),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1251),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1260),
.A2(n_1287),
.B(n_1263),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1170),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1256),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1242),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1170),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1295),
.A2(n_1322),
.B(n_1308),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1219),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_SL g1357 ( 
.A(n_1243),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1286),
.A2(n_1299),
.B1(n_1290),
.B2(n_1300),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1247),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1289),
.B(n_1292),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1166),
.B(n_1305),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1302),
.A2(n_1321),
.B1(n_1316),
.B2(n_1310),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1284),
.B(n_1324),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1274),
.B(n_1264),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1248),
.B(n_1170),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1215),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1284),
.B(n_1171),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_SL g1368 ( 
.A(n_1191),
.B(n_1274),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1217),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1230),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1248),
.B(n_1201),
.Y(n_1371)
);

BUFx10_ASAP7_75t_L g1372 ( 
.A(n_1201),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1264),
.B(n_1248),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1307),
.A2(n_1193),
.B(n_1323),
.C(n_1303),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1309),
.B(n_1317),
.Y(n_1375)
);

OAI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1261),
.A2(n_1308),
.B1(n_1318),
.B2(n_1306),
.C(n_1267),
.Y(n_1376)
);

BUFx2_ASAP7_75t_SL g1377 ( 
.A(n_1201),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1261),
.A2(n_1265),
.B(n_1169),
.C(n_1320),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1238),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1178),
.A2(n_1320),
.B1(n_1280),
.B2(n_1223),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1201),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1185),
.A2(n_1167),
.B1(n_1213),
.B2(n_1212),
.Y(n_1382)
);

OR2x6_ASAP7_75t_L g1383 ( 
.A(n_1235),
.B(n_1185),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1186),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1195),
.B(n_1224),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1176),
.B(n_1280),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1203),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1177),
.B(n_1180),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1204),
.A2(n_1213),
.B1(n_1182),
.B2(n_1231),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1203),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1225),
.A2(n_1222),
.B(n_1184),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1203),
.B(n_1252),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1220),
.B(n_1204),
.Y(n_1394)
);

OAI21xp33_ASAP7_75t_L g1395 ( 
.A1(n_1231),
.A2(n_1221),
.B(n_1188),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1297),
.A2(n_1173),
.B(n_1184),
.C(n_1192),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1203),
.B(n_1252),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1253),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1275),
.B(n_1296),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1226),
.B(n_1253),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1276),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1257),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1255),
.A2(n_1205),
.B1(n_1232),
.B2(n_1254),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1241),
.A2(n_1216),
.B1(n_1239),
.B2(n_1314),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1194),
.B(n_1202),
.Y(n_1405)
);

BUFx4_ASAP7_75t_SL g1406 ( 
.A(n_1257),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1266),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1266),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1196),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1202),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1234),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1294),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1301),
.B(n_1279),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1266),
.B(n_1279),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1266),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1297),
.A2(n_1187),
.B(n_1211),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_L g1418 ( 
.A(n_1189),
.B(n_1216),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1200),
.B(n_1279),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1200),
.B(n_1279),
.Y(n_1420)
);

NAND2xp33_ASAP7_75t_SL g1421 ( 
.A(n_1209),
.B(n_1298),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1200),
.B(n_1174),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1249),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1250),
.B(n_1244),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1198),
.A2(n_1199),
.B1(n_1210),
.B2(n_1227),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1200),
.B(n_1179),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1187),
.B(n_1236),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1233),
.A2(n_1211),
.B(n_1206),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1181),
.B(n_1208),
.Y(n_1429)
);

OAI21xp33_ASAP7_75t_L g1430 ( 
.A1(n_1298),
.A2(n_1237),
.B(n_1183),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1236),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1319),
.A2(n_1172),
.B(n_1311),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1197),
.A2(n_1271),
.B(n_1312),
.C(n_1313),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1271),
.B(n_1262),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1168),
.B(n_751),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1261),
.A2(n_1308),
.B(n_1297),
.Y(n_1436)
);

O2A1O1Ixp5_ASAP7_75t_L g1437 ( 
.A1(n_1297),
.A2(n_830),
.B(n_829),
.C(n_1006),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1166),
.B(n_1305),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1214),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1269),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1214),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1269),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1293),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1278),
.A2(n_1263),
.B(n_1260),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1446)
);

CKINVDCx8_ASAP7_75t_R g1447 ( 
.A(n_1214),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1166),
.B(n_1305),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1262),
.A2(n_1315),
.B1(n_1285),
.B2(n_1272),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1293),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1288),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1288),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1269),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1259),
.B(n_1258),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1256),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1269),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1247),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1278),
.A2(n_829),
.B(n_830),
.C(n_1261),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1278),
.A2(n_1263),
.B(n_1260),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1463)
);

OR2x6_ASAP7_75t_SL g1464 ( 
.A(n_1191),
.B(n_703),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1251),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1262),
.A2(n_1285),
.B1(n_1315),
.B2(n_984),
.Y(n_1467)
);

CKINVDCx16_ASAP7_75t_R g1468 ( 
.A(n_1293),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1293),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1284),
.A2(n_1159),
.B1(n_776),
.B2(n_1160),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1219),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1269),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1219),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1293),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1269),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1271),
.A2(n_1311),
.B(n_1172),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1166),
.B(n_1305),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1278),
.A2(n_829),
.B(n_830),
.C(n_1261),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1218),
.B(n_937),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1261),
.A2(n_1308),
.B(n_1297),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1284),
.A2(n_1159),
.B1(n_776),
.B2(n_1160),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1168),
.B(n_1268),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1278),
.A2(n_1263),
.B(n_1260),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1269),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1251),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1331),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1368),
.A2(n_1363),
.B1(n_1337),
.B2(n_1389),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1453),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1335),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1415),
.B(n_1367),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1334),
.B(n_1446),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1325),
.B(n_1338),
.Y(n_1494)
);

BUFx2_ASAP7_75t_R g1495 ( 
.A(n_1464),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1346),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1348),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1428),
.A2(n_1432),
.B(n_1391),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1440),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1443),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1467),
.A2(n_1449),
.B1(n_1452),
.B2(n_1334),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1400),
.B(n_1436),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1454),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1449),
.A2(n_1452),
.B1(n_1446),
.B2(n_1455),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1436),
.B(n_1482),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1455),
.B(n_1457),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1482),
.B(n_1416),
.Y(n_1508)
);

BUFx10_ASAP7_75t_L g1509 ( 
.A(n_1444),
.Y(n_1509)
);

AO21x1_ASAP7_75t_L g1510 ( 
.A1(n_1389),
.A2(n_1462),
.B(n_1445),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1457),
.B(n_1339),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1473),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1468),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1477),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1451),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1379),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1431),
.Y(n_1518)
);

AO21x1_ASAP7_75t_SL g1519 ( 
.A1(n_1395),
.A2(n_1417),
.B(n_1434),
.Y(n_1519)
);

OAI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1339),
.A2(n_1344),
.B1(n_1368),
.B2(n_1380),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1402),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1344),
.A2(n_1376),
.B1(n_1358),
.B2(n_1362),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1439),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1382),
.A2(n_1483),
.B1(n_1470),
.B2(n_1383),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1419),
.B(n_1420),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1383),
.A2(n_1394),
.B1(n_1328),
.B2(n_1326),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1366),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1384),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1424),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1394),
.A2(n_1360),
.B1(n_1345),
.B2(n_1388),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1383),
.A2(n_1435),
.B1(n_1385),
.B2(n_1472),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1369),
.Y(n_1532)
);

AOI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1391),
.A2(n_1399),
.B(n_1343),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1442),
.Y(n_1534)
);

NAND2x1p5_ASAP7_75t_L g1535 ( 
.A(n_1364),
.B(n_1373),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1419),
.B(n_1420),
.Y(n_1536)
);

INVx6_ASAP7_75t_L g1537 ( 
.A(n_1332),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1336),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1330),
.B(n_1332),
.Y(n_1539)
);

CKINVDCx6p67_ASAP7_75t_R g1540 ( 
.A(n_1450),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1399),
.A2(n_1426),
.B(n_1422),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1341),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1356),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1358),
.B(n_1362),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1347),
.Y(n_1545)
);

BUFx8_ASAP7_75t_SL g1546 ( 
.A(n_1353),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1471),
.Y(n_1547)
);

CKINVDCx11_ASAP7_75t_R g1548 ( 
.A(n_1447),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1405),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1411),
.Y(n_1550)
);

INVx6_ASAP7_75t_L g1551 ( 
.A(n_1349),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1474),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1325),
.B(n_1338),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1345),
.B(n_1360),
.Y(n_1554)
);

BUFx2_ASAP7_75t_SL g1555 ( 
.A(n_1481),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1441),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1460),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1329),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1409),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1463),
.A2(n_1484),
.B1(n_1327),
.B2(n_1476),
.Y(n_1560)
);

INVx5_ASAP7_75t_L g1561 ( 
.A(n_1330),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1388),
.B(n_1375),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1407),
.B(n_1408),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1374),
.B(n_1361),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1412),
.Y(n_1565)
);

AOI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1350),
.A2(n_1485),
.B(n_1445),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1393),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1376),
.A2(n_1461),
.B1(n_1480),
.B2(n_1386),
.Y(n_1568)
);

AOI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1462),
.A2(n_1485),
.B(n_1355),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1364),
.B(n_1373),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1426),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1410),
.Y(n_1572)
);

CKINVDCx11_ASAP7_75t_R g1573 ( 
.A(n_1469),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1465),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1422),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1386),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1411),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1475),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1460),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1456),
.A2(n_1487),
.B1(n_1349),
.B2(n_1466),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1361),
.B(n_1479),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1349),
.Y(n_1582)
);

CKINVDCx6p67_ASAP7_75t_R g1583 ( 
.A(n_1387),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1359),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1411),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1378),
.A2(n_1423),
.B1(n_1355),
.B2(n_1396),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1424),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1414),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1417),
.A2(n_1430),
.B(n_1433),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1414),
.Y(n_1590)
);

BUFx2_ASAP7_75t_R g1591 ( 
.A(n_1370),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1392),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1466),
.A2(n_1487),
.B1(n_1403),
.B2(n_1438),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1403),
.A2(n_1487),
.B1(n_1466),
.B2(n_1479),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1365),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1365),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1438),
.B(n_1448),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1371),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1351),
.Y(n_1599)
);

AOI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1427),
.A2(n_1418),
.B(n_1434),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1340),
.A2(n_1397),
.B1(n_1357),
.B2(n_1421),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1397),
.Y(n_1602)
);

BUFx12f_ASAP7_75t_L g1603 ( 
.A(n_1372),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1390),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1351),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1478),
.Y(n_1606)
);

BUFx2_ASAP7_75t_SL g1607 ( 
.A(n_1352),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1437),
.A2(n_1425),
.B(n_1429),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1398),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1398),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1352),
.A2(n_1458),
.B1(n_1406),
.B2(n_1377),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1351),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1429),
.A2(n_1404),
.B(n_1381),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1372),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1354),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1354),
.B(n_1333),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1354),
.B(n_1333),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1458),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1401),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1401),
.A2(n_1428),
.B(n_1432),
.Y(n_1620)
);

BUFx12f_ASAP7_75t_L g1621 ( 
.A(n_1401),
.Y(n_1621)
);

BUFx8_ASAP7_75t_L g1622 ( 
.A(n_1331),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1351),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1346),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1337),
.B(n_703),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1332),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1382),
.A2(n_1284),
.B1(n_1159),
.B2(n_1185),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1346),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1346),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1431),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1467),
.A2(n_830),
.B1(n_829),
.B2(n_1334),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1413),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1431),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1431),
.Y(n_1634)
);

BUFx8_ASAP7_75t_L g1635 ( 
.A(n_1331),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1346),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1467),
.B(n_1461),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1342),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1325),
.B(n_1338),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1342),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1431),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1346),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1346),
.Y(n_1643)
);

BUFx10_ASAP7_75t_L g1644 ( 
.A(n_1444),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1346),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1467),
.A2(n_1337),
.B1(n_1262),
.B2(n_1315),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1346),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1502),
.B(n_1506),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1502),
.B(n_1506),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1603),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1529),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1498),
.A2(n_1510),
.B(n_1569),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1525),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1525),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1498),
.A2(n_1566),
.B(n_1620),
.Y(n_1655)
);

AOI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1566),
.A2(n_1533),
.B(n_1569),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1536),
.Y(n_1657)
);

OA21x2_ASAP7_75t_L g1658 ( 
.A1(n_1510),
.A2(n_1608),
.B(n_1620),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1536),
.B(n_1508),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1575),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1563),
.B(n_1529),
.Y(n_1661)
);

OA21x2_ASAP7_75t_L g1662 ( 
.A1(n_1606),
.A2(n_1544),
.B(n_1600),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1492),
.B(n_1519),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1613),
.A2(n_1600),
.B(n_1606),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1587),
.B(n_1588),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1523),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1588),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1575),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1571),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1590),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1571),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1541),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1586),
.A2(n_1530),
.B(n_1541),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1613),
.A2(n_1577),
.B(n_1550),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1548),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1554),
.B(n_1505),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1541),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1564),
.B(n_1496),
.Y(n_1679)
);

INVx2_ASAP7_75t_SL g1680 ( 
.A(n_1521),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1517),
.A2(n_1520),
.B(n_1565),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1550),
.A2(n_1585),
.B(n_1577),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1564),
.B(n_1497),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1550),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1528),
.B(n_1640),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1527),
.A2(n_1532),
.B(n_1647),
.Y(n_1686)
);

CKINVDCx14_ASAP7_75t_R g1687 ( 
.A(n_1491),
.Y(n_1687)
);

AO21x2_ASAP7_75t_L g1688 ( 
.A1(n_1499),
.A2(n_1503),
.B(n_1500),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1577),
.A2(n_1585),
.B(n_1589),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1534),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1521),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1637),
.A2(n_1646),
.B(n_1522),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1504),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1512),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1514),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1489),
.A2(n_1625),
.B1(n_1501),
.B2(n_1637),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1558),
.Y(n_1697)
);

AOI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1568),
.A2(n_1630),
.B(n_1641),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1526),
.A2(n_1576),
.B(n_1632),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1589),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1589),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1511),
.B(n_1493),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1515),
.B(n_1624),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1609),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1507),
.B(n_1578),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1518),
.A2(n_1605),
.B(n_1599),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1628),
.B(n_1629),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1636),
.B(n_1642),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1643),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1645),
.Y(n_1710)
);

OA21x2_ASAP7_75t_L g1711 ( 
.A1(n_1531),
.A2(n_1538),
.B(n_1543),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1584),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1518),
.A2(n_1599),
.B(n_1605),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1623),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1547),
.Y(n_1715)
);

AND2x6_ASAP7_75t_L g1716 ( 
.A(n_1518),
.B(n_1582),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1552),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1567),
.B(n_1549),
.Y(n_1718)
);

AO31x2_ASAP7_75t_L g1719 ( 
.A1(n_1549),
.A2(n_1572),
.A3(n_1559),
.B(n_1602),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1599),
.A2(n_1605),
.B(n_1612),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1556),
.B(n_1574),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1610),
.Y(n_1722)
);

AOI222xp33_ASAP7_75t_L g1723 ( 
.A1(n_1524),
.A2(n_1627),
.B1(n_1631),
.B2(n_1560),
.C1(n_1562),
.C2(n_1516),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1619),
.Y(n_1724)
);

AOI21xp33_ASAP7_75t_L g1725 ( 
.A1(n_1630),
.A2(n_1633),
.B(n_1641),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1595),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1604),
.Y(n_1727)
);

AO21x1_ASAP7_75t_SL g1728 ( 
.A1(n_1601),
.A2(n_1593),
.B(n_1580),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1596),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1598),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1488),
.A2(n_1490),
.B(n_1611),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1592),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1612),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1634),
.B(n_1618),
.Y(n_1734)
);

AOI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1634),
.A2(n_1618),
.B(n_1617),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1616),
.B(n_1617),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1546),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1561),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1539),
.B(n_1616),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1603),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1581),
.B(n_1553),
.Y(n_1741)
);

INVxp67_ASAP7_75t_SL g1742 ( 
.A(n_1535),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1597),
.B(n_1579),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1539),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1615),
.Y(n_1745)
);

AO21x2_ASAP7_75t_L g1746 ( 
.A1(n_1494),
.A2(n_1639),
.B(n_1553),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1622),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1570),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1539),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1557),
.B(n_1635),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1582),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1594),
.B(n_1513),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1622),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1546),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1622),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1548),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1582),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1626),
.Y(n_1758)
);

INVxp67_ASAP7_75t_SL g1759 ( 
.A(n_1626),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1677),
.B(n_1635),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1696),
.A2(n_1555),
.B1(n_1607),
.B2(n_1557),
.C(n_1495),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1648),
.B(n_1540),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1659),
.B(n_1540),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1648),
.B(n_1623),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1716),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1649),
.B(n_1635),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1689),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1716),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1659),
.B(n_1513),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1663),
.B(n_1578),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1655),
.A2(n_1614),
.B(n_1537),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1692),
.A2(n_1545),
.B1(n_1551),
.B2(n_1537),
.C(n_1614),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1688),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1663),
.B(n_1583),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1702),
.B(n_1583),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1688),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1728),
.A2(n_1711),
.B1(n_1673),
.B2(n_1699),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1688),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1686),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1679),
.B(n_1644),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1675),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1685),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1683),
.B(n_1509),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1683),
.B(n_1509),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1709),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1661),
.B(n_1626),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1709),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1710),
.Y(n_1788)
);

NOR2x1_ASAP7_75t_SL g1789 ( 
.A(n_1746),
.B(n_1621),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1665),
.B(n_1545),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1665),
.B(n_1491),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1697),
.B(n_1573),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1710),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1752),
.A2(n_1621),
.B1(n_1551),
.B2(n_1537),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1651),
.B(n_1573),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1698),
.A2(n_1542),
.B(n_1591),
.Y(n_1796)
);

NOR2x1_ASAP7_75t_SL g1797 ( 
.A(n_1746),
.B(n_1551),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1653),
.B(n_1542),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1651),
.B(n_1654),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_1722),
.B(n_1723),
.C(n_1733),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1657),
.B(n_1736),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1736),
.B(n_1703),
.Y(n_1802)
);

NAND2x1_ASAP7_75t_L g1803 ( 
.A(n_1716),
.B(n_1662),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1712),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1728),
.A2(n_1711),
.B1(n_1673),
.B2(n_1699),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1673),
.B(n_1727),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1684),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1682),
.B(n_1674),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1707),
.B(n_1708),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1708),
.B(n_1700),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1727),
.B(n_1718),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1701),
.B(n_1662),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1662),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1698),
.B(n_1705),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1718),
.B(n_1732),
.Y(n_1815)
);

BUFx2_ASAP7_75t_SL g1816 ( 
.A(n_1716),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1701),
.B(n_1662),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1684),
.B(n_1722),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1693),
.B(n_1694),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1666),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1734),
.B(n_1695),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1682),
.B(n_1674),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1717),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1800),
.A2(n_1761),
.B1(n_1805),
.B2(n_1777),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1782),
.B(n_1690),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_L g1826 ( 
.A1(n_1814),
.A2(n_1731),
.B1(n_1725),
.B2(n_1743),
.C(n_1734),
.Y(n_1826)
);

NAND4xp25_ASAP7_75t_L g1827 ( 
.A(n_1781),
.B(n_1676),
.C(n_1756),
.D(n_1733),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1802),
.B(n_1680),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1806),
.B(n_1704),
.C(n_1745),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1760),
.A2(n_1691),
.B1(n_1680),
.B2(n_1755),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1794),
.A2(n_1746),
.B1(n_1748),
.B2(n_1742),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1804),
.B(n_1721),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_L g1833 ( 
.A(n_1806),
.B(n_1704),
.C(n_1658),
.Y(n_1833)
);

NOR3xp33_ASAP7_75t_SL g1834 ( 
.A(n_1796),
.B(n_1754),
.C(n_1737),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1812),
.A2(n_1681),
.B1(n_1699),
.B2(n_1743),
.Y(n_1835)
);

NAND4xp25_ASAP7_75t_L g1836 ( 
.A(n_1798),
.B(n_1650),
.C(n_1740),
.D(n_1750),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_L g1837 ( 
.A(n_1812),
.B(n_1658),
.C(n_1678),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1772),
.A2(n_1687),
.B(n_1747),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1765),
.B(n_1735),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1785),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1817),
.A2(n_1789),
.B1(n_1797),
.B2(n_1816),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_SL g1842 ( 
.A1(n_1795),
.A2(n_1753),
.B(n_1735),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1795),
.A2(n_1774),
.B(n_1791),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1809),
.B(n_1741),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1801),
.B(n_1719),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1801),
.B(n_1719),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1763),
.A2(n_1717),
.B1(n_1724),
.B2(n_1715),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1791),
.B(n_1739),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1762),
.A2(n_1716),
.B1(n_1744),
.B2(n_1749),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1763),
.A2(n_1775),
.B1(n_1769),
.B2(n_1766),
.Y(n_1850)
);

NAND3xp33_ASAP7_75t_L g1851 ( 
.A(n_1773),
.B(n_1658),
.C(n_1672),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1791),
.B(n_1739),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_L g1853 ( 
.A(n_1773),
.B(n_1658),
.C(n_1758),
.Y(n_1853)
);

OAI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1818),
.A2(n_1757),
.B(n_1656),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1769),
.A2(n_1650),
.B1(n_1740),
.B2(n_1714),
.Y(n_1855)
);

NOR3xp33_ASAP7_75t_SL g1856 ( 
.A(n_1792),
.B(n_1759),
.C(n_1738),
.Y(n_1856)
);

OAI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1818),
.A2(n_1656),
.B(n_1706),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1799),
.B(n_1667),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1820),
.B(n_1667),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1780),
.B(n_1706),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1810),
.B(n_1652),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1803),
.A2(n_1726),
.B1(n_1730),
.B2(n_1729),
.C(n_1751),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1785),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1821),
.B(n_1670),
.Y(n_1864)
);

OA21x2_ASAP7_75t_L g1865 ( 
.A1(n_1776),
.A2(n_1655),
.B(n_1664),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1776),
.B(n_1652),
.C(n_1730),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1821),
.B(n_1713),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1819),
.B(n_1713),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1823),
.A2(n_1668),
.B1(n_1660),
.B2(n_1669),
.C(n_1671),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1813),
.B(n_1720),
.C(n_1751),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1819),
.B(n_1726),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1787),
.Y(n_1872)
);

OA21x2_ASAP7_75t_L g1873 ( 
.A1(n_1778),
.A2(n_1664),
.B(n_1720),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1861),
.B(n_1764),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1840),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1839),
.B(n_1768),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1863),
.Y(n_1877)
);

INVx2_ASAP7_75t_SL g1878 ( 
.A(n_1868),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1844),
.B(n_1807),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1873),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1873),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1828),
.B(n_1807),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1872),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1856),
.B(n_1790),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1873),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1839),
.B(n_1768),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1851),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1845),
.B(n_1811),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1846),
.B(n_1867),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1837),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1860),
.B(n_1808),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1860),
.B(n_1808),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1865),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1832),
.B(n_1815),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1866),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1824),
.A2(n_1711),
.B1(n_1784),
.B2(n_1783),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1833),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1865),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1848),
.B(n_1822),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1852),
.B(n_1822),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1871),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1841),
.B(n_1771),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1858),
.B(n_1771),
.Y(n_1903)
);

NAND2x1p5_ASAP7_75t_L g1904 ( 
.A(n_1831),
.B(n_1803),
.Y(n_1904)
);

INVxp33_ASAP7_75t_L g1905 ( 
.A(n_1856),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1842),
.B(n_1787),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1865),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1854),
.B(n_1788),
.Y(n_1908)
);

OR2x6_ASAP7_75t_SL g1909 ( 
.A(n_1850),
.B(n_1786),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1853),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1870),
.B(n_1771),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1857),
.B(n_1771),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1829),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1864),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1862),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1847),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1876),
.Y(n_1917)
);

NAND2x1p5_ASAP7_75t_L g1918 ( 
.A(n_1884),
.B(n_1765),
.Y(n_1918)
);

NAND3xp33_ASAP7_75t_SL g1919 ( 
.A(n_1905),
.B(n_1824),
.C(n_1826),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1887),
.B(n_1788),
.Y(n_1920)
);

AOI222xp33_ASAP7_75t_L g1921 ( 
.A1(n_1890),
.A2(n_1835),
.B1(n_1869),
.B2(n_1838),
.C1(n_1779),
.C2(n_1778),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1909),
.B(n_1843),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1875),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1875),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1880),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1905),
.B(n_1827),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1909),
.B(n_1770),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1880),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1888),
.B(n_1825),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1875),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1909),
.B(n_1770),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1913),
.B(n_1836),
.Y(n_1932)
);

OAI21xp33_ASAP7_75t_L g1933 ( 
.A1(n_1897),
.A2(n_1859),
.B(n_1834),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1882),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1890),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1877),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1888),
.B(n_1889),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1877),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1880),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1897),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1877),
.Y(n_1941)
);

CKINVDCx14_ASAP7_75t_R g1942 ( 
.A(n_1879),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1891),
.B(n_1783),
.Y(n_1943)
);

NAND2x1_ASAP7_75t_L g1944 ( 
.A(n_1876),
.B(n_1767),
.Y(n_1944)
);

NOR2x1_ASAP7_75t_L g1945 ( 
.A(n_1887),
.B(n_1830),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1883),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1880),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1897),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1891),
.B(n_1892),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1881),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1883),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1881),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1881),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1876),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1881),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1883),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1901),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1876),
.B(n_1849),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1887),
.B(n_1793),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1882),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1895),
.B(n_1793),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1891),
.B(n_1784),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1889),
.B(n_1823),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1923),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_L g1965 ( 
.A(n_1917),
.B(n_1913),
.Y(n_1965)
);

INVxp33_ASAP7_75t_L g1966 ( 
.A(n_1945),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1923),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1937),
.B(n_1895),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1924),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1924),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1930),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1920),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1945),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1937),
.B(n_1895),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1922),
.B(n_1899),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1925),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1930),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1940),
.B(n_1913),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1936),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1925),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1936),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1938),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1940),
.B(n_1910),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1922),
.B(n_1899),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1948),
.B(n_1935),
.Y(n_1985)
);

A2O1A1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1919),
.A2(n_1896),
.B(n_1916),
.C(n_1910),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1948),
.B(n_1910),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1929),
.B(n_1894),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1938),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1926),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1941),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1949),
.B(n_1910),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1932),
.B(n_1914),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1929),
.B(n_1906),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1941),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1963),
.B(n_1906),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1927),
.B(n_1899),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1946),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1963),
.B(n_1961),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1927),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1931),
.B(n_1900),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1931),
.B(n_1900),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1925),
.Y(n_2003)
);

NAND3xp33_ASAP7_75t_L g2004 ( 
.A(n_1921),
.B(n_1896),
.C(n_1911),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1942),
.Y(n_2005)
);

NAND2x2_ASAP7_75t_L g2006 ( 
.A(n_1934),
.B(n_1878),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1946),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1949),
.B(n_1900),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1961),
.B(n_1914),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1951),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1934),
.B(n_1874),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1944),
.Y(n_2012)
);

INVxp67_ASAP7_75t_SL g2013 ( 
.A(n_1920),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1960),
.B(n_1874),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1959),
.B(n_1914),
.Y(n_2015)
);

NOR2x1p5_ASAP7_75t_SL g2016 ( 
.A(n_1928),
.B(n_1885),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1959),
.B(n_1901),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1964),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1973),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1967),
.Y(n_2020)
);

INVxp67_ASAP7_75t_L g2021 ( 
.A(n_2005),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1966),
.B(n_1919),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1975),
.B(n_1984),
.Y(n_2023)
);

INVx3_ASAP7_75t_SL g2024 ( 
.A(n_1987),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1985),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1969),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1966),
.B(n_1921),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1975),
.B(n_1917),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1970),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1992),
.Y(n_2030)
);

CKINVDCx16_ASAP7_75t_R g2031 ( 
.A(n_1984),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1990),
.B(n_1933),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2008),
.B(n_1917),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1993),
.B(n_1960),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2008),
.B(n_1917),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_L g2036 ( 
.A(n_1987),
.B(n_1954),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1992),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1968),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1971),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1977),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1979),
.Y(n_2041)
);

INVxp67_ASAP7_75t_SL g2042 ( 
.A(n_1983),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1988),
.B(n_1957),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1981),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1968),
.B(n_1957),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1982),
.Y(n_2046)
);

AO22x1_ASAP7_75t_L g2047 ( 
.A1(n_1978),
.A2(n_1916),
.B1(n_1958),
.B2(n_1902),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1974),
.B(n_1933),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1992),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1989),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1991),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1997),
.B(n_1954),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1995),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1965),
.B(n_1918),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_1974),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1998),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_2007),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2057),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2031),
.B(n_2000),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2057),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2018),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2024),
.B(n_2055),
.Y(n_2062)
);

AOI31xp33_ASAP7_75t_L g2063 ( 
.A1(n_2032),
.A2(n_2021),
.A3(n_2048),
.B(n_2022),
.Y(n_2063)
);

AOI32xp33_ASAP7_75t_L g2064 ( 
.A1(n_2027),
.A2(n_1912),
.A3(n_1911),
.B1(n_1902),
.B2(n_2004),
.Y(n_2064)
);

AOI21xp33_ASAP7_75t_L g2065 ( 
.A1(n_2019),
.A2(n_1986),
.B(n_2013),
.Y(n_2065)
);

OAI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2024),
.A2(n_1986),
.B1(n_2042),
.B2(n_2019),
.C(n_1904),
.Y(n_2066)
);

O2A1O1Ixp5_ASAP7_75t_SL g2067 ( 
.A1(n_2038),
.A2(n_2025),
.B(n_2020),
.C(n_2018),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_2030),
.B(n_1997),
.Y(n_2068)
);

AOI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_2047),
.A2(n_1915),
.B1(n_1916),
.B2(n_1902),
.Y(n_2069)
);

AOI332xp33_ASAP7_75t_L g2070 ( 
.A1(n_2020),
.A2(n_2010),
.A3(n_2009),
.B1(n_2015),
.B2(n_1951),
.B3(n_1956),
.C1(n_1939),
.C2(n_1950),
.Y(n_2070)
);

INVx1_ASAP7_75t_SL g2071 ( 
.A(n_2024),
.Y(n_2071)
);

OAI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_2030),
.A2(n_1904),
.B1(n_1915),
.B2(n_2006),
.Y(n_2072)
);

AOI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2047),
.A2(n_1912),
.B1(n_1911),
.B2(n_1885),
.C(n_1972),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2026),
.Y(n_2074)
);

OAI21xp5_ASAP7_75t_SL g2075 ( 
.A1(n_2023),
.A2(n_1918),
.B(n_1904),
.Y(n_2075)
);

OR2x6_ASAP7_75t_L g2076 ( 
.A(n_2037),
.B(n_2049),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_2054),
.A2(n_1994),
.B(n_1915),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2023),
.A2(n_2006),
.B1(n_1918),
.B2(n_1904),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2037),
.A2(n_1915),
.B1(n_1912),
.B2(n_1904),
.Y(n_2079)
);

AOI32xp33_ASAP7_75t_L g2080 ( 
.A1(n_2036),
.A2(n_1994),
.A3(n_1996),
.B1(n_1958),
.B2(n_2001),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_2049),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2026),
.Y(n_2082)
);

AOI222xp33_ASAP7_75t_L g2083 ( 
.A1(n_2029),
.A2(n_2016),
.B1(n_1976),
.B2(n_1980),
.C1(n_2003),
.C2(n_1835),
.Y(n_2083)
);

OA21x2_ASAP7_75t_L g2084 ( 
.A1(n_2029),
.A2(n_1980),
.B(n_1976),
.Y(n_2084)
);

INVxp67_ASAP7_75t_L g2085 ( 
.A(n_2046),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2034),
.A2(n_2028),
.B1(n_2003),
.B2(n_1958),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2062),
.B(n_2043),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2071),
.B(n_2043),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_2063),
.B(n_2065),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2059),
.B(n_2045),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2081),
.B(n_2045),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2061),
.Y(n_2092)
);

INVxp67_ASAP7_75t_L g2093 ( 
.A(n_2076),
.Y(n_2093)
);

NOR2x1_ASAP7_75t_L g2094 ( 
.A(n_2058),
.B(n_2039),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2074),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2084),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_2060),
.B(n_2039),
.Y(n_2097)
);

INVxp67_ASAP7_75t_SL g2098 ( 
.A(n_2084),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2068),
.B(n_2040),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2083),
.A2(n_1928),
.B1(n_1939),
.B2(n_1947),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2068),
.B(n_2028),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_2076),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_2085),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2069),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2082),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_2086),
.Y(n_2106)
);

NAND2x1_ASAP7_75t_L g2107 ( 
.A(n_2078),
.B(n_2012),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2077),
.B(n_1996),
.Y(n_2108)
);

OAI21xp33_ASAP7_75t_SL g2109 ( 
.A1(n_2098),
.A2(n_2067),
.B(n_2080),
.Y(n_2109)
);

NAND4xp25_ASAP7_75t_L g2110 ( 
.A(n_2089),
.B(n_2064),
.C(n_2066),
.D(n_2073),
.Y(n_2110)
);

NAND4xp25_ASAP7_75t_L g2111 ( 
.A(n_2089),
.B(n_2075),
.C(n_2052),
.D(n_2033),
.Y(n_2111)
);

AOI211xp5_ASAP7_75t_L g2112 ( 
.A1(n_2108),
.A2(n_2072),
.B(n_2070),
.C(n_2040),
.Y(n_2112)
);

AOI211xp5_ASAP7_75t_SL g2113 ( 
.A1(n_2103),
.A2(n_2012),
.B(n_2041),
.C(n_2056),
.Y(n_2113)
);

AOI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2104),
.A2(n_2100),
.B1(n_2096),
.B2(n_2106),
.C(n_2093),
.Y(n_2114)
);

OAI322xp33_ASAP7_75t_L g2115 ( 
.A1(n_2104),
.A2(n_2041),
.A3(n_2044),
.B1(n_2050),
.B2(n_2051),
.C1(n_2056),
.C2(n_2053),
.Y(n_2115)
);

OAI211xp5_ASAP7_75t_L g2116 ( 
.A1(n_2094),
.A2(n_2079),
.B(n_2053),
.C(n_2051),
.Y(n_2116)
);

AOI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2100),
.A2(n_1953),
.B1(n_1928),
.B2(n_1955),
.C(n_1952),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2096),
.A2(n_2050),
.B(n_2044),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_2102),
.B(n_1999),
.Y(n_2119)
);

AOI222xp33_ASAP7_75t_L g2120 ( 
.A1(n_2097),
.A2(n_1955),
.B1(n_1939),
.B2(n_1947),
.C1(n_1953),
.C2(n_1952),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_2090),
.A2(n_2097),
.B(n_2088),
.Y(n_2121)
);

OAI211xp5_ASAP7_75t_L g2122 ( 
.A1(n_2099),
.A2(n_2052),
.B(n_2012),
.C(n_2033),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_2109),
.A2(n_2091),
.B(n_2105),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_2121),
.B(n_2087),
.Y(n_2124)
);

NAND4xp25_ASAP7_75t_L g2125 ( 
.A(n_2113),
.B(n_2101),
.C(n_2095),
.D(n_2092),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_2119),
.B(n_2101),
.Y(n_2126)
);

NAND3xp33_ASAP7_75t_L g2127 ( 
.A(n_2114),
.B(n_2105),
.C(n_2107),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_2116),
.A2(n_2017),
.B(n_2035),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2118),
.Y(n_2129)
);

NAND3xp33_ASAP7_75t_L g2130 ( 
.A(n_2112),
.B(n_2035),
.C(n_1999),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2110),
.B(n_2111),
.Y(n_2131)
);

NAND3xp33_ASAP7_75t_SL g2132 ( 
.A(n_2122),
.B(n_1944),
.C(n_2001),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2115),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2126),
.Y(n_2134)
);

AND4x1_ASAP7_75t_L g2135 ( 
.A(n_2127),
.B(n_1834),
.C(n_2120),
.D(n_2117),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_2124),
.B(n_1954),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_SL g2137 ( 
.A(n_2125),
.B(n_2011),
.Y(n_2137)
);

OAI211xp5_ASAP7_75t_L g2138 ( 
.A1(n_2123),
.A2(n_1954),
.B(n_2002),
.C(n_2011),
.Y(n_2138)
);

NAND3xp33_ASAP7_75t_L g2139 ( 
.A(n_2133),
.B(n_1950),
.C(n_1947),
.Y(n_2139)
);

NAND4xp25_ASAP7_75t_SL g2140 ( 
.A(n_2130),
.B(n_2002),
.C(n_2014),
.D(n_1962),
.Y(n_2140)
);

OAI211xp5_ASAP7_75t_SL g2141 ( 
.A1(n_2131),
.A2(n_1884),
.B(n_1950),
.C(n_1952),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2134),
.B(n_2129),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2136),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2139),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2137),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2140),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2138),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2135),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2141),
.A2(n_2132),
.B1(n_2128),
.B2(n_1955),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2142),
.Y(n_2150)
);

AO22x1_ASAP7_75t_L g2151 ( 
.A1(n_2142),
.A2(n_2014),
.B1(n_1958),
.B2(n_1886),
.Y(n_2151)
);

NAND3x1_ASAP7_75t_L g2152 ( 
.A(n_2145),
.B(n_1956),
.C(n_1943),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2144),
.B(n_1953),
.Y(n_2153)
);

AND2x2_ASAP7_75t_SL g2154 ( 
.A(n_2147),
.B(n_1876),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2143),
.B(n_1943),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2150),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2152),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2155),
.B(n_2146),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2153),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2156),
.B(n_2154),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2159),
.A2(n_2148),
.B1(n_2157),
.B2(n_2158),
.Y(n_2161)
);

NAND3xp33_ASAP7_75t_L g2162 ( 
.A(n_2161),
.B(n_2158),
.C(n_2149),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2162),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_2162),
.A2(n_2160),
.B1(n_2151),
.B2(n_1907),
.Y(n_2164)
);

OAI21xp33_ASAP7_75t_L g2165 ( 
.A1(n_2163),
.A2(n_1878),
.B(n_1893),
.Y(n_2165)
);

OR2x6_ASAP7_75t_L g2166 ( 
.A(n_2164),
.B(n_1816),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2166),
.Y(n_2167)
);

OAI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2167),
.A2(n_2165),
.B(n_1885),
.Y(n_2168)
);

AOI322xp5_ASAP7_75t_L g2169 ( 
.A1(n_2168),
.A2(n_1885),
.A3(n_1907),
.B1(n_1893),
.B2(n_1898),
.C1(n_1903),
.C2(n_1908),
.Y(n_2169)
);

AOI221xp5_ASAP7_75t_L g2170 ( 
.A1(n_2169),
.A2(n_1893),
.B1(n_1898),
.B2(n_1907),
.C(n_1878),
.Y(n_2170)
);

AOI211xp5_ASAP7_75t_L g2171 ( 
.A1(n_2170),
.A2(n_1855),
.B(n_1898),
.C(n_1893),
.Y(n_2171)
);


endmodule