module fake_jpeg_29968_n_45 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_7),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_20),
.B(n_19),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_31),
.B(n_23),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_13),
.B1(n_12),
.B2(n_19),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_30),
.B1(n_26),
.B2(n_18),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_32),
.C(n_28),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_26),
.C(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_34),
.C(n_18),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_18),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_42),
.C2(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_8),
.Y(n_45)
);


endmodule