module fake_jpeg_18_n_355 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_4),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_71),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_59),
.Y(n_124)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx2_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_63),
.B(n_77),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_69),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_88),
.Y(n_119)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_19),
.B(n_14),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_23),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_91),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_94),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_25),
.Y(n_94)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_SL g96 ( 
.A(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_20),
.B1(n_47),
.B2(n_25),
.Y(n_115)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_97),
.B(n_0),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_44),
.B1(n_22),
.B2(n_42),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_101),
.B1(n_111),
.B2(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_42),
.B1(n_45),
.B2(n_26),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_26),
.B1(n_45),
.B2(n_34),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_92),
.B1(n_76),
.B2(n_84),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_54),
.A2(n_20),
.B1(n_34),
.B2(n_31),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_31),
.B1(n_29),
.B2(n_27),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_113),
.B(n_12),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_29),
.B1(n_27),
.B2(n_47),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_64),
.A2(n_56),
.B1(n_93),
.B2(n_90),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_144),
.B1(n_67),
.B2(n_52),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_73),
.A2(n_30),
.B1(n_0),
.B2(n_6),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_63),
.B(n_4),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_149),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_6),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_157),
.B1(n_98),
.B2(n_143),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_152),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_59),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_156),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_83),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_86),
.B1(n_68),
.B2(n_66),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_81),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_55),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_9),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_102),
.B(n_62),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_162),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_67),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_9),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_9),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_12),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_142),
.C(n_107),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_99),
.A2(n_12),
.B1(n_13),
.B2(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_178),
.Y(n_186)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_128),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_111),
.A2(n_126),
.B1(n_133),
.B2(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_116),
.B1(n_107),
.B2(n_143),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_178),
.C(n_155),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_209),
.B1(n_157),
.B2(n_150),
.Y(n_216)
);

AOI22x1_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_141),
.B1(n_118),
.B2(n_106),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_174),
.B(n_115),
.Y(n_219)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_160),
.B1(n_173),
.B2(n_184),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_116),
.B1(n_108),
.B2(n_132),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_144),
.B1(n_180),
.B2(n_151),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_153),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_215),
.B(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_232),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_171),
.B(n_179),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_223),
.B(n_233),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_164),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_222),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_166),
.B(n_158),
.C(n_162),
.D(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_162),
.C(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_227),
.C(n_202),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_175),
.B1(n_182),
.B2(n_185),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_181),
.C(n_152),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_175),
.B1(n_108),
.B2(n_132),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_172),
.B1(n_167),
.B2(n_180),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_136),
.B1(n_138),
.B2(n_148),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_234),
.B1(n_207),
.B2(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_136),
.B1(n_138),
.B2(n_120),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_177),
.B(n_165),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_120),
.B1(n_118),
.B2(n_154),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_195),
.B1(n_207),
.B2(n_201),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_188),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_242),
.C(n_250),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_255),
.B(n_256),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_186),
.B(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_220),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_245),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_219),
.B1(n_229),
.B2(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_262),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_235),
.B1(n_222),
.B2(n_223),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_231),
.B1(n_234),
.B2(n_218),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_273),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_200),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_272),
.C(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_200),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_186),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_210),
.B1(n_232),
.B2(n_215),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_212),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_263),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_280),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_277),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_245),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_286),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_262),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_287),
.B1(n_289),
.B2(n_257),
.Y(n_302)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_272),
.C(n_258),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_261),
.C(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_290),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_256),
.B(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_291),
.B(n_303),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_265),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_259),
.B(n_238),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_282),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_238),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_197),
.C(n_190),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_295),
.B(n_285),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_203),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_239),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_285),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_292),
.B(n_284),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_321),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_300),
.C(n_293),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_300),
.C(n_304),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_326),
.C(n_309),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_313),
.A2(n_296),
.B1(n_279),
.B2(n_289),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_266),
.C(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_304),
.C(n_286),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_328),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_329),
.B(n_333),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_316),
.B1(n_318),
.B2(n_311),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_331),
.A2(n_251),
.B1(n_193),
.B2(n_204),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_287),
.C(n_247),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_254),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_332),
.A2(n_326),
.B(n_237),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_335),
.A2(n_337),
.B(n_338),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_336),
.A2(n_339),
.B1(n_205),
.B2(n_197),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_327),
.C(n_190),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_208),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_342),
.B(n_343),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_341),
.A2(n_193),
.B(n_205),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_192),
.B(n_199),
.Y(n_345)
);

NAND3xp33_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_346),
.C(n_199),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_192),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_SL g348 ( 
.A1(n_344),
.A2(n_336),
.B(n_104),
.C(n_204),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_SL g350 ( 
.A(n_348),
.B(n_104),
.C(n_125),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

AOI21x1_ASAP7_75t_L g352 ( 
.A1(n_350),
.A2(n_104),
.B(n_347),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_351),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_353),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_125),
.Y(n_355)
);


endmodule