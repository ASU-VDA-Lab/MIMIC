module fake_jpeg_8141_n_170 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_37),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_15),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_32),
.B1(n_21),
.B2(n_27),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_58),
.B1(n_29),
.B2(n_26),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_56),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_30),
.B1(n_21),
.B2(n_32),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_16),
.Y(n_63)
);

AOI31xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_23),
.A3(n_28),
.B(n_30),
.Y(n_84)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_77),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_82),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_35),
.C(n_22),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_89),
.C(n_90),
.Y(n_92)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_89),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_30),
.B1(n_44),
.B2(n_42),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_84),
.B(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_23),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_62),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_103),
.CI(n_28),
.CON(n_123),
.SN(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_101),
.Y(n_118)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_87),
.Y(n_101)
);

XOR2x2_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_88),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_53),
.C(n_56),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_113),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_119),
.C(n_92),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_77),
.B1(n_70),
.B2(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_120),
.B1(n_95),
.B2(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_115),
.B1(n_65),
.B2(n_17),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_81),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_69),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_60),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_35),
.B1(n_41),
.B2(n_36),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_14),
.C(n_13),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_123),
.A2(n_124),
.B(n_108),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_98),
.B(n_100),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_133),
.B1(n_134),
.B2(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_135),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_137),
.B(n_123),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_137),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_104),
.B1(n_108),
.B2(n_92),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_104),
.B1(n_102),
.B2(n_65),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_105),
.B(n_83),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_111),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_141),
.C(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_122),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_147),
.B(n_80),
.Y(n_154)
);

OAI321xp33_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_130),
.A3(n_123),
.B1(n_133),
.B2(n_126),
.C(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_68),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_28),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_136),
.C(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_140),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_31),
.C(n_17),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_159),
.B(n_31),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_134),
.B1(n_143),
.B2(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_152),
.B1(n_148),
.B2(n_82),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_159),
.A3(n_28),
.B1(n_7),
.B2(n_12),
.C1(n_13),
.C2(n_11),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_163),
.A3(n_11),
.B1(n_2),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_151),
.B1(n_29),
.B2(n_8),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g164 ( 
.A(n_160),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_4),
.B(n_5),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_166),
.B(n_1),
.C(n_4),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_6),
.Y(n_170)
);


endmodule