module fake_jpeg_23411_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_21),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

CKINVDCx12_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx12_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_14),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_21),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_17),
.B(n_15),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_20),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_47),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_24),
.B2(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_33),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_12),
.A3(n_10),
.B1(n_19),
.B2(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_27),
.C(n_28),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_52),
.C(n_39),
.Y(n_68)
);

OAI22x1_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR4xp25_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_45),
.C(n_52),
.D(n_39),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_63),
.C(n_66),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.C(n_72),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_17),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_39),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_22),
.C(n_11),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_14),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_79),
.B(n_84),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_58),
.B(n_30),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_58),
.B1(n_24),
.B2(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_70),
.C(n_13),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_1),
.C(n_2),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_84),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_71),
.B(n_8),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_85),
.B(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_4),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_18),
.B1(n_23),
.B2(n_3),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_9),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_1),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_97),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_104),
.B(n_101),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_2),
.C(n_3),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_23),
.Y(n_108)
);


endmodule