module fake_aes_7690_n_28 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
BUFx6f_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
OAI22xp5_ASAP7_75t_SL g16 ( .A1(n_5), .A2(n_12), .B1(n_4), .B2(n_1), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
A2O1A1Ixp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_17), .B(n_13), .C(n_16), .Y(n_20) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_20), .B(n_18), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
OAI221xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_16), .B1(n_17), .B2(n_13), .C(n_3), .Y(n_24) );
NAND4xp75_ASAP7_75t_L g25 ( .A(n_24), .B(n_0), .C(n_1), .D(n_2), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
OAI22xp5_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_4), .B1(n_7), .B2(n_11), .Y(n_28) );
endmodule