module fake_jpeg_22568_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_7),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_15),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_16),
.B1(n_27),
.B2(n_15),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_19),
.B2(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_0),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_25),
.B(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_19),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_47),
.B1(n_46),
.B2(n_41),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_34),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_63),
.Y(n_84)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_68),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_72),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_54),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_24),
.B1(n_26),
.B2(n_14),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_42),
.B1(n_14),
.B2(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_25),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_50),
.B1(n_39),
.B2(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_39),
.B1(n_42),
.B2(n_53),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_51),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_49),
.B1(n_40),
.B2(n_24),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_51),
.B1(n_44),
.B2(n_40),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_33),
.B(n_24),
.C(n_14),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_60),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_78),
.B1(n_76),
.B2(n_93),
.Y(n_120)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_101),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_74),
.C(n_69),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_105),
.C(n_59),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_77),
.Y(n_101)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_107),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_63),
.Y(n_104)
);

XNOR2x1_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_110),
.Y(n_129)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_64),
.A3(n_62),
.B1(n_61),
.B2(n_44),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_90),
.B(n_95),
.C(n_94),
.D(n_62),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_121),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_113),
.B1(n_106),
.B2(n_95),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_125),
.B1(n_102),
.B2(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_103),
.B1(n_109),
.B2(n_104),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_108),
.B1(n_102),
.B2(n_109),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_80),
.B(n_88),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_62),
.B(n_71),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_89),
.B1(n_87),
.B2(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

AO221x1_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_132),
.B1(n_101),
.B2(n_96),
.C(n_64),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_83),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_139),
.B1(n_140),
.B2(n_148),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_132),
.C(n_128),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_144),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_146),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_142),
.B(n_116),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_44),
.C(n_62),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_122),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_10),
.A3(n_11),
.B1(n_13),
.B2(n_12),
.C1(n_4),
.C2(n_5),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_9),
.C(n_13),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_11),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_75),
.B1(n_51),
.B2(n_61),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_123),
.A3(n_130),
.B1(n_119),
.B2(n_124),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_133),
.C(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_154),
.B(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_145),
.B(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_4),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_135),
.B1(n_131),
.B2(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_153),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_120),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_160),
.C(n_159),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_172),
.B(n_23),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_158),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_174),
.C(n_181),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_152),
.C(n_165),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_180),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_176),
.B(n_178),
.Y(n_186)
);

NOR2xp67_ASAP7_75t_SL g183 ( 
.A(n_179),
.B(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_166),
.A3(n_75),
.B1(n_14),
.B2(n_22),
.C1(n_6),
.C2(n_7),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_22),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_187),
.B(n_8),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_0),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_6),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_174),
.B1(n_175),
.B2(n_22),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_8),
.C(n_11),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_182),
.Y(n_195)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_1),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_1),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_8),
.B(n_2),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_197),
.A2(n_3),
.B(n_1),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_1),
.B1(n_3),
.B2(n_201),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_200),
.A2(n_201),
.B1(n_198),
.B2(n_2),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule