module fake_jpeg_11597_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_9),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_63),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_64),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_72),
.B(n_89),
.Y(n_158)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_75),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_78),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_83),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_94),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_97),
.B(n_98),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_0),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_37),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_99),
.B(n_102),
.Y(n_175)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_37),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_106),
.Y(n_210)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_37),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_42),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_123),
.Y(n_134)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_30),
.B(n_1),
.Y(n_115)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_35),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_53),
.Y(n_141)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_30),
.B(n_2),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_27),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_42),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_45),
.Y(n_124)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_36),
.Y(n_126)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

BUFx4f_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_80),
.A2(n_56),
.B1(n_35),
.B2(n_53),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_130),
.A2(n_176),
.B1(n_202),
.B2(n_67),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_133),
.B(n_141),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_164),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_27),
.B1(n_53),
.B2(n_19),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_137),
.A2(n_48),
.B1(n_46),
.B2(n_29),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_19),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_109),
.A2(n_19),
.B1(n_56),
.B2(n_47),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_162),
.A2(n_177),
.B1(n_215),
.B2(n_76),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_52),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_75),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_182),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_70),
.A2(n_52),
.B(n_47),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_172),
.B(n_73),
.C(n_82),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_71),
.A2(n_24),
.B1(n_40),
.B2(n_38),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_38),
.B1(n_31),
.B2(n_32),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_75),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_81),
.B(n_55),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_106),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_200),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_106),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_116),
.B(n_55),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_121),
.B(n_46),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_221),
.Y(n_232)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_111),
.A2(n_40),
.B1(n_32),
.B2(n_31),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_101),
.Y(n_216)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

BUFx2_ASAP7_75t_R g220 ( 
.A(n_63),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g230 ( 
.A(n_220),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_128),
.B(n_48),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_224),
.Y(n_310)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx4_ASAP7_75t_SL g360 ( 
.A(n_226),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_134),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_264),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_236),
.A2(n_270),
.B1(n_219),
.B2(n_185),
.Y(n_319)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_237),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_29),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_238),
.B(n_267),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_133),
.B(n_25),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_239),
.B(n_255),
.Y(n_308)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_144),
.Y(n_246)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_246),
.Y(n_344)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_150),
.Y(n_249)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_254),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_145),
.B(n_25),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_103),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_256),
.B(n_261),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_130),
.A2(n_95),
.B1(n_94),
.B2(n_88),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_257),
.A2(n_132),
.B1(n_146),
.B2(n_192),
.Y(n_348)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_258),
.Y(n_328)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_156),
.Y(n_259)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_259),
.Y(n_347)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_158),
.B(n_154),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_156),
.Y(n_262)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_147),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_191),
.A2(n_61),
.B1(n_85),
.B2(n_60),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_265),
.A2(n_274),
.B1(n_278),
.B2(n_279),
.Y(n_331)
);

BUFx16f_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx5_ASAP7_75t_SL g353 ( 
.A(n_266),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_158),
.B(n_2),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_162),
.A2(n_84),
.B1(n_62),
.B2(n_77),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_183),
.Y(n_271)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_271),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_275),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_173),
.B(n_152),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_273),
.B(n_283),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_191),
.A2(n_68),
.B1(n_66),
.B2(n_65),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_147),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_281),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_165),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_142),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_292),
.Y(n_335)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_151),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_284),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_173),
.B(n_2),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_289),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_164),
.B(n_3),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_287),
.B(n_290),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_163),
.A2(n_82),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_288),
.A2(n_291),
.B1(n_297),
.B2(n_139),
.Y(n_351)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_135),
.B(n_3),
.Y(n_290)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_174),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_138),
.B(n_4),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_293),
.B(n_294),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_140),
.B(n_4),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_168),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_296),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_177),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_184),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_198),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_298),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_143),
.B(n_4),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_300),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_166),
.B(n_6),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_167),
.B(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_7),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_141),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_306),
.B(n_312),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_270),
.A2(n_215),
.B1(n_176),
.B2(n_203),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_307),
.A2(n_319),
.B1(n_321),
.B2(n_350),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_228),
.A2(n_185),
.B1(n_203),
.B2(n_132),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_232),
.B(n_195),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_327),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_159),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_257),
.A2(n_131),
.B1(n_187),
.B2(n_178),
.Y(n_329)
);

OA22x2_ASAP7_75t_L g396 ( 
.A1(n_329),
.A2(n_338),
.B1(n_354),
.B2(n_244),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_231),
.B(n_157),
.C(n_210),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_330),
.B(n_340),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_229),
.A2(n_131),
.B1(n_187),
.B2(n_178),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_275),
.B(n_210),
.C(n_161),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_233),
.B(n_160),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_346),
.Y(n_374)
);

A2O1A1O1Ixp25_ASAP7_75t_L g343 ( 
.A1(n_223),
.A2(n_188),
.B(n_214),
.C(n_153),
.D(n_161),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_343),
.A2(n_226),
.B(n_227),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_243),
.B(n_219),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_348),
.A2(n_237),
.B1(n_235),
.B2(n_241),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_274),
.A2(n_194),
.B1(n_192),
.B2(n_184),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_351),
.A2(n_249),
.B1(n_259),
.B2(n_247),
.Y(n_383)
);

AO22x2_ASAP7_75t_SL g354 ( 
.A1(n_265),
.A2(n_155),
.B1(n_194),
.B2(n_214),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_288),
.A2(n_155),
.B1(n_42),
.B2(n_10),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_355),
.A2(n_358),
.B1(n_284),
.B2(n_282),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_297),
.A2(n_42),
.B1(n_9),
.B2(n_12),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_230),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_266),
.Y(n_363)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_363),
.B(n_371),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_342),
.A2(n_248),
.B1(n_260),
.B2(n_291),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_364),
.A2(n_383),
.B1(n_387),
.B2(n_397),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_225),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_365),
.B(n_370),
.Y(n_444)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_310),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_369),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_252),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_332),
.B(n_292),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_308),
.B(n_280),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_376),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_345),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_375),
.B(n_390),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_266),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_353),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_381),
.Y(n_411)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_339),
.Y(n_379)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_379),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_240),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_269),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_384),
.B(n_385),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g386 ( 
.A(n_320),
.B(n_269),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_SL g424 ( 
.A1(n_386),
.A2(n_331),
.B(n_360),
.C(n_334),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_244),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_388),
.B(n_398),
.Y(n_413)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_389),
.Y(n_436)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_311),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_392),
.Y(n_423)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_302),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_268),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_394),
.Y(n_426)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_337),
.Y(n_394)
);

OAI21xp33_ASAP7_75t_SL g412 ( 
.A1(n_396),
.A2(n_405),
.B(n_313),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_320),
.A2(n_253),
.B1(n_278),
.B2(n_276),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_246),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_302),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_400),
.Y(n_431)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_336),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_403),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_402),
.A2(n_307),
.B1(n_321),
.B2(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_241),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_406),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_310),
.Y(n_405)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_317),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_347),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_235),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_408),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_410),
.A2(n_416),
.B1(n_418),
.B2(n_425),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_412),
.A2(n_402),
.B1(n_378),
.B2(n_384),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_320),
.B1(n_313),
.B2(n_340),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_306),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_419),
.C(n_422),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_355),
.B1(n_322),
.B2(n_348),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_330),
.C(n_361),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_357),
.C(n_314),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_424),
.A2(n_427),
.B(n_356),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_398),
.B1(n_374),
.B2(n_373),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_385),
.A2(n_324),
.B(n_328),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_393),
.A2(n_404),
.B(n_374),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_398),
.A2(n_333),
.B1(n_352),
.B2(n_318),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_433),
.A2(n_369),
.B1(n_390),
.B2(n_399),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_326),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_419),
.C(n_417),
.Y(n_461)
);

AND2x2_ASAP7_75t_SL g437 ( 
.A(n_367),
.B(n_325),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_437),
.B(n_389),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_362),
.A2(n_326),
.B(n_328),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_436),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_375),
.B(n_333),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_377),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_448),
.A2(n_452),
.B(n_454),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_423),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_465),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_386),
.Y(n_452)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_371),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_455),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_401),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_456),
.B(n_459),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_439),
.A2(n_373),
.B1(n_396),
.B2(n_391),
.Y(n_457)
);

OAI22x1_ASAP7_75t_SL g515 ( 
.A1(n_457),
.A2(n_458),
.B1(n_472),
.B2(n_434),
.Y(n_515)
);

AOI22x1_ASAP7_75t_L g458 ( 
.A1(n_439),
.A2(n_396),
.B1(n_397),
.B2(n_387),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_415),
.B(n_368),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_396),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_463),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_480),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_395),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_462),
.B(n_437),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_395),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_464),
.B(n_413),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_407),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_475),
.Y(n_501)
);

OA22x2_ASAP7_75t_L g468 ( 
.A1(n_410),
.A2(n_425),
.B1(n_418),
.B2(n_424),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_457),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_403),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_429),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_432),
.A2(n_400),
.B1(n_366),
.B2(n_405),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_470),
.A2(n_471),
.B1(n_481),
.B2(n_430),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_420),
.A2(n_405),
.B1(n_392),
.B2(n_347),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_414),
.A2(n_434),
.B1(n_420),
.B2(n_447),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_360),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_476),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_477),
.A2(n_434),
.B(n_446),
.Y(n_496)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_478),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_409),
.A2(n_394),
.B1(n_262),
.B2(n_279),
.Y(n_479)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_479),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_344),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_427),
.A2(n_224),
.B1(n_339),
.B2(n_344),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_461),
.B(n_437),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_513),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_477),
.B(n_455),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_512),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_411),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_489),
.B(n_494),
.Y(n_519)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_493),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_440),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_450),
.B(n_440),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_495),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_496),
.A2(n_507),
.B(n_448),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_441),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_481),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_467),
.B(n_430),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_483),
.B(n_426),
.Y(n_505)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_483),
.B(n_426),
.Y(n_508)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_472),
.B(n_423),
.Y(n_510)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_510),
.Y(n_530)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_511),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_455),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_413),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_464),
.B(n_441),
.Y(n_514)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_514),
.Y(n_538)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_515),
.Y(n_541)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_516),
.Y(n_542)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_518),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_520),
.B(n_539),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_501),
.Y(n_521)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_521),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_523),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_449),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_525),
.B(n_515),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_507),
.A2(n_460),
.B1(n_468),
.B2(n_454),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_528),
.A2(n_541),
.B1(n_536),
.B2(n_535),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_531),
.A2(n_536),
.B(n_537),
.Y(n_552)
);

XOR2x2_ASAP7_75t_L g532 ( 
.A(n_485),
.B(n_463),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_547),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_502),
.A2(n_475),
.B(n_452),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g568 ( 
.A1(n_535),
.A2(n_501),
.B(n_493),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_502),
.A2(n_458),
.B(n_475),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_496),
.A2(n_468),
.B(n_458),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_500),
.B(n_431),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_487),
.B(n_468),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_545),
.Y(n_563)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_503),
.Y(n_543)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_543),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_422),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_431),
.B(n_442),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_546),
.A2(n_501),
.B(n_511),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_505),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_512),
.C(n_499),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_551),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_497),
.C(n_490),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_519),
.Y(n_554)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_544),
.A2(n_500),
.B1(n_517),
.B2(n_490),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_555),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_556),
.A2(n_568),
.B(n_526),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_557),
.B(n_560),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_497),
.C(n_514),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_558),
.B(n_527),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_532),
.B(n_508),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_562),
.B(n_537),
.Y(n_582)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_543),
.Y(n_565)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_565),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_524),
.B(n_510),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g580 ( 
.A(n_566),
.B(n_524),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_528),
.A2(n_533),
.B1(n_541),
.B2(n_530),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_567),
.A2(n_521),
.B1(n_530),
.B2(n_529),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_533),
.A2(n_517),
.B1(n_516),
.B2(n_504),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_569),
.B(n_571),
.Y(n_579)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_570),
.A2(n_527),
.B1(n_529),
.B2(n_526),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_547),
.A2(n_509),
.B1(n_506),
.B2(n_491),
.Y(n_571)
);

CKINVDCx11_ASAP7_75t_R g573 ( 
.A(n_549),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_573),
.B(n_588),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_522),
.Y(n_574)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_574),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_580),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_558),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_578),
.B(n_585),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_582),
.B(n_590),
.Y(n_597)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_584),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_546),
.C(n_542),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_589),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_531),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_552),
.Y(n_602)
);

FAx1_ASAP7_75t_SL g588 ( 
.A(n_550),
.B(n_523),
.CI(n_538),
.CON(n_588),
.SN(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_542),
.C(n_545),
.Y(n_589)
);

XOR2x1_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_560),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_SL g620 ( 
.A(n_591),
.B(n_602),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_572),
.A2(n_562),
.B1(n_567),
.B2(n_559),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_592),
.B(n_600),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_594),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_553),
.C(n_557),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_595),
.B(n_601),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_580),
.B(n_563),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_585),
.B(n_568),
.C(n_559),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_561),
.C(n_556),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_604),
.B(n_606),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_587),
.B(n_569),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_552),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_607),
.B(n_588),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_603),
.B(n_579),
.C(n_576),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_613),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_605),
.Y(n_611)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_611),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_593),
.B(n_590),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_600),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_579),
.C(n_577),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_616),
.B(n_617),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_598),
.A2(n_572),
.B1(n_574),
.B2(n_581),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_593),
.B(n_504),
.C(n_538),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_618),
.B(n_619),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_591),
.B(n_588),
.C(n_509),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_611),
.A2(n_599),
.B(n_597),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_621),
.A2(n_625),
.B(n_626),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_615),
.B(n_597),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_594),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_610),
.A2(n_506),
.B1(n_492),
.B2(n_491),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_628),
.B(n_629),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_608),
.A2(n_492),
.B1(n_486),
.B2(n_328),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_630),
.B(n_258),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_627),
.B(n_609),
.C(n_612),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_634),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_624),
.B(n_620),
.Y(n_634)
);

AOI322xp5_ASAP7_75t_L g635 ( 
.A1(n_623),
.A2(n_626),
.A3(n_624),
.B1(n_622),
.B2(n_620),
.C1(n_258),
.C2(n_316),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_635),
.B(n_305),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_636),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_627),
.B(n_316),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_305),
.B(n_9),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_639),
.Y(n_642)
);

AOI322xp5_ASAP7_75t_L g643 ( 
.A1(n_640),
.A2(n_636),
.A3(n_632),
.B1(n_633),
.B2(n_13),
.C1(n_7),
.C2(n_12),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_641),
.B(n_638),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_644),
.Y(n_645)
);

OAI31xp33_ASAP7_75t_SL g646 ( 
.A1(n_645),
.A2(n_642),
.A3(n_12),
.B(n_13),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_9),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_647),
.B(n_13),
.Y(n_648)
);


endmodule