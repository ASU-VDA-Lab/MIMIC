module fake_jpeg_7952_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_17),
.B1(n_23),
.B2(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_15),
.B1(n_30),
.B2(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_38),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_31),
.C(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_32),
.Y(n_57)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_62),
.CON(n_100),
.SN(n_100)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_74),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_17),
.B1(n_22),
.B2(n_16),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_69),
.B1(n_76),
.B2(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_68),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_15),
.B1(n_19),
.B2(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_82),
.B1(n_47),
.B2(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_30),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_29),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_33),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_18),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_26),
.B1(n_28),
.B2(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_97),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_37),
.C(n_38),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_96),
.B(n_101),
.C(n_97),
.D(n_94),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_131),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_124),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_79),
.B1(n_68),
.B2(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_118),
.B1(n_92),
.B2(n_89),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_72),
.B(n_37),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_92),
.B(n_18),
.Y(n_140)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_119),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_64),
.B1(n_59),
.B2(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_59),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_66),
.Y(n_122)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_108),
.B(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_38),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_73),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_35),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_87),
.C(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_28),
.B(n_18),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_108),
.B(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_63),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_137),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_90),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_89),
.B(n_104),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_18),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_149),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_148),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_112),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_108),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_118),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_121),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_131),
.Y(n_173)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_165),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_140),
.B(n_119),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_123),
.B1(n_146),
.B2(n_113),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_174),
.B1(n_133),
.B2(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_170),
.B(n_160),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_126),
.B1(n_120),
.B2(n_114),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_189),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_138),
.B1(n_151),
.B2(n_145),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_184),
.B1(n_174),
.B2(n_163),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_149),
.C(n_138),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_189),
.C(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_148),
.B1(n_155),
.B2(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_159),
.B1(n_169),
.B2(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_139),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_194),
.C(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_186),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_195),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_172),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_172),
.B(n_158),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_197),
.B(n_201),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_127),
.B(n_13),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_105),
.B(n_98),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_186),
.B1(n_177),
.B2(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_2),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_207),
.C(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_208),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_12),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_200),
.B1(n_4),
.B2(n_5),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_190),
.C(n_201),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_199),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_219),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_212),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_12),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_214),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_207),
.Y(n_221)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_213),
.C(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_11),
.C(n_4),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_3),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_10),
.C2(n_158),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_6),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_232),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_230),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_231),
.B1(n_233),
.B2(n_10),
.C(n_6),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_8),
.Y(n_236)
);


endmodule