module fake_jpeg_22462_n_291 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_35),
.Y(n_72)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_27),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_21),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_23),
.B1(n_26),
.B2(n_21),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_50),
.A2(n_64),
.B1(n_71),
.B2(n_22),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_53),
.B(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_25),
.B1(n_19),
.B2(n_38),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_59),
.A2(n_61),
.B1(n_24),
.B2(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_67),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_34),
.B1(n_23),
.B2(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_62),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_63),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_34),
.B1(n_25),
.B2(n_19),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_72),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_25),
.C(n_38),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_75),
.C(n_58),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_18),
.B1(n_35),
.B2(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_76),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_28),
.B(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_1),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_80),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_46),
.B1(n_24),
.B2(n_29),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_66),
.B1(n_55),
.B2(n_3),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_41),
.B1(n_46),
.B2(n_37),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_87),
.B1(n_83),
.B2(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_37),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_97),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_37),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_118),
.C(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_32),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_50),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_115),
.B1(n_83),
.B2(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_32),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_111),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_31),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_22),
.C(n_2),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_68),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_52),
.B(n_22),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_122),
.B(n_125),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_124),
.B1(n_134),
.B2(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_69),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_64),
.B1(n_77),
.B2(n_86),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_130),
.B1(n_142),
.B2(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_120),
.C(n_117),
.Y(n_159)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_59),
.B1(n_52),
.B2(n_67),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_133),
.Y(n_165)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_94),
.B1(n_90),
.B2(n_93),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_84),
.B1(n_68),
.B2(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_140),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_151),
.B1(n_118),
.B2(n_101),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_145),
.Y(n_182)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_16),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_1),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_55),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_2),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_167),
.B1(n_157),
.B2(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_102),
.B1(n_113),
.B2(n_106),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_176),
.B1(n_133),
.B2(n_149),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_172),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_103),
.Y(n_163)
);

AO21x2_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_93),
.B(n_112),
.Y(n_167)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_93),
.C(n_101),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_181),
.B(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_95),
.B1(n_104),
.B2(n_112),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_95),
.Y(n_179)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_104),
.B(n_6),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_137),
.A2(n_123),
.B(n_130),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_184),
.B(n_142),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_122),
.A2(n_100),
.B(n_7),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_190),
.B(n_191),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_196),
.B1(n_200),
.B2(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_188),
.B(n_192),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_100),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_138),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_162),
.B(n_128),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_177),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_144),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_182),
.B(n_156),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_204),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_165),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_167),
.B1(n_173),
.B2(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_12),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_218),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_201),
.B1(n_200),
.B2(n_194),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_166),
.B(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_215),
.B(n_227),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_167),
.B1(n_166),
.B2(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_189),
.B1(n_197),
.B2(n_156),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_159),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_219),
.B(n_203),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_163),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.C(n_190),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_155),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_208),
.A2(n_183),
.B1(n_158),
.B2(n_184),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_207),
.B1(n_188),
.B2(n_197),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_231),
.C(n_223),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_207),
.C(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_239),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_242),
.B1(n_219),
.B2(n_224),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_238),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_160),
.B1(n_187),
.B2(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_160),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_187),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_225),
.B(n_212),
.C(n_209),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_249),
.B(n_257),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_255),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_258),
.B1(n_248),
.B2(n_234),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_244),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_256),
.B1(n_234),
.B2(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_211),
.B(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_229),
.B1(n_233),
.B2(n_235),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_249),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_232),
.B1(n_237),
.B2(n_231),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_237),
.B1(n_230),
.B2(n_235),
.Y(n_264)
);

NAND4xp25_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_215),
.C(n_221),
.D(n_154),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_252),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_275),
.B(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_251),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_268),
.B(n_254),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_257),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_265),
.B(n_260),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_211),
.B(n_168),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_263),
.B1(n_272),
.B2(n_222),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_279),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_14),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_285),
.C(n_12),
.Y(n_288)
);

OAI21x1_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_289),
.B(n_14),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_14),
.Y(n_291)
);


endmodule