module real_aes_8496_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_10;
INVx1_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
INVx1_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
OAI221xp5_ASAP7_75t_L g25 ( .A1(n_2), .A2(n_4), .B1(n_8), .B2(n_26), .C(n_27), .Y(n_25) );
INVxp67_ASAP7_75t_L g28 ( .A(n_2), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_3), .Y(n_26) );
INVxp67_ASAP7_75t_L g29 ( .A(n_4), .Y(n_29) );
NAND3xp33_ASAP7_75t_SL g12 ( .A(n_5), .B(n_13), .C(n_14), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_6), .B(n_24), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_10), .B(n_21), .Y(n_9) );
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_11), .B(n_17), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
AND2x2_ASAP7_75t_L g21 ( .A(n_18), .B(n_22), .Y(n_21) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_23), .Y(n_22) );
INVxp67_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_28), .B(n_29), .Y(n_27) );
endmodule