module real_jpeg_1907_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_25),
.B1(n_36),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_2),
.A2(n_30),
.B1(n_64),
.B2(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_64),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_125),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_5),
.B(n_56),
.C(n_58),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_55),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_5),
.B(n_40),
.C(n_87),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_5),
.B(n_44),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_5),
.B(n_91),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_5),
.A2(n_25),
.B1(n_34),
.B2(n_36),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_10),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_13),
.A2(n_25),
.B1(n_36),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_13),
.A2(n_30),
.B1(n_52),
.B2(n_69),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_13),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_52),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_14),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_14),
.A2(n_25),
.B1(n_36),
.B2(n_84),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_84),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_15),
.A2(n_30),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_15),
.A2(n_25),
.B1(n_36),
.B2(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_68),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_20),
.B(n_105),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_92),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_21),
.B(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_49),
.C(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_23),
.A2(n_24),
.B1(n_37),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.A3(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_36),
.B1(n_56),
.B2(n_60),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_70)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_69),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_30),
.A2(n_33),
.B(n_34),
.C(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_34),
.A2(n_79),
.B(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_36),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_37),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_149),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_39),
.A2(n_40),
.B1(n_87),
.B2(n_88),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_40),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_42),
.A2(n_43),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_42),
.B(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_42),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_42),
.A2(n_43),
.B1(n_178),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_43),
.A2(n_149),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_43),
.B(n_169),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_46),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_44),
.A2(n_168),
.B(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_65),
.B2(n_76),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_62),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_53),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_53),
.A2(n_62),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_54),
.B(n_63),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_55)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_58),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_58),
.B(n_192),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_71),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_67),
.A2(n_74),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_92),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_82),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_158),
.B(n_160),
.Y(n_157)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_85),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_89),
.A2(n_95),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_89),
.A2(n_159),
.B1(n_186),
.B2(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_91),
.B(n_96),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_102),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_93),
.B(n_102),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_98),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_103),
.A2(n_104),
.B(n_129),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_119),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_130),
.B2(n_131),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_150),
.B(n_230),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_136),
.B(n_138),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_144),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.C(n_148),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_172),
.B(n_229),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_170),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_170),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_162),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_154),
.B(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_162),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_161),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_224),
.B(n_228),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_214),
.B(n_223),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_196),
.B(n_213),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_189),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_189),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_184),
.C(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_207),
.B(n_212),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_202),
.B(n_206),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_205),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_210),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_220),
.C(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_227),
.Y(n_228)
);


endmodule