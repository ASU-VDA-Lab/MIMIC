module fake_jpeg_26023_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_12),
.B(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_50),
.B1(n_57),
.B2(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_24),
.B1(n_33),
.B2(n_18),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_43),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_33),
.B1(n_24),
.B2(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_62),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_24),
.B1(n_33),
.B2(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_16),
.B1(n_18),
.B2(n_32),
.Y(n_87)
);

OAI22x1_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_44),
.B1(n_37),
.B2(n_19),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_74),
.B1(n_87),
.B2(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_76),
.Y(n_95)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_38),
.B1(n_27),
.B2(n_16),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_30),
.B1(n_36),
.B2(n_20),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_80),
.B1(n_85),
.B2(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_32),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_83),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_30),
.B1(n_20),
.B2(n_25),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_59),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_30),
.B1(n_20),
.B2(n_32),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_67),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_65),
.B1(n_46),
.B2(n_45),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_84),
.B1(n_73),
.B2(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_107),
.B1(n_69),
.B2(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_106),
.B(n_109),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_68),
.B(n_54),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_61),
.B(n_45),
.C(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_58),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_63),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_54),
.C(n_63),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_119),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_123),
.B1(n_126),
.B2(n_108),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_86),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_129),
.B1(n_110),
.B2(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_71),
.B1(n_70),
.B2(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_71),
.B1(n_77),
.B2(n_80),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_102),
.B1(n_96),
.B2(n_107),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_91),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_85),
.A3(n_68),
.B1(n_30),
.B2(n_43),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_97),
.B1(n_100),
.B2(n_107),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_109),
.B(n_90),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_131),
.B(n_124),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_145),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_94),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_146),
.B1(n_155),
.B2(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_151),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_93),
.B1(n_68),
.B2(n_86),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_149),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_153),
.Y(n_168)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_0),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_125),
.B1(n_116),
.B2(n_129),
.Y(n_155)
);

XOR2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_117),
.Y(n_156)
);

XOR2x1_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_3),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_170),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_173),
.C(n_174),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_128),
.B1(n_119),
.B2(n_43),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_135),
.B1(n_147),
.B2(n_141),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_41),
.C(n_1),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_41),
.C(n_1),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_0),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_143),
.C(n_152),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_183),
.B1(n_167),
.B2(n_160),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_143),
.A3(n_134),
.B1(n_146),
.B2(n_140),
.C1(n_142),
.C2(n_136),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_134),
.B1(n_151),
.B2(n_5),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_168),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_190),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_15),
.C(n_4),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_187),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_165),
.B(n_4),
.C(n_6),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_191),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_6),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_159),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_164),
.B1(n_166),
.B2(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_205),
.B1(n_201),
.B2(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_172),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_160),
.B1(n_162),
.B2(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_185),
.B(n_171),
.CI(n_175),
.CON(n_204),
.SN(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_174),
.B1(n_167),
.B2(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

AO22x1_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_192),
.B1(n_180),
.B2(n_190),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_189),
.B(n_186),
.Y(n_209)
);

OAI221xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_200),
.B1(n_198),
.B2(n_197),
.C(n_11),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_198),
.B(n_9),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_215),
.A2(n_210),
.B1(n_208),
.B2(n_207),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_14),
.B(n_11),
.C(n_12),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_209),
.B(n_11),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_10),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);


endmodule