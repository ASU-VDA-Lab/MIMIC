module fake_ibex_514_n_3595 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3595);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3595;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_3272;
wire n_3255;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_2230;
wire n_963;
wire n_1782;
wire n_1856;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2333;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_662;
wire n_3097;
wire n_3030;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_709;
wire n_3060;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1806;
wire n_1599;
wire n_2842;
wire n_3070;
wire n_2711;
wire n_3477;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_3557;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_3383;
wire n_2884;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2654;
wire n_2463;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_3314;
wire n_2997;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_961;
wire n_991;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3376;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_3427;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3333;
wire n_3096;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_1455;
wire n_804;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_3044;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_946;
wire n_707;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_645;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_714;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_750;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_665;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3430;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_2928;
wire n_3225;
wire n_2227;
wire n_3380;
wire n_3483;
wire n_1074;
wire n_3067;
wire n_2652;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_704;
wire n_2104;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_683;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_3482;
wire n_2282;
wire n_970;
wire n_2673;
wire n_2430;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

INVx2_ASAP7_75t_L g642 ( 
.A(n_621),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_157),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_450),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_333),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_160),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_338),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_348),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_107),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_111),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_226),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_582),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_421),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_511),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_128),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_297),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_19),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_476),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_307),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_24),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_94),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_543),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_291),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_31),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_105),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_542),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_118),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_563),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_386),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_153),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_41),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_534),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_261),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_553),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_581),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_552),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_282),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_311),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_495),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_503),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_316),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_594),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_27),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_500),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_381),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_600),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_51),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_223),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_492),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_170),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_404),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_399),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_173),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_137),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_225),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_569),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_85),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_513),
.B(n_388),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_49),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_173),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_255),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_527),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_309),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_595),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_518),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_584),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_129),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_29),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_374),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_629),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_603),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_238),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_323),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_526),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_5),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_383),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_387),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_151),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_34),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_604),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_614),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_42),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_150),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_21),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_376),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_305),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_514),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_396),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_512),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_221),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_570),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_70),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_91),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_167),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_354),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_554),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_244),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_206),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_73),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_282),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_412),
.Y(n_742)
);

BUFx5_ASAP7_75t_L g743 ( 
.A(n_519),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_370),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_489),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_533),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_616),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_79),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_132),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_625),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_99),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_639),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_300),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_189),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_467),
.Y(n_755)
);

CKINVDCx16_ASAP7_75t_R g756 ( 
.A(n_459),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_565),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_447),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_64),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_472),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_545),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_256),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_227),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_36),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_183),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_499),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_336),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_355),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_4),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_388),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_365),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_485),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_179),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_567),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_245),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_152),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_180),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_293),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_636),
.Y(n_779)
);

CKINVDCx14_ASAP7_75t_R g780 ( 
.A(n_200),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_314),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_608),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_307),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_428),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_276),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_318),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_607),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_201),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_61),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_227),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_91),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_525),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_360),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_483),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_70),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_151),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_68),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_247),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_178),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_187),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_387),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_22),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_537),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_331),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_98),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_267),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_566),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_89),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_508),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_568),
.B(n_308),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_548),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_369),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_530),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_246),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_481),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_638),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_371),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_487),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_346),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_226),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_609),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_78),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_121),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_294),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_486),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_586),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_403),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_28),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_84),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_478),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_287),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_64),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_377),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_105),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_56),
.B(n_342),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_237),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_339),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_365),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_306),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_141),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_120),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_539),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_97),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_632),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_294),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_259),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_141),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_599),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_463),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_93),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_207),
.B(n_316),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_597),
.B(n_117),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_208),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_540),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_515),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_358),
.Y(n_856)
);

CKINVDCx14_ASAP7_75t_R g857 ( 
.A(n_598),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_602),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_438),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_520),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_615),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_402),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_230),
.Y(n_863)
);

CKINVDCx14_ASAP7_75t_R g864 ( 
.A(n_470),
.Y(n_864)
);

CKINVDCx14_ASAP7_75t_R g865 ( 
.A(n_169),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_640),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_381),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_9),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_613),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_334),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_0),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_356),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_220),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_529),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_521),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_641),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_418),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_457),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_111),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_453),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_386),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_149),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_634),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_460),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_100),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_633),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_350),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_612),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_178),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_48),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_228),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_100),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_314),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_215),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_466),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_398),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_410),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_497),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_237),
.Y(n_899)
);

CKINVDCx14_ASAP7_75t_R g900 ( 
.A(n_301),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_93),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_292),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_502),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_577),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_220),
.Y(n_905)
);

BUFx8_ASAP7_75t_SL g906 ( 
.A(n_309),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_494),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_435),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_87),
.Y(n_909)
);

CKINVDCx16_ASAP7_75t_R g910 ( 
.A(n_364),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_414),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_293),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_253),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_323),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_452),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_15),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_623),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_402),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_578),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_610),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_341),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_310),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_164),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_506),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_207),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_561),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_416),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_451),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_334),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_44),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_218),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_313),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_119),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_490),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_451),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_429),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_247),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_82),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_571),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_618),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_350),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_62),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_268),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_601),
.Y(n_944)
);

CKINVDCx14_ASAP7_75t_R g945 ( 
.A(n_459),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_143),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_52),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_113),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_422),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_433),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_76),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_1),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_538),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_453),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_88),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_624),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_452),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_37),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_415),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_181),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_541),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_45),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_573),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_206),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_239),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_188),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_436),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_510),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_535),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_177),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_278),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_18),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_174),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_522),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_131),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_383),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_362),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_174),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_300),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_159),
.Y(n_980)
);

BUFx8_ASAP7_75t_SL g981 ( 
.A(n_338),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_77),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_83),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_357),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_380),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_547),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_71),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_576),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_56),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_119),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_33),
.Y(n_991)
);

INVx4_ASAP7_75t_R g992 ( 
.A(n_107),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_236),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_325),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_263),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_257),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_375),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_204),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_403),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_155),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_373),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_404),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_596),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_215),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_287),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_346),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_456),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_199),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_190),
.Y(n_1009)
);

CKINVDCx16_ASAP7_75t_R g1010 ( 
.A(n_238),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_339),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_611),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_361),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_116),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_35),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_203),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_289),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_243),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_575),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_587),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_367),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_457),
.Y(n_1022)
);

BUFx2_ASAP7_75t_SL g1023 ( 
.A(n_436),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_332),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_572),
.Y(n_1025)
);

BUFx8_ASAP7_75t_SL g1026 ( 
.A(n_164),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_183),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_115),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_43),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_367),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_716),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_664),
.Y(n_1032)
);

NOR2x1_ASAP7_75t_L g1033 ( 
.A(n_716),
.B(n_462),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_652),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_780),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_732),
.Y(n_1036)
);

BUFx8_ASAP7_75t_SL g1037 ( 
.A(n_906),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_642),
.A2(n_465),
.B(n_464),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_780),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_865),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_743),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_716),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_801),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_743),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_642),
.A2(n_469),
.B(n_468),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_895),
.Y(n_1046)
);

BUFx12f_ASAP7_75t_L g1047 ( 
.A(n_674),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_865),
.Y(n_1048)
);

BUFx8_ASAP7_75t_L g1049 ( 
.A(n_757),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_743),
.Y(n_1050)
);

INVx6_ASAP7_75t_L g1051 ( 
.A(n_674),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_900),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_801),
.B(n_2),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_801),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_652),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_821),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_743),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_821),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_922),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_922),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_900),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_652),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_674),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_652),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_839),
.B(n_3),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_707),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_743),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_686),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_707),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_743),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_945),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_686),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_654),
.A2(n_473),
.B(n_471),
.Y(n_1073)
);

OAI22x1_ASAP7_75t_SL g1074 ( 
.A1(n_700),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_945),
.A2(n_756),
.B1(n_775),
.B2(n_740),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_743),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_686),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_673),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_654),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_697),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_697),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_931),
.B(n_7),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_773),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_970),
.B(n_7),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_673),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_863),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_805),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_664),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_664),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_805),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_686),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1024),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_827),
.Y(n_1093)
);

INVxp33_ASAP7_75t_SL g1094 ( 
.A(n_1029),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_827),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_889),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_707),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_910),
.B(n_6),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_669),
.Y(n_1099)
);

OA21x2_ASAP7_75t_L g1100 ( 
.A1(n_722),
.A2(n_475),
.B(n_474),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_1010),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_669),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_889),
.B(n_8),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_803),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1030),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_671),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_941),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1030),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_671),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_667),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_722),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_941),
.B(n_11),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_995),
.Y(n_1113)
);

BUFx8_ASAP7_75t_L g1114 ( 
.A(n_995),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_803),
.Y(n_1115)
);

BUFx8_ASAP7_75t_SL g1116 ( 
.A(n_906),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_803),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_695),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_794),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_695),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_888),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_888),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_888),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_794),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_830),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_830),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_710),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_1030),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_680),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1030),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_710),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_903),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1053),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1034),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_1069),
.B(n_1097),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1131),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1037),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1048),
.B(n_1061),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1037),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1116),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1116),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_1039),
.B(n_857),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1129),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1131),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1099),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1078),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1129),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1051),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1054),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1085),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1087),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1046),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1101),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1047),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1099),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1047),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1054),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1061),
.B(n_681),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1051),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1102),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1104),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_1040),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_R g1163 ( 
.A(n_1039),
.B(n_1071),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1104),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1069),
.B(n_996),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1121),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1090),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_1052),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1075),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_1121),
.B(n_857),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1122),
.Y(n_1171)
);

CKINVDCx16_ASAP7_75t_R g1172 ( 
.A(n_1122),
.Y(n_1172)
);

AND2x4_ASAP7_75t_SL g1173 ( 
.A(n_1097),
.B(n_1083),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_1123),
.B(n_1088),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1093),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_1123),
.B(n_864),
.Y(n_1176)
);

CKINVDCx16_ASAP7_75t_R g1177 ( 
.A(n_1083),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1092),
.B(n_864),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1036),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1036),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1095),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1096),
.Y(n_1182)
);

INVx11_ASAP7_75t_L g1183 ( 
.A(n_1049),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1049),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1094),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1102),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1086),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1113),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1094),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1114),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1114),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1086),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1051),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1034),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1106),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1063),
.B(n_903),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1106),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1120),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1107),
.A2(n_729),
.B1(n_751),
.B2(n_718),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1120),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1063),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1063),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1066),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_1098),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1109),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1059),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1088),
.B(n_1066),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1034),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1115),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1115),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1115),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1060),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1032),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1089),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1109),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1035),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1117),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1074),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1082),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_1056),
.Y(n_1221)
);

NAND2xp33_ASAP7_75t_R g1222 ( 
.A(n_1100),
.B(n_998),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_1084),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1058),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1103),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1058),
.Y(n_1226)
);

NAND2xp33_ASAP7_75t_R g1227 ( 
.A(n_1100),
.B(n_998),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1031),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1081),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1081),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_SL g1231 ( 
.A(n_1119),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1119),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1124),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1112),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1065),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1042),
.Y(n_1236)
);

INVxp33_ASAP7_75t_SL g1237 ( 
.A(n_1065),
.Y(n_1237)
);

NAND2xp33_ASAP7_75t_R g1238 ( 
.A(n_1100),
.B(n_1002),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1043),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1118),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1127),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1079),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_1033),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1079),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1125),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1080),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1080),
.B(n_897),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1111),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1111),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1126),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1132),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1132),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1041),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1125),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1041),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1125),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1044),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1044),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_R g1259 ( 
.A(n_1105),
.B(n_658),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1050),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1050),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1057),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1057),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1067),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1067),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1070),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1076),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1076),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1105),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1034),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1038),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1105),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1045),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1073),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1105),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1108),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1108),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1108),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_R g1279 ( 
.A(n_1108),
.B(n_1002),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1110),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1110),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1110),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1110),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1130),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1128),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1128),
.B(n_975),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1128),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1130),
.B(n_680),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1128),
.Y(n_1289)
);

INVxp33_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1055),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1055),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1055),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1055),
.Y(n_1294)
);

NAND2xp33_ASAP7_75t_R g1295 ( 
.A(n_1062),
.B(n_1021),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1062),
.B(n_1006),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1062),
.Y(n_1297)
);

NAND2xp33_ASAP7_75t_R g1298 ( 
.A(n_1062),
.B(n_1022),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1064),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1064),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1064),
.B(n_746),
.Y(n_1301)
);

CKINVDCx16_ASAP7_75t_R g1302 ( 
.A(n_1064),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1068),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1068),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1068),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1091),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_R g1307 ( 
.A(n_1072),
.B(n_1027),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1091),
.Y(n_1308)
);

NOR2x1_ASAP7_75t_L g1309 ( 
.A(n_1072),
.B(n_897),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1201),
.B(n_662),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1201),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1225),
.B(n_666),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1234),
.B(n_668),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1248),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1223),
.B(n_997),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1173),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1248),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1224),
.B(n_672),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1135),
.B(n_675),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1149),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1165),
.B(n_676),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1145),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1199),
.B(n_997),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1281),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_L g1326 ( 
.A(n_1190),
.B(n_703),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1244),
.B(n_705),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1226),
.B(n_706),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1246),
.B(n_711),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1149),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1250),
.B(n_1252),
.Y(n_1331)
);

NAND2xp33_ASAP7_75t_L g1332 ( 
.A(n_1191),
.B(n_712),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1157),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1155),
.Y(n_1334)
);

NOR3xp33_ASAP7_75t_L g1335 ( 
.A(n_1177),
.B(n_915),
.C(n_688),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1160),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1157),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1186),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1195),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1229),
.B(n_1230),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1162),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1187),
.B(n_646),
.Y(n_1342)
);

INVx8_ASAP7_75t_L g1343 ( 
.A(n_1193),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1146),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1271),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1150),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1221),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1192),
.B(n_785),
.Y(n_1348)
);

INVxp33_ASAP7_75t_L g1349 ( 
.A(n_1178),
.Y(n_1349)
);

NOR3xp33_ASAP7_75t_L g1350 ( 
.A(n_1200),
.B(n_841),
.C(n_786),
.Y(n_1350)
);

NOR3xp33_ASAP7_75t_L g1351 ( 
.A(n_1185),
.B(n_896),
.C(n_872),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1232),
.B(n_721),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1243),
.B(n_730),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1233),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1273),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1151),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1220),
.B(n_647),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1168),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1240),
.B(n_752),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1167),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1241),
.B(n_755),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1189),
.B(n_1136),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1138),
.B(n_766),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1148),
.B(n_985),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1172),
.B(n_1000),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1158),
.B(n_782),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1198),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1175),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1142),
.B(n_787),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1181),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1159),
.B(n_835),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1183),
.Y(n_1372)
);

BUFx5_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

OR2x6_ASAP7_75t_L g1374 ( 
.A(n_1144),
.B(n_1023),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1206),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1174),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1263),
.B(n_809),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1266),
.B(n_811),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1182),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1231),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1268),
.B(n_813),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1133),
.A2(n_689),
.B1(n_760),
.B2(n_658),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1237),
.B(n_815),
.Y(n_1383)
);

INVxp67_ASAP7_75t_SL g1384 ( 
.A(n_1279),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1255),
.B(n_816),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1218),
.B(n_818),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1142),
.B(n_1174),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1216),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1188),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_SL g1390 ( 
.A(n_1302),
.B(n_826),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1247),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1255),
.B(n_825),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1170),
.B(n_849),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1257),
.B(n_855),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1170),
.B(n_875),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1176),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1257),
.B(n_876),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1247),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1214),
.B(n_886),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1208),
.B(n_898),
.Y(n_1400)
);

AO221x1_ASAP7_75t_L g1401 ( 
.A1(n_1259),
.A2(n_1205),
.B1(n_1176),
.B2(n_1026),
.C(n_981),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1269),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1242),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1249),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1251),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1215),
.B(n_920),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1211),
.B(n_924),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1207),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1235),
.B(n_944),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1213),
.B(n_953),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1228),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_SL g1412 ( 
.A(n_1274),
.B(n_689),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1236),
.B(n_968),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1239),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1245),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1154),
.B(n_986),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1258),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1156),
.B(n_1012),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1276),
.Y(n_1419)
);

INVxp67_ASAP7_75t_L g1420 ( 
.A(n_1231),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1286),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1296),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1202),
.B(n_1025),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1217),
.A2(n_774),
.B1(n_792),
.B2(n_760),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1278),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1203),
.B(n_649),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1161),
.B(n_679),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1164),
.B(n_682),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1258),
.Y(n_1429)
);

NOR3xp33_ASAP7_75t_L g1430 ( 
.A(n_1219),
.B(n_1180),
.C(n_1179),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1166),
.B(n_650),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1288),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1204),
.B(n_655),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1196),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1171),
.B(n_684),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1210),
.B(n_694),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1163),
.B(n_1019),
.Y(n_1437)
);

NOR3xp33_ASAP7_75t_L g1438 ( 
.A(n_1184),
.B(n_657),
.C(n_656),
.Y(n_1438)
);

NAND2xp33_ASAP7_75t_L g1439 ( 
.A(n_1274),
.B(n_907),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1212),
.B(n_659),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1264),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1264),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1197),
.B(n_660),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1283),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1265),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1197),
.B(n_715),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1153),
.Y(n_1447)
);

NOR2xp67_ASAP7_75t_L g1448 ( 
.A(n_1196),
.B(n_484),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1287),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1265),
.B(n_661),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1304),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1309),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1152),
.B(n_728),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1262),
.B(n_665),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1254),
.Y(n_1455)
);

NOR2xp67_ASAP7_75t_L g1456 ( 
.A(n_1256),
.B(n_488),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1143),
.B(n_687),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1259),
.B(n_737),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1279),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1253),
.B(n_690),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1260),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1147),
.B(n_692),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1267),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1301),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1289),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1295),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1291),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1292),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1308),
.B(n_745),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1294),
.B(n_693),
.Y(n_1470)
);

INVxp33_ASAP7_75t_L g1471 ( 
.A(n_1169),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1295),
.Y(n_1472)
);

AND2x2_ASAP7_75t_SL g1473 ( 
.A(n_1137),
.B(n_774),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1297),
.B(n_696),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1299),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1305),
.B(n_747),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_SL g1477 ( 
.A(n_1139),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1306),
.B(n_701),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1277),
.Y(n_1479)
);

NOR2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1480)
);

NAND2xp33_ASAP7_75t_L g1481 ( 
.A(n_1222),
.B(n_907),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1285),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1290),
.B(n_702),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1298),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1304),
.B(n_750),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1275),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1280),
.Y(n_1487)
);

AND2x2_ASAP7_75t_SL g1488 ( 
.A(n_1298),
.B(n_792),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1284),
.A2(n_644),
.B1(n_645),
.B2(n_643),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1222),
.B(n_708),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1307),
.B(n_761),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1227),
.B(n_713),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1272),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1227),
.B(n_714),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1282),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1307),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_SL g1497 ( 
.A(n_1134),
.Y(n_1497)
);

NOR3xp33_ASAP7_75t_L g1498 ( 
.A(n_1293),
.B(n_726),
.C(n_723),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1300),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1303),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1134),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1134),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1134),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1194),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1194),
.B(n_772),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1194),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1209),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1209),
.B(n_779),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1238),
.B(n_733),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1238),
.B(n_734),
.Y(n_1510)
);

AND2x4_ASAP7_75t_SL g1511 ( 
.A(n_1270),
.B(n_883),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1270),
.Y(n_1512)
);

BUFx8_ASAP7_75t_L g1513 ( 
.A(n_1270),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1187),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1201),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1222),
.B(n_842),
.C(n_807),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1201),
.B(n_735),
.Y(n_1517)
);

AO221x1_ASAP7_75t_L g1518 ( 
.A1(n_1192),
.A2(n_1026),
.B1(n_981),
.B2(n_969),
.C(n_940),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1187),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1248),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1201),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1187),
.B(n_736),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1201),
.B(n_739),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1201),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1224),
.B(n_844),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1224),
.B(n_848),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1224),
.B(n_854),
.Y(n_1527)
);

NOR3xp33_ASAP7_75t_L g1528 ( 
.A(n_1177),
.B(n_742),
.C(n_741),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1201),
.B(n_744),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1135),
.B(n_858),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1248),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1224),
.B(n_860),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1201),
.B(n_748),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1201),
.Y(n_1534)
);

INVxp33_ASAP7_75t_L g1535 ( 
.A(n_1187),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1248),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1187),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1201),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1201),
.B(n_749),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1224),
.B(n_861),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1201),
.Y(n_1541)
);

BUFx5_ASAP7_75t_L g1542 ( 
.A(n_1273),
.Y(n_1542)
);

AND2x2_ASAP7_75t_SL g1543 ( 
.A(n_1177),
.B(n_883),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1201),
.B(n_753),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1187),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1201),
.B(n_754),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1248),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1187),
.B(n_759),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1224),
.B(n_866),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1224),
.B(n_869),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1225),
.B(n_874),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1177),
.B(n_1017),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1225),
.B(n_904),
.Y(n_1553)
);

NAND3xp33_ASAP7_75t_L g1554 ( 
.A(n_1222),
.B(n_926),
.C(n_917),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1248),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1201),
.B(n_763),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1201),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1248),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1135),
.B(n_939),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1201),
.B(n_764),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_L g1561 ( 
.A(n_1225),
.B(n_491),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1201),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1344),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1315),
.B(n_940),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1519),
.B(n_1537),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1516),
.A2(n_1003),
.B1(n_1020),
.B2(n_969),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1514),
.B(n_765),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1346),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1513),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1356),
.B(n_1020),
.Y(n_1570)
);

INVx5_ASAP7_75t_L g1571 ( 
.A(n_1402),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1373),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1535),
.B(n_1003),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1360),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1325),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1511),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1545),
.B(n_769),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1373),
.B(n_770),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1345),
.B(n_771),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1513),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1349),
.B(n_833),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1368),
.B(n_777),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1358),
.Y(n_1583)
);

INVxp33_ASAP7_75t_L g1584 ( 
.A(n_1552),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1316),
.B(n_778),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1316),
.B(n_788),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1311),
.B(n_1515),
.Y(n_1587)
);

AND2x6_ASAP7_75t_L g1588 ( 
.A(n_1345),
.B(n_956),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1481),
.A2(n_873),
.B1(n_877),
.B2(n_833),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1521),
.B(n_791),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1524),
.B(n_1534),
.Y(n_1591)
);

BUFx4f_ASAP7_75t_L g1592 ( 
.A(n_1343),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1538),
.A2(n_877),
.B1(n_880),
.B2(n_873),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1370),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1541),
.B(n_1557),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1345),
.B(n_793),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1367),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1562),
.B(n_796),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1331),
.B(n_797),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1355),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1374),
.B(n_851),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1354),
.B(n_1412),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1379),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1412),
.B(n_1402),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1362),
.B(n_880),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1367),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1367),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1389),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1403),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1516),
.A2(n_930),
.B1(n_973),
.B2(n_902),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1343),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1374),
.B(n_648),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1561),
.A2(n_653),
.B(n_663),
.C(n_651),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1391),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1341),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1342),
.B(n_902),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1551),
.B(n_798),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1551),
.B(n_802),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1382),
.A2(n_973),
.B1(n_983),
.B2(n_930),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1522),
.B(n_983),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1355),
.Y(n_1621)
);

BUFx8_ASAP7_75t_SL g1622 ( 
.A(n_1477),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1398),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1554),
.A2(n_994),
.B1(n_1009),
.B2(n_984),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1347),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1355),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1554),
.A2(n_994),
.B1(n_1009),
.B2(n_984),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1382),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1411),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1414),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1408),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1323),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1374),
.B(n_1317),
.Y(n_1633)
);

INVx6_ASAP7_75t_L g1634 ( 
.A(n_1343),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1334),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1336),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_R g1637 ( 
.A(n_1372),
.B(n_1014),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1553),
.B(n_812),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1404),
.Y(n_1639)
);

BUFx2_ASAP7_75t_SL g1640 ( 
.A(n_1477),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1490),
.A2(n_670),
.B1(n_683),
.B2(n_677),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1553),
.B(n_820),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1405),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1338),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1339),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1492),
.A2(n_704),
.B1(n_709),
.B2(n_685),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1402),
.B(n_822),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1494),
.A2(n_719),
.B1(n_720),
.B2(n_717),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1434),
.A2(n_963),
.B(n_961),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1375),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1447),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1388),
.Y(n_1652)
);

AND2x6_ASAP7_75t_SL g1653 ( 
.A(n_1453),
.B(n_810),
.Y(n_1653)
);

INVxp33_ASAP7_75t_SL g1654 ( 
.A(n_1424),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1432),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1417),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1363),
.B(n_824),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1429),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1509),
.A2(n_725),
.B1(n_727),
.B2(n_724),
.Y(n_1659)
);

OR2x6_ASAP7_75t_L g1660 ( 
.A(n_1415),
.B(n_691),
.Y(n_1660)
);

AO21x1_ASAP7_75t_L g1661 ( 
.A1(n_1439),
.A2(n_988),
.B(n_974),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1548),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_SL g1663 ( 
.A(n_1543),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1424),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1419),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1441),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1376),
.B(n_731),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1442),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1365),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1314),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1445),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1318),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1520),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1357),
.B(n_828),
.Y(n_1674)
);

INVx5_ASAP7_75t_L g1675 ( 
.A(n_1419),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1455),
.B(n_738),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1531),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1536),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1419),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1324),
.B(n_829),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_SL g1681 ( 
.A(n_1488),
.B(n_919),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1324),
.B(n_1312),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1547),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1313),
.B(n_831),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1348),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1517),
.B(n_832),
.Y(n_1686)
);

NOR2x2_ASAP7_75t_L g1687 ( 
.A(n_1473),
.B(n_1518),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1425),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1431),
.B(n_834),
.Y(n_1689)
);

INVx5_ASAP7_75t_L g1690 ( 
.A(n_1425),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1523),
.B(n_1529),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1425),
.B(n_837),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1510),
.A2(n_767),
.B1(n_768),
.B2(n_758),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1555),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1364),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1533),
.B(n_1539),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1380),
.B(n_776),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1544),
.B(n_838),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1558),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1457),
.Y(n_1700)
);

BUFx4f_ASAP7_75t_L g1701 ( 
.A(n_1396),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1335),
.A2(n_783),
.B1(n_789),
.B2(n_781),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1350),
.A2(n_795),
.B1(n_799),
.B2(n_790),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_SL g1704 ( 
.A(n_1351),
.B(n_845),
.C(n_840),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1462),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1383),
.B(n_846),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1480),
.Y(n_1707)
);

NOR3xp33_ASAP7_75t_SL g1708 ( 
.A(n_1353),
.B(n_853),
.C(n_850),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1321),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1546),
.B(n_856),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1444),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1420),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1330),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1333),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1498),
.A2(n_804),
.B1(n_806),
.B2(n_800),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1528),
.A2(n_819),
.B1(n_843),
.B2(n_808),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_SL g1717 ( 
.A(n_1393),
.B(n_871),
.C(n_870),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1556),
.B(n_878),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1337),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1560),
.B(n_879),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1463),
.A2(n_859),
.B1(n_862),
.B2(n_847),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1310),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1387),
.B(n_1525),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1450),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1386),
.B(n_885),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_SL g1726 ( 
.A(n_1390),
.B(n_1008),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1479),
.Y(n_1727)
);

BUFx12f_ASAP7_75t_SL g1728 ( 
.A(n_1444),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1444),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1446),
.A2(n_881),
.B1(n_882),
.B2(n_867),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1449),
.B(n_892),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1559),
.A2(n_887),
.B1(n_890),
.B2(n_884),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1449),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1465),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1465),
.B(n_894),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1526),
.B(n_891),
.Y(n_1736)
);

AO22x1_ASAP7_75t_L g1737 ( 
.A1(n_1471),
.A2(n_908),
.B1(n_909),
.B2(n_901),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1530),
.A2(n_899),
.B1(n_911),
.B2(n_893),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1327),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1468),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1366),
.B(n_1454),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1460),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1542),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1491),
.A2(n_913),
.B1(n_927),
.B2(n_912),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1468),
.B(n_918),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1329),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1421),
.Y(n_1747)
);

OR2x2_ASAP7_75t_SL g1748 ( 
.A(n_1401),
.B(n_992),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1527),
.B(n_933),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_R g1750 ( 
.A(n_1326),
.B(n_923),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1532),
.B(n_936),
.Y(n_1751)
);

AND2x2_ASAP7_75t_SL g1752 ( 
.A(n_1430),
.B(n_691),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1468),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1540),
.B(n_942),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1385),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1479),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1542),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1422),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1542),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1392),
.B(n_925),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1497),
.Y(n_1761)
);

INVxp67_ASAP7_75t_SL g1762 ( 
.A(n_1384),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1549),
.B(n_929),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1340),
.B(n_928),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1461),
.A2(n_1496),
.B1(n_1394),
.B2(n_1397),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1438),
.A2(n_948),
.B1(n_950),
.B2(n_947),
.Y(n_1766)
);

BUFx4f_ASAP7_75t_L g1767 ( 
.A(n_1371),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1377),
.A2(n_1028),
.B1(n_935),
.B2(n_937),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1483),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1322),
.B(n_1413),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1378),
.B(n_932),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1484),
.Y(n_1772)
);

CKINVDCx11_ASAP7_75t_R g1773 ( 
.A(n_1484),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1464),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1381),
.B(n_938),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1443),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1459),
.B(n_943),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1399),
.B(n_946),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1416),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1550),
.B(n_949),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1489),
.A2(n_955),
.B1(n_958),
.B2(n_951),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1452),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1406),
.B(n_952),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1418),
.B(n_954),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1466),
.B(n_957),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1352),
.B(n_959),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1437),
.B(n_964),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1409),
.B(n_1359),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1361),
.B(n_960),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1507),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1400),
.B(n_967),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1472),
.A2(n_965),
.B1(n_966),
.B2(n_962),
.Y(n_1792)
);

OR2x2_ASAP7_75t_SL g1793 ( 
.A(n_1426),
.B(n_976),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1427),
.B(n_971),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1507),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1497),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1467),
.B(n_972),
.Y(n_1797)
);

AO22x1_ASAP7_75t_L g1798 ( 
.A1(n_1428),
.A2(n_1435),
.B1(n_977),
.B2(n_979),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_R g1799 ( 
.A(n_1332),
.B(n_978),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1482),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1433),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1436),
.B(n_980),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1440),
.B(n_982),
.Y(n_1803)
);

XNOR2xp5_ASAP7_75t_L g1804 ( 
.A(n_1395),
.B(n_990),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1505),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1475),
.Y(n_1806)
);

OAI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1470),
.A2(n_1004),
.B1(n_1005),
.B2(n_993),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1474),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1485),
.A2(n_989),
.B1(n_991),
.B2(n_987),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1458),
.A2(n_1410),
.B1(n_1320),
.B2(n_1469),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1407),
.Y(n_1811)
);

BUFx5_ASAP7_75t_L g1812 ( 
.A(n_1503),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1478),
.Y(n_1813)
);

INVx5_ASAP7_75t_L g1814 ( 
.A(n_1451),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1423),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1319),
.B(n_999),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1328),
.B(n_1001),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1476),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1369),
.B(n_1007),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1508),
.Y(n_1820)
);

AND2x6_ASAP7_75t_L g1821 ( 
.A(n_1486),
.B(n_919),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1448),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1448),
.A2(n_1015),
.B1(n_1016),
.B2(n_1011),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1456),
.B(n_1018),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1456),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1451),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1487),
.B(n_699),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1495),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1502),
.B(n_698),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1499),
.B(n_934),
.Y(n_1830)
);

OR2x6_ASAP7_75t_L g1831 ( 
.A(n_1500),
.B(n_698),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1493),
.B(n_934),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1501),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1504),
.B(n_762),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1506),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1512),
.B(n_667),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1514),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1345),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1514),
.B(n_784),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1344),
.Y(n_1840)
);

BUFx4f_ASAP7_75t_L g1841 ( 
.A(n_1343),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1344),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1315),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1514),
.B(n_814),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1325),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1344),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1770),
.A2(n_852),
.B(n_817),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1654),
.A2(n_1793),
.B1(n_1664),
.B2(n_1628),
.Y(n_1848)
);

O2A1O1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1691),
.A2(n_817),
.B(n_868),
.C(n_814),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1741),
.A2(n_905),
.B(n_868),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1728),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1634),
.Y(n_1852)
);

A2O1A1Ixp33_ASAP7_75t_SL g1853 ( 
.A1(n_1696),
.A2(n_1710),
.B(n_1794),
.C(n_1580),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1655),
.B(n_905),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1563),
.Y(n_1855)
);

O2A1O1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1682),
.A2(n_916),
.B(n_921),
.C(n_914),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1568),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1566),
.A2(n_916),
.B1(n_921),
.B2(n_914),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1569),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1613),
.A2(n_1809),
.B(n_1662),
.C(n_1582),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1824),
.A2(n_1013),
.B(n_1072),
.Y(n_1861)
);

INVx5_ASAP7_75t_L g1862 ( 
.A(n_1569),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1616),
.A2(n_678),
.B1(n_823),
.B2(n_667),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1580),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1574),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1838),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1765),
.B(n_1091),
.C(n_1077),
.Y(n_1867)
);

AO32x1_ASAP7_75t_L g1868 ( 
.A1(n_1822),
.A2(n_1013),
.A3(n_1091),
.B1(n_1077),
.B2(n_836),
.Y(n_1868)
);

AOI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1825),
.A2(n_1077),
.B(n_823),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1843),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1814),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1584),
.B(n_10),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1605),
.B(n_10),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1573),
.B(n_11),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1594),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1582),
.A2(n_836),
.B(n_479),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1603),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1570),
.B(n_12),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1619),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.C(n_15),
.Y(n_1879)
);

A2O1A1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1776),
.A2(n_16),
.B(n_13),
.C(n_14),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1742),
.A2(n_480),
.B(n_477),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1587),
.B(n_16),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1724),
.A2(n_493),
.B(n_482),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1608),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1840),
.Y(n_1885)
);

INVx3_ASAP7_75t_SL g1886 ( 
.A(n_1634),
.Y(n_1886)
);

BUFx5_ASAP7_75t_L g1887 ( 
.A(n_1588),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1570),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1669),
.B(n_17),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1842),
.Y(n_1890)
);

A2O1A1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1813),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1591),
.B(n_20),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1622),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1809),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_1894)
);

O2A1O1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1627),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1814),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1592),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1564),
.B(n_1700),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1595),
.B(n_26),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1837),
.B(n_27),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1592),
.B(n_29),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1846),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1581),
.B(n_30),
.Y(n_1903)
);

O2A1O1Ixp5_ASAP7_75t_L g1904 ( 
.A1(n_1661),
.A2(n_498),
.B(n_501),
.C(n_496),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1841),
.B(n_30),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1578),
.A2(n_1760),
.B(n_1684),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1705),
.B(n_1722),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1565),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1617),
.A2(n_505),
.B(n_504),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1571),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1755),
.B(n_32),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1618),
.A2(n_509),
.B(n_507),
.Y(n_1912)
);

A2O1A1Ixp33_ASAP7_75t_L g1913 ( 
.A1(n_1823),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1627),
.B(n_35),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1814),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1841),
.B(n_36),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1620),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1566),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1918)
);

A2O1A1Ixp33_ASAP7_75t_SL g1919 ( 
.A1(n_1763),
.A2(n_1780),
.B(n_1649),
.C(n_1788),
.Y(n_1919)
);

BUFx2_ASAP7_75t_L g1920 ( 
.A(n_1615),
.Y(n_1920)
);

OAI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1702),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.C(n_43),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1739),
.B(n_44),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1831),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1637),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1638),
.A2(n_517),
.B(n_516),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1589),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1631),
.A2(n_1649),
.B(n_1629),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1642),
.B(n_49),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1641),
.B(n_50),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1637),
.Y(n_1930)
);

BUFx4_ASAP7_75t_SL g1931 ( 
.A(n_1651),
.Y(n_1931)
);

NOR2x1_ASAP7_75t_L g1932 ( 
.A(n_1640),
.B(n_50),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1571),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1639),
.Y(n_1934)
);

NAND3xp33_ASAP7_75t_SL g1935 ( 
.A(n_1681),
.B(n_51),
.C(n_52),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_SL g1936 ( 
.A(n_1681),
.B(n_1779),
.C(n_1750),
.Y(n_1936)
);

NOR3xp33_ASAP7_75t_SL g1937 ( 
.A(n_1707),
.B(n_53),
.C(n_54),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1600),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1831),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1643),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1646),
.B(n_55),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1743),
.A2(n_524),
.B(n_523),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1633),
.B(n_57),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1630),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1790),
.Y(n_1945)
);

A2O1A1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1823),
.A2(n_1769),
.B(n_1810),
.C(n_1746),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1609),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1757),
.A2(n_531),
.B(n_528),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1589),
.B(n_57),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1609),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_R g1951 ( 
.A(n_1712),
.B(n_58),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1633),
.B(n_58),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1571),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1648),
.B(n_59),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1659),
.B(n_59),
.Y(n_1955)
);

O2A1O1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1718),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1614),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1759),
.A2(n_536),
.B(n_532),
.Y(n_1958)
);

CKINVDCx20_ASAP7_75t_R g1959 ( 
.A(n_1583),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1693),
.B(n_63),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1833),
.A2(n_546),
.B(n_544),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_SL g1962 ( 
.A(n_1600),
.B(n_549),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1610),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1675),
.Y(n_1964)
);

NOR3xp33_ASAP7_75t_L g1965 ( 
.A(n_1704),
.B(n_1602),
.C(n_1798),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1621),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1811),
.B(n_66),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1660),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1811),
.B(n_67),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1583),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1623),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1835),
.A2(n_551),
.B(n_550),
.Y(n_1972)
);

INVx4_ASAP7_75t_L g1973 ( 
.A(n_1675),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1831),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1632),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1718),
.A2(n_556),
.B(n_555),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1621),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1808),
.B(n_1720),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1720),
.B(n_68),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1675),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1732),
.B(n_69),
.Y(n_1981)
);

O2A1O1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1604),
.A2(n_72),
.B(n_69),
.C(n_71),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1635),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1790),
.Y(n_1984)
);

NOR2x1_ASAP7_75t_R g1985 ( 
.A(n_1695),
.B(n_72),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1660),
.Y(n_1986)
);

INVx4_ASAP7_75t_L g1987 ( 
.A(n_1690),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1585),
.A2(n_558),
.B(n_557),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1660),
.Y(n_1989)
);

NAND2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1690),
.B(n_73),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1575),
.Y(n_1991)
);

BUFx4f_ASAP7_75t_L g1992 ( 
.A(n_1611),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1586),
.A2(n_560),
.B(n_559),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1644),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1663),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1995)
);

A2O1A1Ixp33_ASAP7_75t_L g1996 ( 
.A1(n_1709),
.A2(n_77),
.B(n_74),
.C(n_75),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1732),
.B(n_78),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1621),
.Y(n_1998)
);

AO21x1_ASAP7_75t_L g1999 ( 
.A1(n_1762),
.A2(n_564),
.B(n_562),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1834),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_2000)
);

A2O1A1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1713),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1690),
.B(n_83),
.Y(n_2002)
);

BUFx12f_ASAP7_75t_L g2003 ( 
.A(n_1845),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1761),
.B(n_84),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1799),
.B(n_1815),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1801),
.B(n_85),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1790),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1738),
.B(n_86),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1738),
.B(n_86),
.Y(n_2009)
);

BUFx3_ASAP7_75t_L g2010 ( 
.A(n_1665),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1679),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1636),
.Y(n_2012)
);

O2A1O1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_1674),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1663),
.A2(n_94),
.B1(n_90),
.B2(n_92),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1688),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1736),
.B(n_90),
.Y(n_2016)
);

AOI33xp33_ASAP7_75t_L g2017 ( 
.A1(n_1703),
.A2(n_96),
.A3(n_98),
.B1(n_92),
.B2(n_95),
.B3(n_97),
.Y(n_2017)
);

A2O1A1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1714),
.A2(n_99),
.B(n_95),
.C(n_96),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1761),
.B(n_101),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1834),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1689),
.B(n_102),
.Y(n_2021)
);

NAND3xp33_ASAP7_75t_SL g2022 ( 
.A(n_1716),
.B(n_103),
.C(n_104),
.Y(n_2022)
);

NOR3xp33_ASAP7_75t_SL g2023 ( 
.A(n_1726),
.B(n_104),
.C(n_106),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1736),
.B(n_108),
.Y(n_2024)
);

NAND3xp33_ASAP7_75t_SL g2025 ( 
.A(n_1766),
.B(n_108),
.C(n_109),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1834),
.A2(n_112),
.B1(n_109),
.B2(n_110),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_1796),
.B(n_110),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1729),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1749),
.B(n_1751),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1749),
.B(n_112),
.Y(n_2030)
);

BUFx6f_ASAP7_75t_L g2031 ( 
.A(n_1626),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1751),
.B(n_113),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1768),
.B(n_114),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1771),
.A2(n_579),
.B(n_574),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1650),
.Y(n_2035)
);

BUFx2_ASAP7_75t_L g2036 ( 
.A(n_1667),
.Y(n_2036)
);

OR2x6_ASAP7_75t_L g2037 ( 
.A(n_1576),
.B(n_114),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1588),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1839),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_2039)
);

NAND3xp33_ASAP7_75t_SL g2040 ( 
.A(n_1708),
.B(n_118),
.C(n_120),
.Y(n_2040)
);

INVx1_ASAP7_75t_SL g2041 ( 
.A(n_1588),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1625),
.B(n_121),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1775),
.A2(n_583),
.B(n_580),
.Y(n_2043)
);

O2A1O1Ixp33_ASAP7_75t_L g2044 ( 
.A1(n_1680),
.A2(n_1698),
.B(n_1686),
.C(n_1844),
.Y(n_2044)
);

NOR2x1p5_ASAP7_75t_L g2045 ( 
.A(n_1612),
.B(n_122),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1645),
.Y(n_2046)
);

OAI22x1_ASAP7_75t_L g2047 ( 
.A1(n_1612),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1652),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1774),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1624),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1577),
.B(n_125),
.Y(n_2051)
);

AND2x2_ASAP7_75t_SL g2052 ( 
.A(n_1593),
.B(n_1767),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1754),
.B(n_126),
.Y(n_2053)
);

O2A1O1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1802),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1828),
.A2(n_130),
.B1(n_127),
.B2(n_129),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1740),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1676),
.A2(n_133),
.B1(n_130),
.B2(n_131),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1719),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1753),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1747),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_1802),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1656),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_1786),
.A2(n_588),
.B(n_585),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_1803),
.B(n_1706),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1725),
.B(n_134),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1758),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1754),
.B(n_135),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1723),
.B(n_136),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1723),
.B(n_136),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1806),
.B(n_137),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1784),
.B(n_138),
.Y(n_2071)
);

OAI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1792),
.A2(n_1744),
.B1(n_1818),
.B2(n_1781),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1626),
.A2(n_590),
.B(n_589),
.Y(n_2073)
);

CKINVDCx20_ASAP7_75t_R g2074 ( 
.A(n_1773),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_1782),
.B(n_138),
.Y(n_2075)
);

BUFx10_ASAP7_75t_L g2076 ( 
.A(n_1588),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1658),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1781),
.B(n_139),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1626),
.A2(n_592),
.B(n_591),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1666),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1795),
.Y(n_2081)
);

NAND2xp33_ASAP7_75t_L g2082 ( 
.A(n_1821),
.B(n_593),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1730),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1807),
.B(n_144),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1567),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_1711),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_R g2087 ( 
.A(n_1767),
.B(n_145),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_SL g2088 ( 
.A(n_1717),
.B(n_146),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1821),
.Y(n_2089)
);

OAI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1730),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1676),
.B(n_148),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1789),
.B(n_150),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1701),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1670),
.Y(n_2094)
);

AOI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_1791),
.A2(n_606),
.B(n_605),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1697),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1657),
.A2(n_157),
.B1(n_154),
.B2(n_156),
.Y(n_2097)
);

INVx4_ASAP7_75t_L g2098 ( 
.A(n_1795),
.Y(n_2098)
);

AOI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_1789),
.A2(n_1697),
.B1(n_1816),
.B2(n_1601),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1817),
.B(n_158),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_L g2101 ( 
.A(n_1778),
.B(n_158),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1673),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1701),
.B(n_159),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1816),
.B(n_160),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1677),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_1734),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1590),
.B(n_161),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1678),
.Y(n_2108)
);

INVx4_ASAP7_75t_L g2109 ( 
.A(n_1727),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_1737),
.Y(n_2110)
);

BUFx12f_ASAP7_75t_L g2111 ( 
.A(n_1748),
.Y(n_2111)
);

OAI22x1_ASAP7_75t_L g2112 ( 
.A1(n_1601),
.A2(n_165),
.B1(n_162),
.B2(n_163),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1598),
.B(n_165),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_1653),
.Y(n_2114)
);

INVx4_ASAP7_75t_L g2115 ( 
.A(n_1727),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1721),
.B(n_166),
.Y(n_2116)
);

NAND3xp33_ASAP7_75t_L g2117 ( 
.A(n_1827),
.B(n_166),
.C(n_167),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1727),
.Y(n_2118)
);

A2O1A1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_1819),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1715),
.B(n_168),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1752),
.A2(n_175),
.B1(n_171),
.B2(n_172),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_1821),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1804),
.B(n_176),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_1821),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1699),
.Y(n_2125)
);

O2A1O1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_1783),
.A2(n_179),
.B(n_176),
.C(n_177),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_1733),
.Y(n_2127)
);

OAI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_1572),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1668),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_SL g2130 ( 
.A1(n_1687),
.A2(n_185),
.B1(n_182),
.B2(n_184),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1671),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1672),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1756),
.B(n_186),
.Y(n_2133)
);

OAI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_1772),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_1647),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1777),
.A2(n_619),
.B(n_617),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1787),
.B(n_189),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_1599),
.B(n_190),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1683),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1694),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1764),
.B(n_191),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1797),
.B(n_191),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1653),
.B(n_192),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1785),
.A2(n_626),
.B(n_620),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1829),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_1692),
.B(n_195),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1731),
.B(n_196),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_R g2148 ( 
.A(n_1756),
.B(n_196),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1820),
.A2(n_628),
.B(n_627),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1830),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1597),
.B(n_197),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1597),
.B(n_197),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1800),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1735),
.B(n_198),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1745),
.B(n_198),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_1606),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1579),
.B(n_199),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1832),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_1606),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1826),
.B(n_200),
.Y(n_2160)
);

OAI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1805),
.A2(n_201),
.B(n_202),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1596),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_1607),
.A2(n_205),
.B(n_202),
.C(n_204),
.Y(n_2163)
);

INVx2_ASAP7_75t_SL g2164 ( 
.A(n_1607),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1836),
.A2(n_631),
.B(n_630),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_1812),
.B(n_205),
.Y(n_2166)
);

NOR2x1_ASAP7_75t_L g2167 ( 
.A(n_1812),
.B(n_208),
.Y(n_2167)
);

OAI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_1812),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2168)
);

OAI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_1812),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1838),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_1584),
.B(n_212),
.Y(n_2171)
);

NAND2x1p5_ASAP7_75t_L g2172 ( 
.A(n_1571),
.B(n_212),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1655),
.B(n_213),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1843),
.B(n_213),
.Y(n_2174)
);

CKINVDCx20_ASAP7_75t_R g2175 ( 
.A(n_1622),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1655),
.B(n_214),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1563),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_1584),
.B(n_214),
.Y(n_2178)
);

AO32x1_ASAP7_75t_L g2179 ( 
.A1(n_1822),
.A2(n_216),
.A3(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1566),
.A2(n_219),
.B1(n_216),
.B2(n_217),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1843),
.B(n_221),
.Y(n_2181)
);

O2A1O1Ixp33_ASAP7_75t_L g2182 ( 
.A1(n_1691),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_1584),
.B(n_222),
.Y(n_2183)
);

INVx4_ASAP7_75t_L g2184 ( 
.A(n_1569),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1685),
.B(n_224),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_1728),
.Y(n_2186)
);

INVx4_ASAP7_75t_L g2187 ( 
.A(n_1569),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1563),
.Y(n_2188)
);

NAND3xp33_ASAP7_75t_SL g2189 ( 
.A(n_1681),
.B(n_228),
.C(n_229),
.Y(n_2189)
);

BUFx4f_ASAP7_75t_SL g2190 ( 
.A(n_1651),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1655),
.B(n_229),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1655),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1655),
.B(n_230),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1843),
.B(n_231),
.Y(n_2194)
);

O2A1O1Ixp33_ASAP7_75t_L g2195 ( 
.A1(n_1691),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1584),
.B(n_232),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_1570),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1655),
.B(n_234),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_1770),
.A2(n_637),
.B(n_635),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_SL g2200 ( 
.A1(n_1654),
.A2(n_239),
.B1(n_235),
.B2(n_236),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_1570),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1655),
.B(n_240),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1843),
.B(n_241),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1655),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1655),
.Y(n_2205)
);

O2A1O1Ixp33_ASAP7_75t_L g2206 ( 
.A1(n_1691),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1563),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1655),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1655),
.B(n_248),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1584),
.B(n_249),
.Y(n_2210)
);

O2A1O1Ixp33_ASAP7_75t_L g2211 ( 
.A1(n_1691),
.A2(n_250),
.B(n_251),
.C(n_252),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1655),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1655),
.B(n_251),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1838),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1685),
.B(n_252),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_1728),
.Y(n_2216)
);

O2A1O1Ixp33_ASAP7_75t_L g2217 ( 
.A1(n_1691),
.A2(n_253),
.B(n_254),
.C(n_255),
.Y(n_2217)
);

OAI21xp33_ASAP7_75t_L g2218 ( 
.A1(n_1696),
.A2(n_258),
.B(n_259),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1569),
.Y(n_2219)
);

AND2x4_ASAP7_75t_L g2220 ( 
.A(n_1655),
.B(n_258),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1655),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_1728),
.Y(n_2222)
);

OAI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_1823),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_2223)
);

OAI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_1682),
.A2(n_263),
.B(n_264),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1570),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_2225)
);

A2O1A1Ixp33_ASAP7_75t_L g2226 ( 
.A1(n_1696),
.A2(n_265),
.B(n_266),
.C(n_267),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1843),
.B(n_268),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1655),
.B(n_269),
.Y(n_2228)
);

NAND2x1_ASAP7_75t_L g2229 ( 
.A(n_1588),
.B(n_270),
.Y(n_2229)
);

OR2x6_ASAP7_75t_L g2230 ( 
.A(n_1634),
.B(n_461),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1843),
.B(n_270),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_1770),
.A2(n_271),
.B(n_272),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1584),
.B(n_271),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1655),
.B(n_272),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1569),
.Y(n_2235)
);

BUFx8_ASAP7_75t_L g2236 ( 
.A(n_1663),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1843),
.B(n_273),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1655),
.B(n_273),
.Y(n_2238)
);

INVx1_ASAP7_75t_SL g2239 ( 
.A(n_1634),
.Y(n_2239)
);

AOI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_1566),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_2240)
);

NAND2x1p5_ASAP7_75t_L g2241 ( 
.A(n_1571),
.B(n_274),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1655),
.B(n_277),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_1634),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_1570),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1634),
.Y(n_2245)
);

AOI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_1770),
.A2(n_279),
.B(n_280),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1655),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1843),
.B(n_281),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1622),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1655),
.B(n_281),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1843),
.B(n_283),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1838),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2192),
.Y(n_2253)
);

BUFx3_ASAP7_75t_L g2254 ( 
.A(n_1886),
.Y(n_2254)
);

OA21x2_ASAP7_75t_L g2255 ( 
.A1(n_1867),
.A2(n_283),
.B(n_284),
.Y(n_2255)
);

BUFx2_ASAP7_75t_L g2256 ( 
.A(n_1959),
.Y(n_2256)
);

NAND2x1p5_ASAP7_75t_L g2257 ( 
.A(n_1973),
.B(n_284),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_2098),
.Y(n_2258)
);

NAND2x1p5_ASAP7_75t_L g2259 ( 
.A(n_1973),
.B(n_285),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1946),
.B(n_1927),
.Y(n_2260)
);

OA21x2_ASAP7_75t_L g2261 ( 
.A1(n_1867),
.A2(n_1999),
.B(n_1904),
.Y(n_2261)
);

INVx1_ASAP7_75t_SL g2262 ( 
.A(n_1870),
.Y(n_2262)
);

OAI21x1_ASAP7_75t_SL g2263 ( 
.A1(n_1927),
.A2(n_285),
.B(n_286),
.Y(n_2263)
);

BUFx5_ASAP7_75t_L g2264 ( 
.A(n_2076),
.Y(n_2264)
);

INVx4_ASAP7_75t_L g2265 ( 
.A(n_2230),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2204),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2205),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2029),
.B(n_1978),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2208),
.Y(n_2269)
);

BUFx12f_ASAP7_75t_L g2270 ( 
.A(n_1893),
.Y(n_2270)
);

NAND2x1p5_ASAP7_75t_L g2271 ( 
.A(n_1987),
.B(n_288),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_1970),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1855),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1875),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1907),
.B(n_289),
.Y(n_2275)
);

NOR2x1_ASAP7_75t_R g2276 ( 
.A(n_2249),
.B(n_290),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2212),
.B(n_290),
.Y(n_2277)
);

HB1xp67_ASAP7_75t_L g2278 ( 
.A(n_2230),
.Y(n_2278)
);

BUFx2_ASAP7_75t_R g2279 ( 
.A(n_2114),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1884),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2044),
.A2(n_291),
.B(n_292),
.Y(n_2281)
);

OR2x6_ASAP7_75t_L g2282 ( 
.A(n_2230),
.B(n_295),
.Y(n_2282)
);

BUFx3_ASAP7_75t_L g2283 ( 
.A(n_1851),
.Y(n_2283)
);

AOI22x1_ASAP7_75t_L g2284 ( 
.A1(n_1876),
.A2(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_2284)
);

INVx1_ASAP7_75t_SL g2285 ( 
.A(n_2222),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_2003),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2064),
.B(n_299),
.Y(n_2287)
);

OA21x2_ASAP7_75t_L g2288 ( 
.A1(n_2161),
.A2(n_299),
.B(n_301),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2177),
.B(n_302),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_2245),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2221),
.Y(n_2291)
);

NAND2x1_ASAP7_75t_L g2292 ( 
.A(n_2109),
.B(n_302),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_1906),
.A2(n_303),
.B(n_304),
.Y(n_2293)
);

INVx2_ASAP7_75t_SL g2294 ( 
.A(n_1992),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_2036),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2188),
.Y(n_2296)
);

NAND2x1p5_ASAP7_75t_L g2297 ( 
.A(n_1987),
.B(n_305),
.Y(n_2297)
);

INVxp67_ASAP7_75t_SL g2298 ( 
.A(n_2075),
.Y(n_2298)
);

BUFx8_ASAP7_75t_L g2299 ( 
.A(n_1920),
.Y(n_2299)
);

BUFx3_ASAP7_75t_L g2300 ( 
.A(n_1991),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2247),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2207),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1857),
.Y(n_2303)
);

AO21x2_ASAP7_75t_L g2304 ( 
.A1(n_2224),
.A2(n_312),
.B(n_313),
.Y(n_2304)
);

AO21x2_ASAP7_75t_L g2305 ( 
.A1(n_2224),
.A2(n_312),
.B(n_315),
.Y(n_2305)
);

BUFx5_ASAP7_75t_L g2306 ( 
.A(n_1934),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_1897),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_1861),
.A2(n_315),
.B(n_317),
.Y(n_2308)
);

BUFx2_ASAP7_75t_SL g2309 ( 
.A(n_2175),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1865),
.Y(n_2310)
);

BUFx2_ASAP7_75t_R g2311 ( 
.A(n_2005),
.Y(n_2311)
);

BUFx12f_ASAP7_75t_L g2312 ( 
.A(n_2236),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2099),
.B(n_319),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_1887),
.B(n_319),
.Y(n_2314)
);

BUFx10_ASAP7_75t_L g2315 ( 
.A(n_2070),
.Y(n_2315)
);

OA21x2_ASAP7_75t_L g2316 ( 
.A1(n_2161),
.A2(n_320),
.B(n_321),
.Y(n_2316)
);

OAI21x1_ASAP7_75t_SL g2317 ( 
.A1(n_2167),
.A2(n_322),
.B(n_324),
.Y(n_2317)
);

BUFx2_ASAP7_75t_L g2318 ( 
.A(n_2186),
.Y(n_2318)
);

INVx1_ASAP7_75t_SL g2319 ( 
.A(n_2216),
.Y(n_2319)
);

AOI21xp5_ASAP7_75t_L g2320 ( 
.A1(n_1919),
.A2(n_322),
.B(n_324),
.Y(n_2320)
);

BUFx2_ASAP7_75t_L g2321 ( 
.A(n_2087),
.Y(n_2321)
);

INVxp33_ASAP7_75t_L g2322 ( 
.A(n_1898),
.Y(n_2322)
);

NAND2x1p5_ASAP7_75t_L g2323 ( 
.A(n_2098),
.B(n_326),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_1949),
.B(n_327),
.Y(n_2324)
);

BUFx3_ASAP7_75t_L g2325 ( 
.A(n_1871),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1877),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1885),
.Y(n_2327)
);

AO21x2_ASAP7_75t_L g2328 ( 
.A1(n_2218),
.A2(n_327),
.B(n_328),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1890),
.Y(n_2329)
);

AOI22x1_ASAP7_75t_L g2330 ( 
.A1(n_1976),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_2330)
);

INVx4_ASAP7_75t_L g2331 ( 
.A(n_1862),
.Y(n_2331)
);

INVx4_ASAP7_75t_L g2332 ( 
.A(n_1862),
.Y(n_2332)
);

AO21x2_ASAP7_75t_L g2333 ( 
.A1(n_1869),
.A2(n_329),
.B(n_330),
.Y(n_2333)
);

INVx4_ASAP7_75t_L g2334 ( 
.A(n_1862),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_1871),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_1896),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1994),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1902),
.Y(n_2338)
);

AO21x2_ASAP7_75t_L g2339 ( 
.A1(n_1935),
.A2(n_335),
.B(n_336),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2035),
.Y(n_2340)
);

BUFx12f_ASAP7_75t_L g2341 ( 
.A(n_2236),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_1938),
.Y(n_2342)
);

BUFx12f_ASAP7_75t_L g2343 ( 
.A(n_2111),
.Y(n_2343)
);

AOI22x1_ASAP7_75t_L g2344 ( 
.A1(n_2034),
.A2(n_337),
.B1(n_340),
.B2(n_341),
.Y(n_2344)
);

INVx3_ASAP7_75t_SL g2345 ( 
.A(n_2239),
.Y(n_2345)
);

AOI22x1_ASAP7_75t_L g2346 ( 
.A1(n_2043),
.A2(n_337),
.B1(n_340),
.B2(n_342),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_1896),
.Y(n_2347)
);

OR2x6_ASAP7_75t_L g2348 ( 
.A(n_2070),
.B(n_343),
.Y(n_2348)
);

OAI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_1860),
.A2(n_343),
.B(n_344),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1938),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1957),
.B(n_1971),
.Y(n_2351)
);

INVx2_ASAP7_75t_SL g2352 ( 
.A(n_1992),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2075),
.Y(n_2353)
);

BUFx3_ASAP7_75t_L g2354 ( 
.A(n_1915),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_1915),
.Y(n_2355)
);

INVx5_ASAP7_75t_L g2356 ( 
.A(n_1966),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2109),
.Y(n_2357)
);

INVx4_ASAP7_75t_L g2358 ( 
.A(n_2190),
.Y(n_2358)
);

BUFx2_ASAP7_75t_L g2359 ( 
.A(n_1968),
.Y(n_2359)
);

INVx1_ASAP7_75t_SL g2360 ( 
.A(n_2015),
.Y(n_2360)
);

BUFx4f_ASAP7_75t_L g2361 ( 
.A(n_2037),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1944),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2010),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2185),
.B(n_344),
.Y(n_2364)
);

AO21x2_ASAP7_75t_L g2365 ( 
.A1(n_2189),
.A2(n_345),
.B(n_347),
.Y(n_2365)
);

BUFx12f_ASAP7_75t_L g2366 ( 
.A(n_2045),
.Y(n_2366)
);

INVx3_ASAP7_75t_L g2367 ( 
.A(n_2115),
.Y(n_2367)
);

BUFx12f_ASAP7_75t_L g2368 ( 
.A(n_1852),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1975),
.Y(n_2369)
);

BUFx12f_ASAP7_75t_L g2370 ( 
.A(n_2243),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_1868),
.A2(n_345),
.B(n_347),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2028),
.Y(n_2372)
);

INVx3_ASAP7_75t_L g2373 ( 
.A(n_2115),
.Y(n_2373)
);

OAI21x1_ASAP7_75t_L g2374 ( 
.A1(n_2199),
.A2(n_348),
.B(n_349),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_1848),
.B(n_349),
.Y(n_2375)
);

BUFx12f_ASAP7_75t_SL g2376 ( 
.A(n_2037),
.Y(n_2376)
);

BUFx12f_ASAP7_75t_L g2377 ( 
.A(n_2037),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_1931),
.Y(n_2378)
);

BUFx2_ASAP7_75t_SL g2379 ( 
.A(n_2074),
.Y(n_2379)
);

INVx5_ASAP7_75t_L g2380 ( 
.A(n_1966),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1983),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_SL g2382 ( 
.A1(n_2000),
.A2(n_351),
.B(n_352),
.Y(n_2382)
);

NAND2x1p5_ASAP7_75t_L g2383 ( 
.A(n_2038),
.B(n_353),
.Y(n_2383)
);

BUFx3_ASAP7_75t_L g2384 ( 
.A(n_1964),
.Y(n_2384)
);

BUFx3_ASAP7_75t_L g2385 ( 
.A(n_2127),
.Y(n_2385)
);

HB1xp67_ASAP7_75t_L g2386 ( 
.A(n_2198),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1977),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2012),
.B(n_359),
.Y(n_2388)
);

BUFx4f_ASAP7_75t_L g2389 ( 
.A(n_1990),
.Y(n_2389)
);

BUFx2_ASAP7_75t_R g2390 ( 
.A(n_2143),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1977),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1977),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_1986),
.Y(n_2393)
);

OAI21x1_ASAP7_75t_L g2394 ( 
.A1(n_1942),
.A2(n_1958),
.B(n_1948),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2046),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1998),
.Y(n_2396)
);

OAI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_1979),
.A2(n_361),
.B(n_362),
.Y(n_2397)
);

CKINVDCx14_ASAP7_75t_R g2398 ( 
.A(n_2148),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2048),
.B(n_363),
.Y(n_2399)
);

AOI22x1_ASAP7_75t_L g2400 ( 
.A1(n_2063),
.A2(n_363),
.B1(n_364),
.B2(n_366),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2058),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2215),
.B(n_2123),
.Y(n_2402)
);

AO21x2_ASAP7_75t_L g2403 ( 
.A1(n_2166),
.A2(n_366),
.B(n_368),
.Y(n_2403)
);

AOI21x1_ASAP7_75t_L g2404 ( 
.A1(n_2133),
.A2(n_372),
.B(n_373),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_1974),
.B(n_372),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_1998),
.Y(n_2406)
);

BUFx12f_ASAP7_75t_L g2407 ( 
.A(n_1989),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2049),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_1856),
.A2(n_376),
.B(n_377),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_1974),
.B(n_378),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_1998),
.Y(n_2411)
);

BUFx12f_ASAP7_75t_L g2412 ( 
.A(n_2052),
.Y(n_2412)
);

INVx5_ASAP7_75t_L g2413 ( 
.A(n_2031),
.Y(n_2413)
);

OR2x6_ASAP7_75t_SL g2414 ( 
.A(n_1914),
.B(n_378),
.Y(n_2414)
);

AO21x2_ASAP7_75t_L g2415 ( 
.A1(n_1850),
.A2(n_379),
.B(n_380),
.Y(n_2415)
);

INVx5_ASAP7_75t_SL g2416 ( 
.A(n_2198),
.Y(n_2416)
);

BUFx12f_ASAP7_75t_L g2417 ( 
.A(n_2093),
.Y(n_2417)
);

INVx6_ASAP7_75t_L g2418 ( 
.A(n_2184),
.Y(n_2418)
);

BUFx2_ASAP7_75t_R g2419 ( 
.A(n_1901),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2031),
.Y(n_2420)
);

OAI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_1849),
.A2(n_379),
.B(n_382),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2094),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2072),
.B(n_382),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2031),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_1910),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2102),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_SL g2427 ( 
.A(n_1985),
.B(n_384),
.Y(n_2427)
);

INVxp67_ASAP7_75t_L g2428 ( 
.A(n_2220),
.Y(n_2428)
);

OR3x4_ASAP7_75t_SL g2429 ( 
.A(n_2130),
.B(n_384),
.C(n_385),
.Y(n_2429)
);

INVx5_ASAP7_75t_L g2430 ( 
.A(n_1866),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_1945),
.Y(n_2431)
);

AO21x2_ASAP7_75t_L g2432 ( 
.A1(n_1847),
.A2(n_385),
.B(n_389),
.Y(n_2432)
);

OAI21x1_ASAP7_75t_SL g2433 ( 
.A1(n_2000),
.A2(n_389),
.B(n_390),
.Y(n_2433)
);

AOI22x1_ASAP7_75t_L g2434 ( 
.A1(n_1988),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_2434)
);

OAI21x1_ASAP7_75t_L g2435 ( 
.A1(n_1993),
.A2(n_391),
.B(n_392),
.Y(n_2435)
);

OAI21x1_ASAP7_75t_L g2436 ( 
.A1(n_1909),
.A2(n_393),
.B(n_394),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1940),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_1933),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2062),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2105),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_1990),
.Y(n_2441)
);

BUFx12f_ASAP7_75t_L g2442 ( 
.A(n_2184),
.Y(n_2442)
);

AO21x2_ASAP7_75t_L g2443 ( 
.A1(n_1912),
.A2(n_393),
.B(n_394),
.Y(n_2443)
);

INVx3_ASAP7_75t_L g2444 ( 
.A(n_1945),
.Y(n_2444)
);

OR2x6_ASAP7_75t_L g2445 ( 
.A(n_2220),
.B(n_395),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2108),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_1984),
.Y(n_2447)
);

INVx6_ASAP7_75t_L g2448 ( 
.A(n_2187),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2073),
.A2(n_397),
.B(n_398),
.Y(n_2449)
);

CKINVDCx20_ASAP7_75t_R g2450 ( 
.A(n_1924),
.Y(n_2450)
);

NAND2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2041),
.B(n_397),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2125),
.Y(n_2452)
);

INVx4_ASAP7_75t_L g2453 ( 
.A(n_2172),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2015),
.Y(n_2454)
);

INVx3_ASAP7_75t_L g2455 ( 
.A(n_1984),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2056),
.B(n_399),
.Y(n_2456)
);

OAI21x1_ASAP7_75t_SL g2457 ( 
.A1(n_2223),
.A2(n_2090),
.B(n_2083),
.Y(n_2457)
);

AND2x4_ASAP7_75t_L g2458 ( 
.A(n_1947),
.B(n_400),
.Y(n_2458)
);

INVx1_ASAP7_75t_SL g2459 ( 
.A(n_2239),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2060),
.Y(n_2460)
);

OAI21x1_ASAP7_75t_L g2461 ( 
.A1(n_2079),
.A2(n_400),
.B(n_401),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2059),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2007),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_SL g2464 ( 
.A(n_2187),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2021),
.B(n_405),
.Y(n_2465)
);

INVxp67_ASAP7_75t_SL g2466 ( 
.A(n_2252),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_1922),
.B(n_406),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2066),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2017),
.Y(n_2469)
);

OAI21x1_ASAP7_75t_L g2470 ( 
.A1(n_1925),
.A2(n_406),
.B(n_407),
.Y(n_2470)
);

OA21x2_ASAP7_75t_L g2471 ( 
.A1(n_1881),
.A2(n_1883),
.B(n_1961),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2081),
.Y(n_2472)
);

OAI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_1882),
.A2(n_407),
.B(n_408),
.Y(n_2473)
);

CKINVDCx16_ASAP7_75t_R g2474 ( 
.A(n_1951),
.Y(n_2474)
);

INVx3_ASAP7_75t_L g2475 ( 
.A(n_2081),
.Y(n_2475)
);

INVxp33_ASAP7_75t_L g2476 ( 
.A(n_1848),
.Y(n_2476)
);

AOI22x1_ASAP7_75t_L g2477 ( 
.A1(n_2095),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2173),
.Y(n_2478)
);

CKINVDCx14_ASAP7_75t_R g2479 ( 
.A(n_1936),
.Y(n_2479)
);

NAND2x1_ASAP7_75t_L g2480 ( 
.A(n_2118),
.B(n_409),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_1889),
.B(n_2065),
.Y(n_2481)
);

OA21x2_ASAP7_75t_L g2482 ( 
.A1(n_1972),
.A2(n_411),
.B(n_413),
.Y(n_2482)
);

INVx3_ASAP7_75t_L g2483 ( 
.A(n_2252),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_1953),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2176),
.Y(n_2485)
);

AND2x4_ASAP7_75t_L g2486 ( 
.A(n_1950),
.B(n_461),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_1980),
.Y(n_2487)
);

AOI22x1_ASAP7_75t_L g2488 ( 
.A1(n_2136),
.A2(n_415),
.B1(n_417),
.B2(n_418),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2129),
.B(n_417),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_1868),
.A2(n_419),
.B(n_420),
.Y(n_2490)
);

OAI21x1_ASAP7_75t_L g2491 ( 
.A1(n_2149),
.A2(n_2156),
.B(n_2144),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2071),
.B(n_419),
.Y(n_2492)
);

NAND2x1_ASAP7_75t_L g2493 ( 
.A(n_2252),
.B(n_420),
.Y(n_2493)
);

AND2x6_ASAP7_75t_L g2494 ( 
.A(n_2041),
.B(n_421),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_1911),
.B(n_422),
.Y(n_2495)
);

OAI21x1_ASAP7_75t_L g2496 ( 
.A1(n_2172),
.A2(n_423),
.B(n_424),
.Y(n_2496)
);

OAI21x1_ASAP7_75t_L g2497 ( 
.A1(n_2156),
.A2(n_423),
.B(n_424),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2077),
.Y(n_2498)
);

OAI21x1_ASAP7_75t_L g2499 ( 
.A1(n_2165),
.A2(n_425),
.B(n_426),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_1908),
.B(n_425),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2080),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_2011),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_SL g2503 ( 
.A(n_2135),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2191),
.Y(n_2504)
);

NAND2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2089),
.B(n_426),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2193),
.Y(n_2506)
);

INVx5_ASAP7_75t_L g2507 ( 
.A(n_2170),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2241),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_1858),
.B(n_427),
.Y(n_2509)
);

OAI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2241),
.A2(n_427),
.B(n_428),
.Y(n_2510)
);

AO21x2_ASAP7_75t_L g2511 ( 
.A1(n_1928),
.A2(n_430),
.B(n_431),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2131),
.Y(n_2512)
);

NAND2x1p5_ASAP7_75t_L g2513 ( 
.A(n_2122),
.B(n_430),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_1873),
.B(n_431),
.Y(n_2514)
);

OAI21x1_ASAP7_75t_L g2515 ( 
.A1(n_1982),
.A2(n_432),
.B(n_433),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2139),
.Y(n_2516)
);

BUFx4f_ASAP7_75t_SL g2517 ( 
.A(n_1859),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2202),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_1878),
.B(n_2091),
.Y(n_2519)
);

CKINVDCx20_ASAP7_75t_R g2520 ( 
.A(n_1930),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2132),
.B(n_432),
.Y(n_2521)
);

BUFx2_ASAP7_75t_L g2522 ( 
.A(n_2110),
.Y(n_2522)
);

AO21x2_ASAP7_75t_L g2523 ( 
.A1(n_2025),
.A2(n_434),
.B(n_435),
.Y(n_2523)
);

NAND2x1p5_ASAP7_75t_L g2524 ( 
.A(n_2124),
.B(n_434),
.Y(n_2524)
);

INVx2_ASAP7_75t_SL g2525 ( 
.A(n_1859),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2214),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2209),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_1872),
.B(n_437),
.Y(n_2528)
);

NOR2x1_ASAP7_75t_R g2529 ( 
.A(n_1887),
.B(n_437),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2213),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2228),
.Y(n_2531)
);

INVx1_ASAP7_75t_SL g2532 ( 
.A(n_1864),
.Y(n_2532)
);

BUFx4f_ASAP7_75t_L g2533 ( 
.A(n_2004),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2234),
.Y(n_2534)
);

CKINVDCx16_ASAP7_75t_R g2535 ( 
.A(n_2200),
.Y(n_2535)
);

AND2x6_ASAP7_75t_L g2536 ( 
.A(n_2214),
.B(n_438),
.Y(n_2536)
);

BUFx12f_ASAP7_75t_L g2537 ( 
.A(n_2004),
.Y(n_2537)
);

OAI21x1_ASAP7_75t_SL g2538 ( 
.A1(n_2223),
.A2(n_439),
.B(n_440),
.Y(n_2538)
);

OR2x6_ASAP7_75t_L g2539 ( 
.A(n_2229),
.B(n_439),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2171),
.B(n_440),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2238),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2100),
.B(n_441),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_1887),
.Y(n_2543)
);

AO21x2_ASAP7_75t_L g2544 ( 
.A1(n_2232),
.A2(n_441),
.B(n_442),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2140),
.B(n_442),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2178),
.B(n_443),
.Y(n_2546)
);

AO21x2_ASAP7_75t_L g2547 ( 
.A1(n_2246),
.A2(n_443),
.B(n_444),
.Y(n_2547)
);

OAI21x1_ASAP7_75t_L g2548 ( 
.A1(n_2151),
.A2(n_444),
.B(n_445),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_1864),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2214),
.Y(n_2550)
);

AO21x2_ASAP7_75t_L g2551 ( 
.A1(n_2022),
.A2(n_2082),
.B(n_2107),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2162),
.B(n_2219),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_2219),
.Y(n_2553)
);

OAI21x1_ASAP7_75t_L g2554 ( 
.A1(n_2152),
.A2(n_446),
.B(n_447),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_1892),
.B(n_448),
.Y(n_2555)
);

OAI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_1899),
.A2(n_448),
.B(n_449),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2130),
.Y(n_2557)
);

OR2x6_ASAP7_75t_L g2558 ( 
.A(n_2200),
.B(n_449),
.Y(n_2558)
);

BUFx2_ASAP7_75t_SL g2559 ( 
.A(n_1887),
.Y(n_2559)
);

INVx3_ASAP7_75t_SL g2560 ( 
.A(n_2235),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2235),
.Y(n_2561)
);

AO21x1_ASAP7_75t_L g2562 ( 
.A1(n_2054),
.A2(n_450),
.B(n_454),
.Y(n_2562)
);

INVxp67_ASAP7_75t_L g2563 ( 
.A(n_2016),
.Y(n_2563)
);

INVx4_ASAP7_75t_L g2564 ( 
.A(n_2159),
.Y(n_2564)
);

BUFx10_ASAP7_75t_L g2565 ( 
.A(n_1952),
.Y(n_2565)
);

INVx5_ASAP7_75t_SL g2566 ( 
.A(n_2159),
.Y(n_2566)
);

BUFx2_ASAP7_75t_SL g2567 ( 
.A(n_2086),
.Y(n_2567)
);

AND2x4_ASAP7_75t_L g2568 ( 
.A(n_2153),
.B(n_460),
.Y(n_2568)
);

OAI21x1_ASAP7_75t_L g2569 ( 
.A1(n_2002),
.A2(n_454),
.B(n_455),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2242),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2106),
.Y(n_2571)
);

BUFx3_ASAP7_75t_L g2572 ( 
.A(n_2164),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2250),
.Y(n_2573)
);

AOI22x1_ASAP7_75t_L g2574 ( 
.A1(n_2047),
.A2(n_458),
.B1(n_455),
.B2(n_456),
.Y(n_2574)
);

BUFx3_ASAP7_75t_L g2575 ( 
.A(n_2160),
.Y(n_2575)
);

INVx3_ASAP7_75t_SL g2576 ( 
.A(n_1905),
.Y(n_2576)
);

BUFx2_ASAP7_75t_L g2577 ( 
.A(n_2088),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2138),
.Y(n_2578)
);

OAI21x1_ASAP7_75t_L g2579 ( 
.A1(n_1854),
.A2(n_2158),
.B(n_2150),
.Y(n_2579)
);

OAI21x1_ASAP7_75t_L g2580 ( 
.A1(n_2113),
.A2(n_1956),
.B(n_2182),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2183),
.B(n_2196),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_1853),
.B(n_2101),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_1868),
.Y(n_2583)
);

INVx3_ASAP7_75t_L g2584 ( 
.A(n_2154),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2273),
.Y(n_2585)
);

INVx6_ASAP7_75t_L g2586 ( 
.A(n_2358),
.Y(n_2586)
);

BUFx2_ASAP7_75t_L g2587 ( 
.A(n_2442),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2273),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2442),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2351),
.Y(n_2590)
);

BUFx12f_ASAP7_75t_L g2591 ( 
.A(n_2312),
.Y(n_2591)
);

OAI21x1_ASAP7_75t_L g2592 ( 
.A1(n_2394),
.A2(n_2206),
.B(n_2195),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2274),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2351),
.Y(n_2594)
);

AO21x1_ASAP7_75t_L g2595 ( 
.A1(n_2349),
.A2(n_2083),
.B(n_2090),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2385),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2262),
.B(n_2092),
.Y(n_2597)
);

CKINVDCx11_ASAP7_75t_R g2598 ( 
.A(n_2312),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2253),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2476),
.A2(n_1965),
.B1(n_1874),
.B2(n_1903),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_SL g2601 ( 
.A1(n_2535),
.A2(n_1918),
.B1(n_1923),
.B2(n_1939),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2274),
.Y(n_2602)
);

OAI22xp5_ASAP7_75t_L g2603 ( 
.A1(n_2282),
.A2(n_2180),
.B1(n_2240),
.B2(n_1926),
.Y(n_2603)
);

HB1xp67_ASAP7_75t_L g2604 ( 
.A(n_2385),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_L g2605 ( 
.A1(n_2476),
.A2(n_2457),
.B1(n_2412),
.B2(n_2558),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2266),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2462),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2280),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2267),
.Y(n_2609)
);

INVx3_ASAP7_75t_L g2610 ( 
.A(n_2441),
.Y(n_2610)
);

NOR2xp33_ASAP7_75t_L g2611 ( 
.A(n_2322),
.B(n_2210),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2462),
.Y(n_2612)
);

INVx1_ASAP7_75t_SL g2613 ( 
.A(n_2360),
.Y(n_2613)
);

OAI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2282),
.A2(n_2121),
.B1(n_1963),
.B2(n_1981),
.Y(n_2614)
);

INVx2_ASAP7_75t_SL g2615 ( 
.A(n_2254),
.Y(n_2615)
);

AOI22xp33_ASAP7_75t_SL g2616 ( 
.A1(n_2558),
.A2(n_2026),
.B1(n_2020),
.B2(n_2055),
.Y(n_2616)
);

AO21x1_ASAP7_75t_L g2617 ( 
.A1(n_2349),
.A2(n_2281),
.B(n_2451),
.Y(n_2617)
);

OAI21x1_ASAP7_75t_L g2618 ( 
.A1(n_2491),
.A2(n_2211),
.B(n_2217),
.Y(n_2618)
);

OR2x2_ASAP7_75t_L g2619 ( 
.A(n_2416),
.B(n_2268),
.Y(n_2619)
);

OAI22xp33_ASAP7_75t_L g2620 ( 
.A1(n_2558),
.A2(n_2096),
.B1(n_2008),
.B2(n_2009),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2269),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2291),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2282),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_L g2624 ( 
.A1(n_2412),
.A2(n_1879),
.B1(n_2040),
.B2(n_2233),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2301),
.Y(n_2625)
);

BUFx2_ASAP7_75t_SL g2626 ( 
.A(n_2358),
.Y(n_2626)
);

BUFx3_ASAP7_75t_L g2627 ( 
.A(n_2254),
.Y(n_2627)
);

CKINVDCx11_ASAP7_75t_R g2628 ( 
.A(n_2341),
.Y(n_2628)
);

AOI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2557),
.A2(n_2197),
.B1(n_2244),
.B2(n_2225),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2303),
.Y(n_2630)
);

CKINVDCx11_ASAP7_75t_R g2631 ( 
.A(n_2341),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2310),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2376),
.Y(n_2633)
);

BUFx6f_ASAP7_75t_L g2634 ( 
.A(n_2356),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_2378),
.Y(n_2635)
);

OAI22xp33_ASAP7_75t_L g2636 ( 
.A1(n_2445),
.A2(n_2427),
.B1(n_2361),
.B2(n_2348),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2326),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2260),
.B(n_2068),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_2286),
.Y(n_2639)
);

AOI22xp33_ASAP7_75t_SL g2640 ( 
.A1(n_2361),
.A2(n_2134),
.B1(n_1921),
.B2(n_2168),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2327),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2441),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2329),
.Y(n_2643)
);

AND2x2_ASAP7_75t_L g2644 ( 
.A(n_2445),
.B(n_1937),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2445),
.B(n_2112),
.Y(n_2645)
);

OA21x2_ASAP7_75t_L g2646 ( 
.A1(n_2583),
.A2(n_2490),
.B(n_2371),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2378),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2338),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2296),
.Y(n_2649)
);

BUFx6f_ASAP7_75t_L g2650 ( 
.A(n_2356),
.Y(n_2650)
);

INVx6_ASAP7_75t_L g2651 ( 
.A(n_2299),
.Y(n_2651)
);

NOR2x1_ASAP7_75t_SL g2652 ( 
.A(n_2537),
.B(n_1916),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2453),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2375),
.A2(n_2051),
.B1(n_2033),
.B2(n_2084),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2401),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2270),
.Y(n_2656)
);

AO21x1_ASAP7_75t_L g2657 ( 
.A1(n_2281),
.A2(n_2169),
.B(n_1895),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_2453),
.Y(n_2658)
);

INVx4_ASAP7_75t_L g2659 ( 
.A(n_2464),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2375),
.A2(n_2251),
.B1(n_2194),
.B2(n_2248),
.Y(n_2660)
);

BUFx12f_ASAP7_75t_L g2661 ( 
.A(n_2270),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2389),
.Y(n_2662)
);

INVx6_ASAP7_75t_L g2663 ( 
.A(n_2299),
.Y(n_2663)
);

INVxp67_ASAP7_75t_L g2664 ( 
.A(n_2567),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2408),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2557),
.A2(n_2201),
.B1(n_1888),
.B2(n_1997),
.Y(n_2666)
);

OAI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2348),
.A2(n_2050),
.B1(n_1917),
.B2(n_2078),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_SL g2668 ( 
.A1(n_2416),
.A2(n_2061),
.B1(n_2117),
.B2(n_2039),
.Y(n_2668)
);

AOI22xp33_ASAP7_75t_L g2669 ( 
.A1(n_2376),
.A2(n_2237),
.B1(n_2174),
.B2(n_2231),
.Y(n_2669)
);

INVx6_ASAP7_75t_L g2670 ( 
.A(n_2286),
.Y(n_2670)
);

HB1xp67_ASAP7_75t_L g2671 ( 
.A(n_2348),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2460),
.Y(n_2672)
);

CKINVDCx11_ASAP7_75t_R g2673 ( 
.A(n_2343),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2468),
.Y(n_2674)
);

BUFx2_ASAP7_75t_R g2675 ( 
.A(n_2309),
.Y(n_2675)
);

NOR2xp67_ASAP7_75t_R g2676 ( 
.A(n_2265),
.B(n_2023),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_SL g2677 ( 
.A1(n_2398),
.A2(n_2085),
.B1(n_2104),
.B2(n_2097),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2260),
.B(n_2069),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2437),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2362),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2369),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2437),
.Y(n_2682)
);

BUFx3_ASAP7_75t_L g2683 ( 
.A(n_2300),
.Y(n_2683)
);

INVx4_ASAP7_75t_L g2684 ( 
.A(n_2464),
.Y(n_2684)
);

BUFx2_ASAP7_75t_SL g2685 ( 
.A(n_2321),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2381),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2395),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2422),
.Y(n_2688)
);

AOI21x1_ASAP7_75t_L g2689 ( 
.A1(n_2261),
.A2(n_2006),
.B(n_1967),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2571),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2426),
.Y(n_2691)
);

CKINVDCx20_ASAP7_75t_R g2692 ( 
.A(n_2474),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2469),
.B(n_1969),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2440),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2379),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2446),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2402),
.B(n_2155),
.Y(n_2697)
);

OR2x2_ASAP7_75t_L g2698 ( 
.A(n_2416),
.B(n_2024),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2452),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2302),
.Y(n_2700)
);

BUFx10_ASAP7_75t_L g2701 ( 
.A(n_2536),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_SL g2702 ( 
.A1(n_2377),
.A2(n_2117),
.B1(n_2145),
.B2(n_2030),
.Y(n_2702)
);

INVx3_ASAP7_75t_L g2703 ( 
.A(n_2389),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2571),
.Y(n_2704)
);

BUFx3_ASAP7_75t_L g2705 ( 
.A(n_2300),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2366),
.A2(n_2227),
.B1(n_2203),
.B2(n_2181),
.Y(n_2706)
);

OAI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2414),
.A2(n_2067),
.B1(n_2032),
.B2(n_2053),
.Y(n_2707)
);

INVx3_ASAP7_75t_L g2708 ( 
.A(n_2533),
.Y(n_2708)
);

INVx1_ASAP7_75t_SL g2709 ( 
.A(n_2454),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2298),
.A2(n_2120),
.B1(n_1955),
.B2(n_1960),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_SL g2711 ( 
.A1(n_2377),
.A2(n_2146),
.B1(n_2141),
.B2(n_2042),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2277),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2366),
.A2(n_1943),
.B1(n_1954),
.B2(n_1941),
.Y(n_2713)
);

INVx2_ASAP7_75t_SL g2714 ( 
.A(n_2537),
.Y(n_2714)
);

BUFx10_ASAP7_75t_L g2715 ( 
.A(n_2536),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_2363),
.Y(n_2716)
);

HB1xp67_ASAP7_75t_L g2717 ( 
.A(n_2295),
.Y(n_2717)
);

INVx3_ASAP7_75t_L g2718 ( 
.A(n_2533),
.Y(n_2718)
);

AOI22xp33_ASAP7_75t_L g2719 ( 
.A1(n_2265),
.A2(n_1929),
.B1(n_2137),
.B2(n_2103),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2287),
.B(n_1932),
.Y(n_2720)
);

NAND2x1p5_ASAP7_75t_L g2721 ( 
.A(n_2331),
.B(n_2019),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2363),
.Y(n_2722)
);

NOR2x1_ASAP7_75t_R g2723 ( 
.A(n_2343),
.B(n_2116),
.Y(n_2723)
);

INVxp67_ASAP7_75t_SL g2724 ( 
.A(n_2298),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2277),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_SL g2726 ( 
.A1(n_2386),
.A2(n_2128),
.B1(n_1900),
.B2(n_2147),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2386),
.A2(n_1913),
.B1(n_2057),
.B2(n_2226),
.Y(n_2727)
);

BUFx8_ASAP7_75t_L g2728 ( 
.A(n_2256),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2388),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2278),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2388),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2581),
.A2(n_2027),
.B1(n_1863),
.B2(n_2014),
.Y(n_2732)
);

AOI21xp33_ASAP7_75t_L g2733 ( 
.A1(n_2582),
.A2(n_2126),
.B(n_2013),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2324),
.B(n_1995),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2337),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2570),
.B(n_1894),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2388),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2399),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2399),
.Y(n_2739)
);

BUFx4f_ASAP7_75t_SL g2740 ( 
.A(n_2417),
.Y(n_2740)
);

AND2x6_ASAP7_75t_L g2741 ( 
.A(n_2289),
.B(n_2157),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2275),
.B(n_2142),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2337),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2399),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2489),
.Y(n_2745)
);

INVx3_ASAP7_75t_L g2746 ( 
.A(n_2418),
.Y(n_2746)
);

NAND2x1p5_ASAP7_75t_L g2747 ( 
.A(n_2331),
.B(n_2332),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2489),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2570),
.B(n_1891),
.Y(n_2749)
);

OAI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2428),
.A2(n_1880),
.B1(n_2018),
.B2(n_1996),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2489),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2568),
.Y(n_2752)
);

BUFx3_ASAP7_75t_L g2753 ( 
.A(n_2372),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2340),
.Y(n_2754)
);

OAI22xp33_ASAP7_75t_L g2755 ( 
.A1(n_2278),
.A2(n_1962),
.B1(n_2119),
.B2(n_2001),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2568),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2568),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2521),
.Y(n_2758)
);

CKINVDCx20_ASAP7_75t_R g2759 ( 
.A(n_2398),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2340),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2418),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2372),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2521),
.Y(n_2763)
);

OR2x2_ASAP7_75t_L g2764 ( 
.A(n_2484),
.B(n_2163),
.Y(n_2764)
);

BUFx3_ASAP7_75t_L g2765 ( 
.A(n_2290),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2418),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2364),
.B(n_2456),
.Y(n_2767)
);

AO21x1_ASAP7_75t_L g2768 ( 
.A1(n_2451),
.A2(n_2179),
.B(n_2320),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2478),
.B(n_2179),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2439),
.Y(n_2770)
);

NAND2x1p5_ASAP7_75t_L g2771 ( 
.A(n_2332),
.B(n_2179),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2545),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2545),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_2487),
.Y(n_2774)
);

INVx6_ASAP7_75t_L g2775 ( 
.A(n_2368),
.Y(n_2775)
);

NAND2x1p5_ASAP7_75t_L g2776 ( 
.A(n_2334),
.B(n_2356),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2448),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2325),
.B(n_2354),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2439),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2289),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2289),
.Y(n_2781)
);

AOI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2509),
.A2(n_2313),
.B1(n_2542),
.B2(n_2481),
.Y(n_2782)
);

AOI22xp33_ASAP7_75t_SL g2783 ( 
.A1(n_2574),
.A2(n_2494),
.B1(n_2508),
.B2(n_2479),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2498),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2322),
.A2(n_2578),
.B1(n_2584),
.B2(n_2514),
.Y(n_2785)
);

INVx3_ASAP7_75t_L g2786 ( 
.A(n_2448),
.Y(n_2786)
);

INVx8_ASAP7_75t_L g2787 ( 
.A(n_2536),
.Y(n_2787)
);

BUFx2_ASAP7_75t_L g2788 ( 
.A(n_2407),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2498),
.Y(n_2789)
);

OR2x6_ASAP7_75t_L g2790 ( 
.A(n_2257),
.B(n_2259),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_2356),
.Y(n_2791)
);

OAI22xp33_ASAP7_75t_SL g2792 ( 
.A1(n_2257),
.A2(n_2259),
.B1(n_2297),
.B2(n_2271),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2501),
.Y(n_2793)
);

BUFx2_ASAP7_75t_R g2794 ( 
.A(n_2272),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_SL g2795 ( 
.A1(n_2494),
.A2(n_2508),
.B1(n_2479),
.B2(n_2536),
.Y(n_2795)
);

BUFx12f_ASAP7_75t_L g2796 ( 
.A(n_2417),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_L g2797 ( 
.A1(n_2578),
.A2(n_2584),
.B1(n_2542),
.B2(n_2465),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2501),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2512),
.Y(n_2799)
);

OA21x2_ASAP7_75t_L g2800 ( 
.A1(n_2490),
.A2(n_2320),
.B(n_2580),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2577),
.A2(n_2528),
.B1(n_2546),
.B2(n_2540),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2512),
.Y(n_2802)
);

AOI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_2261),
.A2(n_2471),
.B(n_2551),
.Y(n_2803)
);

NAND2x1p5_ASAP7_75t_L g2804 ( 
.A(n_2334),
.B(n_2380),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2492),
.B(n_2405),
.Y(n_2805)
);

OAI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2428),
.A2(n_2539),
.B1(n_2271),
.B2(n_2297),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2502),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2516),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2380),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2516),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2380),
.Y(n_2811)
);

INVx3_ASAP7_75t_L g2812 ( 
.A(n_2448),
.Y(n_2812)
);

BUFx4f_ASAP7_75t_L g2813 ( 
.A(n_2536),
.Y(n_2813)
);

BUFx4f_ASAP7_75t_SL g2814 ( 
.A(n_2368),
.Y(n_2814)
);

BUFx2_ASAP7_75t_L g2815 ( 
.A(n_2407),
.Y(n_2815)
);

INVx1_ASAP7_75t_SL g2816 ( 
.A(n_2345),
.Y(n_2816)
);

CKINVDCx20_ASAP7_75t_R g2817 ( 
.A(n_2450),
.Y(n_2817)
);

INVxp33_ASAP7_75t_L g2818 ( 
.A(n_2276),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2485),
.B(n_2504),
.Y(n_2819)
);

CKINVDCx11_ASAP7_75t_R g2820 ( 
.A(n_2450),
.Y(n_2820)
);

INVx6_ASAP7_75t_L g2821 ( 
.A(n_2370),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2458),
.Y(n_2822)
);

AOI22xp33_ASAP7_75t_L g2823 ( 
.A1(n_2467),
.A2(n_2538),
.B1(n_2518),
.B2(n_2527),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2306),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2279),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2458),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2458),
.Y(n_2827)
);

AO21x1_ASAP7_75t_L g2828 ( 
.A1(n_2314),
.A2(n_2323),
.B(n_2383),
.Y(n_2828)
);

CKINVDCx11_ASAP7_75t_R g2829 ( 
.A(n_2520),
.Y(n_2829)
);

HB1xp67_ASAP7_75t_L g2830 ( 
.A(n_2425),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2306),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2306),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2306),
.Y(n_2833)
);

OR2x6_ASAP7_75t_L g2834 ( 
.A(n_2383),
.B(n_2539),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2306),
.Y(n_2835)
);

BUFx3_ASAP7_75t_L g2836 ( 
.A(n_2290),
.Y(n_2836)
);

BUFx2_ASAP7_75t_L g2837 ( 
.A(n_2517),
.Y(n_2837)
);

BUFx12f_ASAP7_75t_L g2838 ( 
.A(n_2370),
.Y(n_2838)
);

INVx2_ASAP7_75t_SL g2839 ( 
.A(n_2307),
.Y(n_2839)
);

AOI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2423),
.A2(n_2530),
.B1(n_2531),
.B2(n_2506),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2306),
.Y(n_2841)
);

OAI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2539),
.A2(n_2576),
.B1(n_2505),
.B2(n_2524),
.Y(n_2842)
);

AO21x1_ASAP7_75t_SL g2843 ( 
.A1(n_2409),
.A2(n_2421),
.B(n_2423),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2486),
.Y(n_2844)
);

INVx2_ASAP7_75t_SL g2845 ( 
.A(n_2307),
.Y(n_2845)
);

AOI22xp33_ASAP7_75t_SL g2846 ( 
.A1(n_2494),
.A2(n_2433),
.B1(n_2382),
.B2(n_2315),
.Y(n_2846)
);

OA21x2_ASAP7_75t_L g2847 ( 
.A1(n_2374),
.A2(n_2436),
.B(n_2435),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2486),
.Y(n_2848)
);

HB1xp67_ASAP7_75t_L g2849 ( 
.A(n_2438),
.Y(n_2849)
);

INVx3_ASAP7_75t_L g2850 ( 
.A(n_2264),
.Y(n_2850)
);

BUFx3_ASAP7_75t_L g2851 ( 
.A(n_2345),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2486),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2380),
.Y(n_2853)
);

AOI22xp5_ASAP7_75t_SL g2854 ( 
.A1(n_2494),
.A2(n_2429),
.B1(n_2520),
.B2(n_2288),
.Y(n_2854)
);

OAI21x1_ASAP7_75t_L g2855 ( 
.A1(n_2579),
.A2(n_2350),
.B(n_2342),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2534),
.B(n_2541),
.Y(n_2856)
);

INVx6_ASAP7_75t_L g2857 ( 
.A(n_2315),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2410),
.B(n_2560),
.Y(n_2858)
);

BUFx2_ASAP7_75t_L g2859 ( 
.A(n_2517),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2497),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2323),
.Y(n_2861)
);

HB1xp67_ASAP7_75t_L g2862 ( 
.A(n_2283),
.Y(n_2862)
);

INVx1_ASAP7_75t_SL g2863 ( 
.A(n_2359),
.Y(n_2863)
);

INVx3_ASAP7_75t_L g2864 ( 
.A(n_2264),
.Y(n_2864)
);

BUFx12f_ASAP7_75t_L g2865 ( 
.A(n_2318),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_SL g2866 ( 
.A1(n_2494),
.A2(n_2505),
.B1(n_2513),
.B2(n_2524),
.Y(n_2866)
);

A2O1A1Ixp33_ASAP7_75t_L g2867 ( 
.A1(n_2854),
.A2(n_2496),
.B(n_2510),
.C(n_2421),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2662),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2598),
.Y(n_2869)
);

BUFx12f_ASAP7_75t_L g2870 ( 
.A(n_2628),
.Y(n_2870)
);

OR2x2_ASAP7_75t_SL g2871 ( 
.A(n_2651),
.B(n_2429),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2679),
.Y(n_2872)
);

CKINVDCx16_ASAP7_75t_R g2873 ( 
.A(n_2591),
.Y(n_2873)
);

NOR3xp33_ASAP7_75t_SL g2874 ( 
.A(n_2636),
.B(n_2825),
.C(n_2656),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2690),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_2631),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2599),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2590),
.B(n_2393),
.Y(n_2878)
);

O2A1O1Ixp33_ASAP7_75t_L g2879 ( 
.A1(n_2707),
.A2(n_2563),
.B(n_2519),
.C(n_2573),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2682),
.Y(n_2880)
);

NOR2x1_ASAP7_75t_L g2881 ( 
.A(n_2834),
.B(n_2384),
.Y(n_2881)
);

CKINVDCx16_ASAP7_75t_R g2882 ( 
.A(n_2796),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2606),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2673),
.Y(n_2884)
);

NOR2x1p5_ASAP7_75t_L g2885 ( 
.A(n_2659),
.B(n_2292),
.Y(n_2885)
);

NAND2xp33_ASAP7_75t_R g2886 ( 
.A(n_2587),
.B(n_2522),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2585),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2594),
.B(n_2353),
.Y(n_2888)
);

NAND3xp33_ASAP7_75t_L g2889 ( 
.A(n_2600),
.B(n_2500),
.C(n_2293),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2588),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2819),
.B(n_2563),
.Y(n_2891)
);

OR2x2_ASAP7_75t_L g2892 ( 
.A(n_2607),
.B(n_2459),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2616),
.A2(n_2576),
.B1(n_2575),
.B2(n_2500),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_2820),
.Y(n_2894)
);

OR2x2_ASAP7_75t_L g2895 ( 
.A(n_2612),
.B(n_2384),
.Y(n_2895)
);

OR2x6_ASAP7_75t_L g2896 ( 
.A(n_2626),
.B(n_2294),
.Y(n_2896)
);

O2A1O1Ixp33_ASAP7_75t_SL g2897 ( 
.A1(n_2842),
.A2(n_2314),
.B(n_2556),
.C(n_2473),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2834),
.A2(n_2513),
.B1(n_2311),
.B2(n_2575),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2697),
.B(n_2560),
.Y(n_2899)
);

INVxp33_ASAP7_75t_SL g2900 ( 
.A(n_2829),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2767),
.B(n_2258),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2593),
.Y(n_2902)
);

INVxp67_ASAP7_75t_L g2903 ( 
.A(n_2830),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2602),
.Y(n_2904)
);

NAND2xp33_ASAP7_75t_R g2905 ( 
.A(n_2589),
.B(n_2288),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_R g2906 ( 
.A(n_2740),
.B(n_2352),
.Y(n_2906)
);

HB1xp67_ASAP7_75t_L g2907 ( 
.A(n_2704),
.Y(n_2907)
);

HB1xp67_ASAP7_75t_L g2908 ( 
.A(n_2596),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_R g2909 ( 
.A(n_2814),
.B(n_2817),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2819),
.B(n_2552),
.Y(n_2910)
);

INVx2_ASAP7_75t_SL g2911 ( 
.A(n_2670),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2792),
.B(n_2264),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2616),
.A2(n_2317),
.B1(n_2556),
.B2(n_2473),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_2792),
.B(n_2264),
.Y(n_2914)
);

INVx2_ASAP7_75t_SL g2915 ( 
.A(n_2670),
.Y(n_2915)
);

CKINVDCx16_ASAP7_75t_R g2916 ( 
.A(n_2838),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2608),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2661),
.Y(n_2918)
);

OR2x6_ASAP7_75t_L g2919 ( 
.A(n_2787),
.B(n_2496),
.Y(n_2919)
);

CKINVDCx5p33_ASAP7_75t_R g2920 ( 
.A(n_2635),
.Y(n_2920)
);

AND2x2_ASAP7_75t_SL g2921 ( 
.A(n_2813),
.B(n_2288),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2647),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2834),
.Y(n_2923)
);

CKINVDCx16_ASAP7_75t_R g2924 ( 
.A(n_2759),
.Y(n_2924)
);

NOR2xp33_ASAP7_75t_R g2925 ( 
.A(n_2714),
.B(n_2258),
.Y(n_2925)
);

CKINVDCx5p33_ASAP7_75t_R g2926 ( 
.A(n_2651),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2805),
.B(n_2325),
.Y(n_2927)
);

OR2x6_ASAP7_75t_L g2928 ( 
.A(n_2787),
.B(n_2510),
.Y(n_2928)
);

AOI22xp33_ASAP7_75t_L g2929 ( 
.A1(n_2601),
.A2(n_2397),
.B1(n_2562),
.B2(n_2409),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2663),
.Y(n_2930)
);

BUFx3_ASAP7_75t_L g2931 ( 
.A(n_2639),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_R g2932 ( 
.A(n_2662),
.B(n_2503),
.Y(n_2932)
);

OR2x6_ASAP7_75t_L g2933 ( 
.A(n_2787),
.B(n_2283),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2856),
.B(n_2552),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2604),
.B(n_2354),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2609),
.Y(n_2936)
);

INVx6_ASAP7_75t_L g2937 ( 
.A(n_2775),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2858),
.B(n_2532),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2663),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2621),
.Y(n_2940)
);

AO31x2_ASAP7_75t_L g2941 ( 
.A1(n_2768),
.A2(n_2293),
.A3(n_2543),
.B(n_2411),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2622),
.Y(n_2942)
);

CKINVDCx16_ASAP7_75t_R g2943 ( 
.A(n_2692),
.Y(n_2943)
);

INVx2_ASAP7_75t_SL g2944 ( 
.A(n_2775),
.Y(n_2944)
);

OR2x6_ASAP7_75t_L g2945 ( 
.A(n_2821),
.B(n_2790),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2862),
.B(n_2553),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2625),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2630),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_R g2949 ( 
.A(n_2703),
.B(n_2503),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_2695),
.Y(n_2950)
);

HB1xp67_ASAP7_75t_L g2951 ( 
.A(n_2807),
.Y(n_2951)
);

AOI22xp33_ASAP7_75t_L g2952 ( 
.A1(n_2595),
.A2(n_2605),
.B1(n_2603),
.B2(n_2640),
.Y(n_2952)
);

INVx3_ASAP7_75t_L g2953 ( 
.A(n_2703),
.Y(n_2953)
);

OAI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2614),
.A2(n_2515),
.B(n_2397),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2856),
.B(n_2319),
.Y(n_2955)
);

OR2x2_ASAP7_75t_SL g2956 ( 
.A(n_2633),
.B(n_2316),
.Y(n_2956)
);

CKINVDCx20_ASAP7_75t_R g2957 ( 
.A(n_2728),
.Y(n_2957)
);

OR2x2_ASAP7_75t_L g2958 ( 
.A(n_2613),
.B(n_2285),
.Y(n_2958)
);

AOI211xp5_ASAP7_75t_SL g2959 ( 
.A1(n_2806),
.A2(n_2308),
.B(n_2357),
.C(n_2367),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2632),
.Y(n_2960)
);

INVx3_ASAP7_75t_L g2961 ( 
.A(n_2708),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2603),
.A2(n_2614),
.B1(n_2620),
.B2(n_2645),
.Y(n_2962)
);

NAND2xp33_ASAP7_75t_R g2963 ( 
.A(n_2708),
.B(n_2316),
.Y(n_2963)
);

OAI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2702),
.A2(n_2515),
.B(n_2308),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2634),
.Y(n_2965)
);

BUFx3_ASAP7_75t_L g2966 ( 
.A(n_2627),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_SL g2967 ( 
.A1(n_2854),
.A2(n_2316),
.B1(n_2263),
.B2(n_2305),
.Y(n_2967)
);

NAND2xp33_ASAP7_75t_R g2968 ( 
.A(n_2718),
.B(n_2255),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2637),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2641),
.Y(n_2970)
);

AOI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2667),
.A2(n_2403),
.B1(n_2565),
.B2(n_2432),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2839),
.B(n_2561),
.Y(n_2972)
);

INVxp67_ASAP7_75t_L g2973 ( 
.A(n_2849),
.Y(n_2973)
);

NOR2x1_ASAP7_75t_SL g2974 ( 
.A(n_2790),
.B(n_2559),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2845),
.B(n_2572),
.Y(n_2975)
);

BUFx10_ASAP7_75t_L g2976 ( 
.A(n_2821),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2683),
.B(n_2572),
.Y(n_2977)
);

NAND2xp33_ASAP7_75t_R g2978 ( 
.A(n_2718),
.B(n_2255),
.Y(n_2978)
);

BUFx2_ASAP7_75t_L g2979 ( 
.A(n_2851),
.Y(n_2979)
);

NAND2xp33_ASAP7_75t_R g2980 ( 
.A(n_2837),
.B(n_2859),
.Y(n_2980)
);

BUFx4f_ASAP7_75t_SL g2981 ( 
.A(n_2728),
.Y(n_2981)
);

OR2x2_ASAP7_75t_L g2982 ( 
.A(n_2613),
.B(n_2335),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2643),
.Y(n_2983)
);

OR2x2_ASAP7_75t_L g2984 ( 
.A(n_2709),
.B(n_2335),
.Y(n_2984)
);

NAND2x1p5_ASAP7_75t_L g2985 ( 
.A(n_2659),
.B(n_2413),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2782),
.B(n_2511),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2675),
.Y(n_2987)
);

AO31x2_ASAP7_75t_L g2988 ( 
.A1(n_2617),
.A2(n_2424),
.A3(n_2342),
.B(n_2350),
.Y(n_2988)
);

AOI22xp33_ASAP7_75t_SL g2989 ( 
.A1(n_2623),
.A2(n_2304),
.B1(n_2305),
.B2(n_2403),
.Y(n_2989)
);

NAND2xp33_ASAP7_75t_SL g2990 ( 
.A(n_2671),
.B(n_2304),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2648),
.Y(n_2991)
);

INVxp67_ASAP7_75t_L g2992 ( 
.A(n_2774),
.Y(n_2992)
);

NAND2xp33_ASAP7_75t_R g2993 ( 
.A(n_2788),
.B(n_2815),
.Y(n_2993)
);

OAI22xp5_ASAP7_75t_L g2994 ( 
.A1(n_2866),
.A2(n_2311),
.B1(n_2419),
.B2(n_2390),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2705),
.B(n_2336),
.Y(n_2995)
);

HB1xp67_ASAP7_75t_L g2996 ( 
.A(n_2863),
.Y(n_2996)
);

NOR2x1p5_ASAP7_75t_L g2997 ( 
.A(n_2684),
.B(n_2480),
.Y(n_2997)
);

AND2x4_ASAP7_75t_L g2998 ( 
.A(n_2790),
.B(n_2778),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2675),
.Y(n_2999)
);

INVxp67_ASAP7_75t_L g3000 ( 
.A(n_2717),
.Y(n_3000)
);

OR2x6_ASAP7_75t_L g3001 ( 
.A(n_2684),
.B(n_2685),
.Y(n_3001)
);

AND2x4_ASAP7_75t_SL g3002 ( 
.A(n_2701),
.B(n_2357),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2709),
.B(n_2863),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_2794),
.Y(n_3004)
);

HB1xp67_ASAP7_75t_L g3005 ( 
.A(n_2730),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2655),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2665),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2778),
.B(n_2367),
.Y(n_3008)
);

HB1xp67_ASAP7_75t_L g3009 ( 
.A(n_2649),
.Y(n_3009)
);

AND2x4_ASAP7_75t_L g3010 ( 
.A(n_2610),
.B(n_2373),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2782),
.B(n_2511),
.Y(n_3011)
);

CKINVDCx16_ASAP7_75t_R g3012 ( 
.A(n_2865),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2794),
.Y(n_3013)
);

AOI22xp33_ASAP7_75t_L g3014 ( 
.A1(n_2667),
.A2(n_2734),
.B1(n_2644),
.B2(n_2702),
.Y(n_3014)
);

AND2x4_ASAP7_75t_L g3015 ( 
.A(n_2610),
.B(n_2373),
.Y(n_3015)
);

INVxp67_ASAP7_75t_SL g3016 ( 
.A(n_2724),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2716),
.B(n_2336),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_R g3018 ( 
.A(n_2642),
.B(n_2347),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2672),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2664),
.Y(n_3020)
);

BUFx6f_ASAP7_75t_L g3021 ( 
.A(n_2634),
.Y(n_3021)
);

CKINVDCx5p33_ASAP7_75t_R g3022 ( 
.A(n_2586),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2611),
.A2(n_2565),
.B1(n_2432),
.B2(n_2434),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_2624),
.A2(n_2344),
.B1(n_2346),
.B2(n_2400),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2722),
.B(n_2347),
.Y(n_3025)
);

INVx4_ASAP7_75t_L g3026 ( 
.A(n_2650),
.Y(n_3026)
);

BUFx3_ASAP7_75t_L g3027 ( 
.A(n_2753),
.Y(n_3027)
);

OR2x6_ASAP7_75t_L g3028 ( 
.A(n_2586),
.B(n_2525),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2674),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2680),
.B(n_2555),
.Y(n_3030)
);

AND2x4_ASAP7_75t_SL g3031 ( 
.A(n_2701),
.B(n_2355),
.Y(n_3031)
);

AO32x2_ASAP7_75t_L g3032 ( 
.A1(n_2727),
.A2(n_2549),
.A3(n_2564),
.B1(n_2328),
.B2(n_2415),
.Y(n_3032)
);

NAND2xp33_ASAP7_75t_R g3033 ( 
.A(n_2642),
.B(n_2255),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2762),
.B(n_2355),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2681),
.B(n_2555),
.Y(n_3035)
);

NAND2xp33_ASAP7_75t_SL g3036 ( 
.A(n_2653),
.B(n_2529),
.Y(n_3036)
);

OR2x2_ASAP7_75t_L g3037 ( 
.A(n_2816),
.B(n_2495),
.Y(n_3037)
);

CKINVDCx16_ASAP7_75t_R g3038 ( 
.A(n_2765),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_2816),
.B(n_2431),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2686),
.Y(n_3040)
);

NAND3xp33_ASAP7_75t_SL g3041 ( 
.A(n_2818),
.B(n_2493),
.C(n_2390),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2687),
.Y(n_3042)
);

BUFx2_ASAP7_75t_L g3043 ( 
.A(n_2653),
.Y(n_3043)
);

BUFx6f_ASAP7_75t_L g3044 ( 
.A(n_2650),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_2742),
.B(n_2415),
.Y(n_3045)
);

NAND2xp33_ASAP7_75t_R g3046 ( 
.A(n_2658),
.B(n_2482),
.Y(n_3046)
);

CKINVDCx5p33_ASAP7_75t_R g3047 ( 
.A(n_2615),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2836),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_R g3049 ( 
.A(n_2658),
.B(n_2264),
.Y(n_3049)
);

NOR3xp33_ASAP7_75t_SL g3050 ( 
.A(n_2861),
.B(n_2279),
.C(n_2419),
.Y(n_3050)
);

AO31x2_ASAP7_75t_L g3051 ( 
.A1(n_2803),
.A2(n_2392),
.A3(n_2387),
.B(n_2526),
.Y(n_3051)
);

AND2x2_ASAP7_75t_SL g3052 ( 
.A(n_2791),
.B(n_2809),
.Y(n_3052)
);

NAND3xp33_ASAP7_75t_L g3053 ( 
.A(n_2801),
.B(n_2284),
.C(n_2488),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2720),
.B(n_2544),
.Y(n_3054)
);

AOI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2654),
.A2(n_2330),
.B1(n_2477),
.B2(n_2523),
.Y(n_3055)
);

OAI21xp5_ASAP7_75t_SL g3056 ( 
.A1(n_2795),
.A2(n_2404),
.B(n_2447),
.Y(n_3056)
);

NOR3xp33_ASAP7_75t_SL g3057 ( 
.A(n_2727),
.B(n_2466),
.C(n_2544),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2688),
.B(n_2547),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2691),
.Y(n_3059)
);

AO31x2_ASAP7_75t_L g3060 ( 
.A1(n_2803),
.A2(n_2391),
.A3(n_2392),
.B(n_2396),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_2857),
.Y(n_3061)
);

NOR2xp33_ASAP7_75t_R g3062 ( 
.A(n_2715),
.B(n_2264),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2694),
.B(n_2547),
.Y(n_3063)
);

NAND2xp33_ASAP7_75t_SL g3064 ( 
.A(n_2791),
.B(n_2339),
.Y(n_3064)
);

OAI22xp5_ASAP7_75t_L g3065 ( 
.A1(n_2629),
.A2(n_2430),
.B1(n_2507),
.B2(n_2413),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_R g3066 ( 
.A(n_2715),
.B(n_2857),
.Y(n_3066)
);

NAND2xp33_ASAP7_75t_SL g3067 ( 
.A(n_2791),
.B(n_2339),
.Y(n_3067)
);

NAND2xp33_ASAP7_75t_R g3068 ( 
.A(n_2850),
.B(n_2482),
.Y(n_3068)
);

AND2x4_ASAP7_75t_L g3069 ( 
.A(n_2729),
.B(n_2413),
.Y(n_3069)
);

HB1xp67_ASAP7_75t_L g3070 ( 
.A(n_2784),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2696),
.B(n_2523),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2699),
.B(n_2431),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2700),
.Y(n_3073)
);

CKINVDCx16_ASAP7_75t_R g3074 ( 
.A(n_2619),
.Y(n_3074)
);

AO32x1_ASAP7_75t_L g3075 ( 
.A1(n_2860),
.A2(n_2564),
.A3(n_2406),
.B1(n_2420),
.B2(n_2550),
.Y(n_3075)
);

OAI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_2629),
.A2(n_2507),
.B1(n_2413),
.B2(n_2430),
.Y(n_3076)
);

CKINVDCx16_ASAP7_75t_R g3077 ( 
.A(n_2809),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2789),
.Y(n_3078)
);

OAI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2666),
.A2(n_2507),
.B1(n_2430),
.B2(n_2475),
.Y(n_3079)
);

AND2x4_ASAP7_75t_L g3080 ( 
.A(n_2731),
.B(n_2430),
.Y(n_3080)
);

BUFx3_ASAP7_75t_L g3081 ( 
.A(n_2776),
.Y(n_3081)
);

INVx3_ASAP7_75t_L g3082 ( 
.A(n_2747),
.Y(n_3082)
);

AOI222xp33_ASAP7_75t_L g3083 ( 
.A1(n_2723),
.A2(n_2548),
.B1(n_2569),
.B2(n_2554),
.C1(n_2374),
.C2(n_2435),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2597),
.B(n_2785),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2798),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2747),
.B(n_2444),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2799),
.Y(n_3087)
);

OR2x6_ASAP7_75t_L g3088 ( 
.A(n_2776),
.B(n_2548),
.Y(n_3088)
);

NAND2x1p5_ASAP7_75t_L g3089 ( 
.A(n_2811),
.B(n_2507),
.Y(n_3089)
);

INVx3_ASAP7_75t_L g3090 ( 
.A(n_2804),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2668),
.A2(n_2365),
.B1(n_2333),
.B2(n_2443),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2797),
.B(n_2444),
.Y(n_3092)
);

OR2x2_ASAP7_75t_L g3093 ( 
.A(n_2802),
.B(n_2447),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2808),
.Y(n_3094)
);

NAND2xp33_ASAP7_75t_R g3095 ( 
.A(n_2850),
.B(n_2482),
.Y(n_3095)
);

NAND2xp33_ASAP7_75t_R g3096 ( 
.A(n_2864),
.B(n_2483),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2804),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2746),
.B(n_2455),
.Y(n_3098)
);

AND2x4_ASAP7_75t_L g3099 ( 
.A(n_3016),
.B(n_2864),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2938),
.B(n_2810),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2877),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2927),
.B(n_2737),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2887),
.Y(n_3103)
);

AND2x4_ASAP7_75t_SL g3104 ( 
.A(n_2933),
.B(n_2811),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2901),
.B(n_2738),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_3009),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_3058),
.B(n_2840),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2962),
.A2(n_2657),
.B1(n_2843),
.B2(n_2666),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2872),
.Y(n_3109)
);

INVx3_ASAP7_75t_L g3110 ( 
.A(n_2998),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3045),
.B(n_2769),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2880),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2883),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2936),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_3054),
.B(n_2769),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_2899),
.B(n_2739),
.Y(n_3116)
);

INVx5_ASAP7_75t_L g3117 ( 
.A(n_3001),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2890),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_3084),
.B(n_2744),
.Y(n_3119)
);

OR2x2_ASAP7_75t_L g3120 ( 
.A(n_2875),
.B(n_2735),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2998),
.B(n_2780),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2986),
.B(n_2712),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2907),
.B(n_2745),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2897),
.A2(n_2828),
.B(n_2847),
.Y(n_3124)
);

INVxp67_ASAP7_75t_L g3125 ( 
.A(n_2908),
.Y(n_3125)
);

HB1xp67_ASAP7_75t_L g3126 ( 
.A(n_3070),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3011),
.B(n_2725),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2902),
.Y(n_3128)
);

AND2x2_ASAP7_75t_L g3129 ( 
.A(n_2946),
.B(n_2748),
.Y(n_3129)
);

BUFx3_ASAP7_75t_L g3130 ( 
.A(n_3097),
.Y(n_3130)
);

BUFx2_ASAP7_75t_L g3131 ( 
.A(n_3018),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2940),
.Y(n_3132)
);

BUFx3_ASAP7_75t_L g3133 ( 
.A(n_3081),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_2935),
.B(n_2751),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2942),
.Y(n_3135)
);

HB1xp67_ASAP7_75t_L g3136 ( 
.A(n_3005),
.Y(n_3136)
);

OR2x2_ASAP7_75t_L g3137 ( 
.A(n_3003),
.B(n_2743),
.Y(n_3137)
);

AND2x2_ASAP7_75t_L g3138 ( 
.A(n_2996),
.B(n_2752),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_3063),
.B(n_2758),
.Y(n_3139)
);

INVxp67_ASAP7_75t_SL g3140 ( 
.A(n_2912),
.Y(n_3140)
);

OR2x2_ASAP7_75t_L g3141 ( 
.A(n_2951),
.B(n_2754),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_3074),
.B(n_2756),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2947),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2948),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2904),
.Y(n_3145)
);

OR2x2_ASAP7_75t_L g3146 ( 
.A(n_2955),
.B(n_2760),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2960),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_3014),
.A2(n_2783),
.B1(n_2823),
.B2(n_2846),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2969),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2952),
.B(n_2763),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2970),
.Y(n_3151)
);

NAND3xp33_ASAP7_75t_SL g3152 ( 
.A(n_2925),
.B(n_2721),
.C(n_2669),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2972),
.B(n_2757),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2917),
.Y(n_3154)
);

BUFx3_ASAP7_75t_L g3155 ( 
.A(n_2966),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_3072),
.B(n_2770),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_3078),
.B(n_2772),
.Y(n_3157)
);

OR2x2_ASAP7_75t_L g3158 ( 
.A(n_2892),
.B(n_2779),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_3043),
.B(n_2992),
.Y(n_3159)
);

BUFx3_ASAP7_75t_L g3160 ( 
.A(n_3027),
.Y(n_3160)
);

OA21x2_ASAP7_75t_L g3161 ( 
.A1(n_2867),
.A2(n_2592),
.B(n_2618),
.Y(n_3161)
);

BUFx3_ASAP7_75t_L g3162 ( 
.A(n_3048),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_2895),
.B(n_2793),
.Y(n_3163)
);

OR2x2_ASAP7_75t_L g3164 ( 
.A(n_2958),
.B(n_2781),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2983),
.Y(n_3165)
);

BUFx6f_ASAP7_75t_L g3166 ( 
.A(n_2965),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2977),
.B(n_2822),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_3085),
.B(n_2773),
.Y(n_3168)
);

BUFx10_ASAP7_75t_L g3169 ( 
.A(n_2896),
.Y(n_3169)
);

INVx5_ASAP7_75t_SL g3170 ( 
.A(n_2896),
.Y(n_3170)
);

AOI221xp5_ASAP7_75t_L g3171 ( 
.A1(n_2879),
.A2(n_2660),
.B1(n_2706),
.B2(n_2733),
.C(n_2711),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2991),
.Y(n_3172)
);

AOI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_2889),
.A2(n_2750),
.B1(n_2726),
.B2(n_2733),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3006),
.B(n_2826),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3007),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_3019),
.B(n_2827),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3029),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3040),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3042),
.Y(n_3179)
);

AND2x4_ASAP7_75t_SL g3180 ( 
.A(n_2933),
.B(n_2811),
.Y(n_3180)
);

OR2x2_ASAP7_75t_L g3181 ( 
.A(n_3038),
.B(n_2844),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_3059),
.B(n_2975),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3073),
.Y(n_3183)
);

NAND4xp25_ASAP7_75t_L g3184 ( 
.A(n_2893),
.B(n_2677),
.C(n_2732),
.D(n_2713),
.Y(n_3184)
);

INVx3_ASAP7_75t_L g3185 ( 
.A(n_3026),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2976),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_3000),
.B(n_2848),
.Y(n_3187)
);

BUFx2_ASAP7_75t_L g3188 ( 
.A(n_3049),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3087),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3077),
.B(n_2852),
.Y(n_3190)
);

AND2x4_ASAP7_75t_L g3191 ( 
.A(n_2881),
.B(n_2853),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3094),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2903),
.B(n_2771),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2878),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_2973),
.B(n_3092),
.Y(n_3195)
);

AND2x4_ASAP7_75t_L g3196 ( 
.A(n_2923),
.B(n_2853),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_2995),
.B(n_2771),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3017),
.B(n_2764),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_3025),
.B(n_2824),
.Y(n_3199)
);

HB1xp67_ASAP7_75t_L g3200 ( 
.A(n_3051),
.Y(n_3200)
);

INVx5_ASAP7_75t_L g3201 ( 
.A(n_3001),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_3034),
.B(n_2831),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2979),
.B(n_2832),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_3020),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2891),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_2982),
.B(n_2833),
.Y(n_3206)
);

INVx2_ASAP7_75t_SL g3207 ( 
.A(n_2976),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_3093),
.Y(n_3208)
);

AOI322xp5_ASAP7_75t_L g3209 ( 
.A1(n_2874),
.A2(n_2736),
.A3(n_2719),
.B1(n_2755),
.B2(n_2726),
.C1(n_2693),
.C2(n_2749),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2888),
.Y(n_3210)
);

INVxp67_ASAP7_75t_L g3211 ( 
.A(n_2914),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_3071),
.B(n_2638),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2984),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2971),
.B(n_2638),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_3037),
.B(n_3008),
.Y(n_3215)
);

AO21x2_ASAP7_75t_L g3216 ( 
.A1(n_3057),
.A2(n_2689),
.B(n_2855),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3008),
.B(n_2835),
.Y(n_3217)
);

NOR2x1_ASAP7_75t_R g3218 ( 
.A(n_2870),
.B(n_2853),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_3060),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2910),
.B(n_2678),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3039),
.B(n_2841),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2931),
.B(n_2746),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_2909),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3030),
.Y(n_3224)
);

OR2x2_ASAP7_75t_L g3225 ( 
.A(n_2934),
.B(n_2736),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3035),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_3010),
.B(n_3015),
.Y(n_3227)
);

INVx2_ASAP7_75t_SL g3228 ( 
.A(n_2937),
.Y(n_3228)
);

INVx3_ASAP7_75t_L g3229 ( 
.A(n_3026),
.Y(n_3229)
);

AND2x2_ASAP7_75t_L g3230 ( 
.A(n_3010),
.B(n_2761),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2954),
.B(n_2678),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3015),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3088),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3088),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_2937),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2945),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2913),
.B(n_2749),
.Y(n_3237)
);

AND2x2_ASAP7_75t_L g3238 ( 
.A(n_3195),
.B(n_2988),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3115),
.B(n_2988),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3126),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3103),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3115),
.B(n_2988),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3126),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3111),
.B(n_2941),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3136),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_3136),
.Y(n_3246)
);

OA211x2_ASAP7_75t_L g3247 ( 
.A1(n_3152),
.A2(n_3041),
.B(n_2964),
.C(n_3091),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3101),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_SL g3249 ( 
.A1(n_3131),
.A2(n_2898),
.B1(n_2994),
.B2(n_2974),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_3125),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3113),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3205),
.B(n_2929),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_3125),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_3103),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3114),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3111),
.B(n_2941),
.Y(n_3256)
);

INVx1_ASAP7_75t_SL g3257 ( 
.A(n_3155),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3132),
.Y(n_3258)
);

NAND3xp33_ASAP7_75t_L g3259 ( 
.A(n_3173),
.B(n_2959),
.C(n_3023),
.Y(n_3259)
);

NAND3xp33_ASAP7_75t_L g3260 ( 
.A(n_3173),
.B(n_2989),
.C(n_2905),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3135),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3194),
.B(n_2967),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3143),
.Y(n_3263)
);

AND2x4_ASAP7_75t_L g3264 ( 
.A(n_3233),
.B(n_2919),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_3234),
.B(n_2919),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3144),
.Y(n_3266)
);

INVxp67_ASAP7_75t_L g3267 ( 
.A(n_3155),
.Y(n_3267)
);

HB1xp67_ASAP7_75t_L g3268 ( 
.A(n_3106),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3215),
.B(n_3052),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3147),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3224),
.B(n_2710),
.Y(n_3271)
);

HB1xp67_ASAP7_75t_L g3272 ( 
.A(n_3120),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_3145),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3184),
.A2(n_3036),
.B1(n_3053),
.B2(n_2921),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3226),
.B(n_3210),
.Y(n_3275)
);

BUFx6f_ASAP7_75t_L g3276 ( 
.A(n_3166),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3119),
.B(n_3213),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3198),
.B(n_3159),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3149),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3151),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_3141),
.B(n_3012),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_3182),
.B(n_3098),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3220),
.B(n_2710),
.Y(n_3283)
);

AOI21xp33_ASAP7_75t_L g3284 ( 
.A1(n_3148),
.A2(n_3108),
.B(n_3150),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3122),
.B(n_2941),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_3211),
.B(n_2928),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3145),
.Y(n_3287)
);

CKINVDCx20_ASAP7_75t_R g3288 ( 
.A(n_3160),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3165),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3109),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3220),
.B(n_2741),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3122),
.B(n_3127),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3237),
.B(n_3100),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3172),
.Y(n_3294)
);

INVx2_ASAP7_75t_SL g3295 ( 
.A(n_3130),
.Y(n_3295)
);

NAND3xp33_ASAP7_75t_L g3296 ( 
.A(n_3209),
.B(n_3108),
.C(n_3171),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_3127),
.B(n_3032),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3237),
.B(n_2741),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3212),
.B(n_3032),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3212),
.B(n_3032),
.Y(n_3300)
);

INVxp67_ASAP7_75t_L g3301 ( 
.A(n_3160),
.Y(n_3301)
);

AND2x4_ASAP7_75t_L g3302 ( 
.A(n_3211),
.B(n_3110),
.Y(n_3302)
);

BUFx2_ASAP7_75t_L g3303 ( 
.A(n_3188),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3204),
.B(n_2741),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3175),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3112),
.Y(n_3306)
);

OR2x2_ASAP7_75t_L g3307 ( 
.A(n_3208),
.B(n_3047),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3225),
.B(n_2741),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3118),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3107),
.B(n_2646),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3107),
.B(n_2646),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3139),
.B(n_3206),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_3130),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_3139),
.B(n_2928),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3128),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3231),
.B(n_2800),
.Y(n_3316)
);

INVxp67_ASAP7_75t_L g3317 ( 
.A(n_3246),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3240),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3292),
.B(n_3177),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3241),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3278),
.B(n_3197),
.Y(n_3321)
);

OR2x2_ASAP7_75t_L g3322 ( 
.A(n_3272),
.B(n_3137),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3243),
.Y(n_3323)
);

OR2x2_ASAP7_75t_L g3324 ( 
.A(n_3312),
.B(n_3158),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_3249),
.A2(n_2871),
.B1(n_3148),
.B2(n_3117),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3248),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3241),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3312),
.B(n_3193),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3292),
.B(n_3178),
.Y(n_3329)
);

INVx3_ASAP7_75t_L g3330 ( 
.A(n_3295),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3251),
.Y(n_3331)
);

OR2x2_ASAP7_75t_L g3332 ( 
.A(n_3293),
.B(n_3146),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3277),
.B(n_3227),
.Y(n_3333)
);

AND2x4_ASAP7_75t_L g3334 ( 
.A(n_3286),
.B(n_3099),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3255),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3254),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3258),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3261),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_3295),
.B(n_3303),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3263),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3239),
.B(n_3179),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3266),
.Y(n_3342)
);

CKINVDCx16_ASAP7_75t_R g3343 ( 
.A(n_3288),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3277),
.B(n_3282),
.Y(n_3344)
);

OR2x2_ASAP7_75t_L g3345 ( 
.A(n_3268),
.B(n_3163),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3270),
.Y(n_3346)
);

NAND2x1p5_ASAP7_75t_L g3347 ( 
.A(n_3257),
.B(n_3117),
.Y(n_3347)
);

OR2x2_ASAP7_75t_L g3348 ( 
.A(n_3245),
.B(n_3164),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3314),
.B(n_3110),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3314),
.B(n_3221),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3254),
.Y(n_3351)
);

NOR3xp33_ASAP7_75t_L g3352 ( 
.A(n_3296),
.B(n_3152),
.C(n_3171),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3273),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_3250),
.B(n_3231),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3253),
.B(n_3142),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3279),
.Y(n_3356)
);

OR2x2_ASAP7_75t_L g3357 ( 
.A(n_3275),
.B(n_3183),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3313),
.B(n_3129),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_3288),
.B(n_3117),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3269),
.B(n_3199),
.Y(n_3360)
);

O2A1O1Ixp33_ASAP7_75t_L g3361 ( 
.A1(n_3284),
.A2(n_3184),
.B(n_3207),
.C(n_3186),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3280),
.Y(n_3362)
);

INVx1_ASAP7_75t_SL g3363 ( 
.A(n_3281),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3239),
.B(n_3189),
.Y(n_3364)
);

OR2x2_ASAP7_75t_L g3365 ( 
.A(n_3290),
.B(n_3192),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3242),
.B(n_3214),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3289),
.Y(n_3367)
);

INVx2_ASAP7_75t_L g3368 ( 
.A(n_3273),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3238),
.B(n_3202),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3238),
.B(n_3116),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3294),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3287),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3305),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3290),
.Y(n_3374)
);

OR2x2_ASAP7_75t_L g3375 ( 
.A(n_3306),
.B(n_3154),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3302),
.B(n_3264),
.Y(n_3376)
);

OR2x2_ASAP7_75t_L g3377 ( 
.A(n_3306),
.B(n_3309),
.Y(n_3377)
);

NAND2x1_ASAP7_75t_SL g3378 ( 
.A(n_3330),
.B(n_3185),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3366),
.B(n_3242),
.Y(n_3379)
);

OR2x2_ASAP7_75t_L g3380 ( 
.A(n_3366),
.B(n_3310),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3354),
.Y(n_3381)
);

O2A1O1Ixp5_ASAP7_75t_R g3382 ( 
.A1(n_3352),
.A2(n_3262),
.B(n_3252),
.C(n_3283),
.Y(n_3382)
);

AOI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3325),
.A2(n_3274),
.B1(n_3259),
.B2(n_3247),
.Y(n_3383)
);

NAND4xp25_ASAP7_75t_L g3384 ( 
.A(n_3352),
.B(n_3325),
.C(n_3361),
.D(n_3274),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3365),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3341),
.B(n_3244),
.Y(n_3386)
);

OR2x2_ASAP7_75t_L g3387 ( 
.A(n_3345),
.B(n_3310),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3324),
.B(n_3311),
.Y(n_3388)
);

NAND2x2_ASAP7_75t_L g3389 ( 
.A(n_3361),
.B(n_2939),
.Y(n_3389)
);

AOI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3343),
.A2(n_3260),
.B1(n_3170),
.B2(n_3150),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3377),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_3332),
.B(n_3311),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3326),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3376),
.B(n_3369),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3320),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3320),
.Y(n_3396)
);

OAI222xp33_ASAP7_75t_L g3397 ( 
.A1(n_3339),
.A2(n_3267),
.B1(n_3301),
.B2(n_3201),
.C1(n_3117),
.C2(n_3236),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3331),
.Y(n_3398)
);

INVx1_ASAP7_75t_SL g3399 ( 
.A(n_3363),
.Y(n_3399)
);

OAI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_3339),
.A2(n_3201),
.B1(n_3170),
.B2(n_3162),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3327),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3341),
.B(n_3244),
.Y(n_3402)
);

AOI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_3363),
.A2(n_3170),
.B1(n_2993),
.B2(n_3271),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3335),
.Y(n_3404)
);

INVx1_ASAP7_75t_SL g3405 ( 
.A(n_3322),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3337),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3338),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3327),
.Y(n_3408)
);

INVx1_ASAP7_75t_SL g3409 ( 
.A(n_3358),
.Y(n_3409)
);

OR2x2_ASAP7_75t_L g3410 ( 
.A(n_3364),
.B(n_3256),
.Y(n_3410)
);

OAI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3317),
.A2(n_2900),
.B(n_3201),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3353),
.Y(n_3412)
);

AOI32xp33_ASAP7_75t_L g3413 ( 
.A1(n_3330),
.A2(n_3162),
.A3(n_3133),
.B1(n_3286),
.B2(n_3302),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3340),
.Y(n_3414)
);

NAND4xp75_ASAP7_75t_SL g3415 ( 
.A(n_3359),
.B(n_3161),
.C(n_2981),
.D(n_3050),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3342),
.Y(n_3416)
);

NOR3xp33_ASAP7_75t_L g3417 ( 
.A(n_3317),
.B(n_2873),
.C(n_2882),
.Y(n_3417)
);

OAI22xp33_ASAP7_75t_L g3418 ( 
.A1(n_3347),
.A2(n_3201),
.B1(n_3133),
.B2(n_2945),
.Y(n_3418)
);

OAI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_3347),
.A2(n_3307),
.B1(n_3013),
.B2(n_3004),
.Y(n_3419)
);

OR3x2_ASAP7_75t_L g3420 ( 
.A(n_3348),
.B(n_2916),
.C(n_3218),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3359),
.A2(n_3286),
.B1(n_3308),
.B2(n_2957),
.Y(n_3421)
);

AOI22xp5_ASAP7_75t_L g3422 ( 
.A1(n_3355),
.A2(n_3291),
.B1(n_3169),
.B2(n_2980),
.Y(n_3422)
);

OAI22xp5_ASAP7_75t_L g3423 ( 
.A1(n_3344),
.A2(n_3334),
.B1(n_3321),
.B2(n_3329),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3346),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3349),
.A2(n_3265),
.B1(n_3264),
.B2(n_3298),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3356),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3362),
.Y(n_3427)
);

INVxp67_ASAP7_75t_L g3428 ( 
.A(n_3318),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3367),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3364),
.B(n_3256),
.Y(n_3430)
);

XOR2x2_ASAP7_75t_L g3431 ( 
.A(n_3417),
.B(n_3419),
.Y(n_3431)
);

AOI221xp5_ASAP7_75t_L g3432 ( 
.A1(n_3384),
.A2(n_3319),
.B1(n_3329),
.B2(n_3373),
.C(n_3371),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3420),
.A2(n_3389),
.B1(n_3403),
.B2(n_3383),
.Y(n_3433)
);

AOI22xp33_ASAP7_75t_L g3434 ( 
.A1(n_3383),
.A2(n_3265),
.B1(n_3264),
.B2(n_3302),
.Y(n_3434)
);

AOI21xp33_ASAP7_75t_L g3435 ( 
.A1(n_3382),
.A2(n_2886),
.B(n_2723),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3387),
.Y(n_3436)
);

AOI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3390),
.A2(n_3265),
.B1(n_3319),
.B2(n_3334),
.Y(n_3437)
);

NOR3xp33_ASAP7_75t_L g3438 ( 
.A(n_3397),
.B(n_2943),
.C(n_2924),
.Y(n_3438)
);

AOI221xp5_ASAP7_75t_L g3439 ( 
.A1(n_3423),
.A2(n_3405),
.B1(n_3399),
.B2(n_3428),
.C(n_3381),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3392),
.Y(n_3440)
);

OAI22xp33_ASAP7_75t_L g3441 ( 
.A1(n_3390),
.A2(n_3140),
.B1(n_3229),
.B2(n_3185),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3400),
.A2(n_3140),
.B(n_3229),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3394),
.B(n_3328),
.Y(n_3443)
);

NOR2xp33_ASAP7_75t_L g3444 ( 
.A(n_3409),
.B(n_3223),
.Y(n_3444)
);

AOI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3403),
.A2(n_3360),
.B1(n_3350),
.B2(n_3323),
.Y(n_3445)
);

OAI22xp5_ASAP7_75t_SL g3446 ( 
.A1(n_3422),
.A2(n_3223),
.B1(n_2926),
.B2(n_2930),
.Y(n_3446)
);

OAI21xp5_ASAP7_75t_SL g3447 ( 
.A1(n_3413),
.A2(n_3180),
.B(n_3104),
.Y(n_3447)
);

OAI21xp5_ASAP7_75t_L g3448 ( 
.A1(n_3422),
.A2(n_3124),
.B(n_3228),
.Y(n_3448)
);

OAI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3411),
.A2(n_3124),
.B(n_3235),
.Y(n_3449)
);

BUFx2_ASAP7_75t_SL g3450 ( 
.A(n_3421),
.Y(n_3450)
);

OAI221xp5_ASAP7_75t_SL g3451 ( 
.A1(n_3425),
.A2(n_3181),
.B1(n_3357),
.B2(n_3056),
.C(n_3299),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_3388),
.A2(n_3370),
.B1(n_3333),
.B2(n_2999),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3380),
.B(n_3285),
.Y(n_3453)
);

INVx1_ASAP7_75t_SL g3454 ( 
.A(n_3378),
.Y(n_3454)
);

OAI21xp33_ASAP7_75t_L g3455 ( 
.A1(n_3379),
.A2(n_3300),
.B(n_3299),
.Y(n_3455)
);

NOR3xp33_ASAP7_75t_L g3456 ( 
.A(n_3418),
.B(n_2944),
.C(n_2915),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3393),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3385),
.B(n_3300),
.Y(n_3458)
);

XOR2x2_ASAP7_75t_L g3459 ( 
.A(n_3415),
.B(n_2869),
.Y(n_3459)
);

INVx1_ASAP7_75t_SL g3460 ( 
.A(n_3398),
.Y(n_3460)
);

OAI21xp33_ASAP7_75t_L g3461 ( 
.A1(n_3386),
.A2(n_3297),
.B(n_3285),
.Y(n_3461)
);

NAND3xp33_ASAP7_75t_L g3462 ( 
.A(n_3404),
.B(n_2990),
.C(n_3083),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3406),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3402),
.B(n_3297),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3457),
.Y(n_3465)
);

NAND2xp33_ASAP7_75t_L g3466 ( 
.A(n_3438),
.B(n_2987),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_SL g3467 ( 
.A1(n_3450),
.A2(n_2884),
.B1(n_2876),
.B2(n_2894),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3454),
.B(n_3169),
.Y(n_3468)
);

OR2x2_ASAP7_75t_L g3469 ( 
.A(n_3458),
.B(n_3410),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3463),
.Y(n_3470)
);

OAI22xp33_ASAP7_75t_L g3471 ( 
.A1(n_3437),
.A2(n_3447),
.B1(n_3433),
.B2(n_3445),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3440),
.Y(n_3472)
);

INVxp67_ASAP7_75t_L g3473 ( 
.A(n_3446),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3460),
.Y(n_3474)
);

AOI221xp5_ASAP7_75t_L g3475 ( 
.A1(n_3432),
.A2(n_3424),
.B1(n_3429),
.B2(n_3427),
.C(n_3426),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3460),
.Y(n_3476)
);

OAI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3434),
.A2(n_3430),
.B1(n_3391),
.B2(n_3414),
.Y(n_3477)
);

AOI221xp5_ASAP7_75t_SL g3478 ( 
.A1(n_3439),
.A2(n_3448),
.B1(n_3435),
.B2(n_3441),
.C(n_3454),
.Y(n_3478)
);

INVx1_ASAP7_75t_SL g3479 ( 
.A(n_3431),
.Y(n_3479)
);

OAI21xp33_ASAP7_75t_L g3480 ( 
.A1(n_3451),
.A2(n_3407),
.B(n_3416),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3436),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3453),
.B(n_3395),
.Y(n_3482)
);

O2A1O1Ixp5_ASAP7_75t_L g3483 ( 
.A1(n_3444),
.A2(n_3401),
.B(n_3408),
.C(n_3396),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3464),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3455),
.B(n_3412),
.Y(n_3485)
);

OR2x2_ASAP7_75t_L g3486 ( 
.A(n_3461),
.B(n_3375),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3452),
.Y(n_3487)
);

OAI31xp33_ASAP7_75t_L g3488 ( 
.A1(n_3456),
.A2(n_2885),
.A3(n_2997),
.B(n_3104),
.Y(n_3488)
);

AOI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_3462),
.A2(n_3232),
.B1(n_3304),
.B2(n_3222),
.Y(n_3489)
);

OAI21xp33_ASAP7_75t_L g3490 ( 
.A1(n_3449),
.A2(n_3214),
.B(n_3316),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3443),
.B(n_3374),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3442),
.B(n_3316),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3459),
.B(n_3353),
.Y(n_3493)
);

NAND3xp33_ASAP7_75t_L g3494 ( 
.A(n_3433),
.B(n_3024),
.C(n_2677),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3432),
.B(n_3368),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3457),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3457),
.Y(n_3497)
);

INVx1_ASAP7_75t_SL g3498 ( 
.A(n_3460),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3450),
.B(n_3230),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3457),
.Y(n_3500)
);

AOI211xp5_ASAP7_75t_L g3501 ( 
.A1(n_3479),
.A2(n_2918),
.B(n_2906),
.C(n_3022),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3474),
.Y(n_3502)
);

AOI221xp5_ASAP7_75t_L g3503 ( 
.A1(n_3479),
.A2(n_3187),
.B1(n_3168),
.B2(n_3157),
.C(n_3167),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3476),
.Y(n_3504)
);

AND2x2_ASAP7_75t_L g3505 ( 
.A(n_3499),
.B(n_3203),
.Y(n_3505)
);

HB1xp67_ASAP7_75t_L g3506 ( 
.A(n_3498),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_L g3507 ( 
.A(n_3473),
.B(n_2950),
.Y(n_3507)
);

INVx1_ASAP7_75t_SL g3508 ( 
.A(n_3467),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3481),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_3487),
.B(n_2920),
.Y(n_3510)
);

NOR3xp33_ASAP7_75t_L g3511 ( 
.A(n_3471),
.B(n_2911),
.C(n_2868),
.Y(n_3511)
);

AOI221xp5_ASAP7_75t_L g3512 ( 
.A1(n_3478),
.A2(n_3168),
.B1(n_3157),
.B2(n_3123),
.C(n_3153),
.Y(n_3512)
);

NOR2x1_ASAP7_75t_L g3513 ( 
.A(n_3494),
.B(n_3028),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3468),
.B(n_3493),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_SL g3515 ( 
.A(n_3488),
.B(n_3061),
.Y(n_3515)
);

AOI211xp5_ASAP7_75t_L g3516 ( 
.A1(n_3478),
.A2(n_3466),
.B(n_3480),
.C(n_3477),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_3483),
.B(n_3066),
.Y(n_3517)
);

NOR3xp33_ASAP7_75t_L g3518 ( 
.A(n_3498),
.B(n_2961),
.C(n_2953),
.Y(n_3518)
);

NAND3xp33_ASAP7_75t_L g3519 ( 
.A(n_3475),
.B(n_3055),
.C(n_3064),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3484),
.B(n_2922),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3495),
.A2(n_2676),
.B(n_3028),
.Y(n_3521)
);

NOR2x1_ASAP7_75t_L g3522 ( 
.A(n_3465),
.B(n_3082),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3470),
.B(n_3368),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3472),
.B(n_3372),
.Y(n_3524)
);

NOR3x1_ASAP7_75t_L g3525 ( 
.A(n_3492),
.B(n_3076),
.C(n_3065),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3508),
.B(n_3496),
.Y(n_3526)
);

AOI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3511),
.A2(n_3489),
.B1(n_3490),
.B2(n_3500),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3517),
.A2(n_3497),
.B(n_3485),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3506),
.B(n_3469),
.Y(n_3529)
);

AOI21xp5_ASAP7_75t_L g3530 ( 
.A1(n_3515),
.A2(n_3491),
.B(n_3486),
.Y(n_3530)
);

AOI211x1_ASAP7_75t_L g3531 ( 
.A1(n_3521),
.A2(n_3502),
.B(n_3504),
.C(n_3516),
.Y(n_3531)
);

OA22x2_ASAP7_75t_L g3532 ( 
.A1(n_3509),
.A2(n_3513),
.B1(n_3525),
.B2(n_3523),
.Y(n_3532)
);

AOI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3514),
.A2(n_3482),
.B1(n_3121),
.B2(n_2963),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3503),
.B(n_3372),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3510),
.Y(n_3535)
);

NAND2x1_ASAP7_75t_L g3536 ( 
.A(n_3522),
.B(n_3099),
.Y(n_3536)
);

AOI221x1_ASAP7_75t_SL g3537 ( 
.A1(n_3507),
.A2(n_2750),
.B1(n_3079),
.B2(n_3196),
.C(n_3191),
.Y(n_3537)
);

AOI211x1_ASAP7_75t_L g3538 ( 
.A1(n_3519),
.A2(n_3174),
.B(n_3176),
.C(n_2676),
.Y(n_3538)
);

NOR3x1_ASAP7_75t_L g3539 ( 
.A(n_3501),
.B(n_3523),
.C(n_3520),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3524),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3512),
.A2(n_3067),
.B(n_3180),
.Y(n_3541)
);

OA22x2_ASAP7_75t_L g3542 ( 
.A1(n_3505),
.A2(n_3191),
.B1(n_3002),
.B2(n_3031),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3518),
.B(n_3336),
.Y(n_3543)
);

AOI211xp5_ASAP7_75t_L g3544 ( 
.A1(n_3508),
.A2(n_2949),
.B(n_2932),
.C(n_3062),
.Y(n_3544)
);

OAI22xp5_ASAP7_75t_L g3545 ( 
.A1(n_3516),
.A2(n_2956),
.B1(n_3351),
.B2(n_3196),
.Y(n_3545)
);

AOI222xp33_ASAP7_75t_L g3546 ( 
.A1(n_3526),
.A2(n_2652),
.B1(n_2693),
.B2(n_3138),
.C1(n_3219),
.C2(n_3200),
.Y(n_3546)
);

AOI211xp5_ASAP7_75t_L g3547 ( 
.A1(n_3545),
.A2(n_2698),
.B(n_3086),
.C(n_3090),
.Y(n_3547)
);

OAI21xp5_ASAP7_75t_SL g3548 ( 
.A1(n_3535),
.A2(n_2985),
.B(n_2721),
.Y(n_3548)
);

NAND4xp25_ASAP7_75t_L g3549 ( 
.A(n_3531),
.B(n_3046),
.C(n_2978),
.D(n_2968),
.Y(n_3549)
);

OAI22xp33_ASAP7_75t_L g3550 ( 
.A1(n_3532),
.A2(n_3033),
.B1(n_3276),
.B2(n_3095),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_3544),
.B(n_3530),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3537),
.B(n_3105),
.Y(n_3552)
);

OAI211xp5_ASAP7_75t_SL g3553 ( 
.A1(n_3528),
.A2(n_2761),
.B(n_2786),
.C(n_2777),
.Y(n_3553)
);

NAND3xp33_ASAP7_75t_L g3554 ( 
.A(n_3538),
.B(n_2777),
.C(n_2766),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3529),
.B(n_3102),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3540),
.B(n_3134),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3527),
.B(n_3543),
.Y(n_3557)
);

O2A1O1Ixp33_ASAP7_75t_SL g3558 ( 
.A1(n_3536),
.A2(n_3534),
.B(n_3539),
.C(n_3533),
.Y(n_3558)
);

NOR3x1_ASAP7_75t_L g3559 ( 
.A(n_3542),
.B(n_2436),
.C(n_2449),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3541),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3526),
.A2(n_3216),
.B(n_3075),
.Y(n_3561)
);

NOR3xp33_ASAP7_75t_L g3562 ( 
.A(n_3551),
.B(n_3553),
.C(n_3550),
.Y(n_3562)
);

NOR2x1_ASAP7_75t_L g3563 ( 
.A(n_3560),
.B(n_2443),
.Y(n_3563)
);

OR2x6_ASAP7_75t_L g3564 ( 
.A(n_3548),
.B(n_3089),
.Y(n_3564)
);

AOI22xp5_ASAP7_75t_L g3565 ( 
.A1(n_3557),
.A2(n_3121),
.B1(n_3190),
.B2(n_3068),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3546),
.B(n_3552),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3555),
.Y(n_3567)
);

AND2x4_ASAP7_75t_L g3568 ( 
.A(n_3554),
.B(n_3156),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3556),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_L g3570 ( 
.A(n_3558),
.B(n_2766),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3561),
.B(n_3559),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_3547),
.A2(n_3315),
.B1(n_3309),
.B2(n_3287),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_3549),
.Y(n_3573)
);

NAND4xp25_ASAP7_75t_L g3574 ( 
.A(n_3562),
.B(n_2786),
.C(n_2812),
.D(n_3096),
.Y(n_3574)
);

NOR2x1_ASAP7_75t_L g3575 ( 
.A(n_3573),
.B(n_2333),
.Y(n_3575)
);

NAND2x1_ASAP7_75t_L g3576 ( 
.A(n_3570),
.B(n_2812),
.Y(n_3576)
);

INVxp67_ASAP7_75t_L g3577 ( 
.A(n_3571),
.Y(n_3577)
);

NAND4xp75_ASAP7_75t_L g3578 ( 
.A(n_3566),
.B(n_3161),
.C(n_2800),
.D(n_3217),
.Y(n_3578)
);

NOR3xp33_ASAP7_75t_L g3579 ( 
.A(n_3567),
.B(n_2499),
.C(n_2461),
.Y(n_3579)
);

AND3x4_ASAP7_75t_L g3580 ( 
.A(n_3563),
.B(n_3069),
.C(n_3080),
.Y(n_3580)
);

NOR2xp33_ASAP7_75t_R g3581 ( 
.A(n_3569),
.B(n_3021),
.Y(n_3581)
);

NOR3xp33_ASAP7_75t_L g3582 ( 
.A(n_3565),
.B(n_2470),
.C(n_2463),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3577),
.B(n_3568),
.Y(n_3583)
);

XOR2xp5_ASAP7_75t_L g3584 ( 
.A(n_3574),
.B(n_3572),
.Y(n_3584)
);

AND2x4_ASAP7_75t_L g3585 ( 
.A(n_3576),
.B(n_3564),
.Y(n_3585)
);

BUFx12f_ASAP7_75t_L g3586 ( 
.A(n_3581),
.Y(n_3586)
);

INVx1_ASAP7_75t_SL g3587 ( 
.A(n_3575),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3583),
.Y(n_3588)
);

AOI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_3588),
.A2(n_3586),
.B1(n_3585),
.B2(n_3584),
.Y(n_3589)
);

XNOR2xp5_ASAP7_75t_L g3590 ( 
.A(n_3589),
.B(n_3587),
.Y(n_3590)
);

O2A1O1Ixp33_ASAP7_75t_L g3591 ( 
.A1(n_3590),
.A2(n_3564),
.B(n_3582),
.C(n_3579),
.Y(n_3591)
);

XNOR2xp5_ASAP7_75t_L g3592 ( 
.A(n_3591),
.B(n_3578),
.Y(n_3592)
);

AOI222xp33_ASAP7_75t_L g3593 ( 
.A1(n_3592),
.A2(n_3580),
.B1(n_3276),
.B2(n_2566),
.C1(n_2475),
.C2(n_2472),
.Y(n_3593)
);

OR2x6_ASAP7_75t_L g3594 ( 
.A(n_3593),
.B(n_3021),
.Y(n_3594)
);

AOI22xp33_ASAP7_75t_L g3595 ( 
.A1(n_3594),
.A2(n_3276),
.B1(n_3021),
.B2(n_3044),
.Y(n_3595)
);


endmodule