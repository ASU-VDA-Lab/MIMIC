module real_jpeg_4527_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_213;
wire n_179;
wire n_128;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.C(n_35),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_43),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_35),
.B1(n_43),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_43),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_56),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_191),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_196),
.B(n_198),
.C(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_209),
.C(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_2),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_2),
.B(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_5),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_13)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_11),
.A2(n_115),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_12),
.Y(n_134)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_168),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_167),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_150),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_150),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_104),
.C(n_144),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_25),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_53),
.B2(n_54),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_27),
.A2(n_77),
.B(n_146),
.C(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_28),
.A2(n_29),
.B1(n_38),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_36),
.A2(n_80),
.B1(n_84),
.B2(n_86),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_37),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_38),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_38),
.B(n_147),
.C(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_38),
.A2(n_176),
.B1(n_195),
.B2(n_202),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_38),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_38),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_38),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_38),
.B(n_195),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_43),
.A2(n_90),
.B(n_93),
.Y(n_198)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_49),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_49),
.A2(n_109),
.B1(n_156),
.B2(n_160),
.Y(n_155)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_51),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_54),
.B(n_166),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_77),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_55),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_55),
.B(n_118),
.Y(n_149)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_55),
.A2(n_152),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_65),
.B(n_74),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_66),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_77),
.A2(n_117),
.B1(n_118),
.B2(n_147),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_77),
.A2(n_147),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

AO21x2_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_101),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

OA22x2_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_104),
.A2(n_144),
.B1(n_145),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_117),
.B1(n_118),
.B2(n_143),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_118),
.Y(n_166)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_118),
.B1(n_155),
.B2(n_164),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_117),
.B(n_176),
.C(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_117),
.A2(n_118),
.B1(n_190),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_117),
.A2(n_118),
.B1(n_206),
.B2(n_207),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_117),
.A2(n_118),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_117),
.B(n_232),
.C(n_237),
.Y(n_242)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_118),
.B(n_206),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_118),
.A2(n_147),
.B(n_194),
.C(n_239),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.Y(n_118)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_121),
.Y(n_211)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.Y(n_125)
);

NAND2x1_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_126),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_134),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_127),
.B(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_142),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AND3x1_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_149),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_165),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_183),
.B(n_247),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_170),
.B(n_180),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_173),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_176),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_241),
.B(n_246),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_230),
.B(n_240),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_203),
.B(n_229),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_215),
.B(n_228),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_212),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_238),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);


endmodule