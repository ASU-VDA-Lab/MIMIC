module fake_netlist_6_1675_n_1755 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1755);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1755;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_75),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_36),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_68),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_88),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_73),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_51),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_62),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_30),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_49),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_14),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_74),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_58),
.Y(n_178)
);

BUFx2_ASAP7_75t_SL g179 ( 
.A(n_119),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_41),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_91),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_70),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_103),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_64),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_10),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_56),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_67),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_118),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_112),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_50),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_65),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_38),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_138),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_153),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_96),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_85),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_34),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_59),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_9),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_139),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_50),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_122),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_12),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_47),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_98),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_18),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_126),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_108),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_8),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_20),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_151),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_149),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_80),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_53),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_76),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_3),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_12),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_63),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_69),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_142),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_89),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_127),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_46),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_100),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_21),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_147),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_41),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_106),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_39),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_97),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_44),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_116),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_60),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_158),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_5),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_133),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_31),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_84),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_156),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_46),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_150),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_24),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_37),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_0),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_49),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_55),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_102),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_154),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_31),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_130),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_82),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_90),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_48),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_20),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_22),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_25),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_40),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_87),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_5),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_61),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_21),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_22),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_9),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_2),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_28),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_39),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_131),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_86),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_23),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_30),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_18),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_77),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_105),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_78),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_2),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_R g318 ( 
.A(n_165),
.B(n_113),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_201),
.B(n_0),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_199),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_206),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_164),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_238),
.B(n_1),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_208),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_214),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_215),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_217),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_196),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_216),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_180),
.B(n_238),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_1),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_195),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_226),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_244),
.B(n_4),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_221),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_243),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_241),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_193),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_243),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_4),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_242),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_164),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_245),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_172),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_317),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_162),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_213),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_250),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_248),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_218),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_247),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_314),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_290),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_249),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_256),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_222),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_265),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_266),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_267),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_271),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_211),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_233),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_185),
.B(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_236),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_251),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_311),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_272),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_273),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_276),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_288),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_262),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_293),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_275),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_204),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_212),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_285),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_224),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_323),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_202),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_325),
.B(n_160),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_322),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_163),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_320),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_333),
.B(n_163),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_389),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_336),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_330),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_166),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_324),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_331),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_185),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_344),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_353),
.B(n_231),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_344),
.B(n_166),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_347),
.Y(n_428)
);

CKINVDCx6p67_ASAP7_75t_R g429 ( 
.A(n_349),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_354),
.B(n_168),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_332),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_334),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_354),
.B(n_168),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_257),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_359),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_338),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_329),
.B(n_161),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_346),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_355),
.B(n_170),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_342),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_348),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_361),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_352),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_363),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_356),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_368),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_369),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_R g457 ( 
.A(n_391),
.B(n_170),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_371),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_370),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_R g463 ( 
.A(n_380),
.B(n_169),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_372),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_376),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_360),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_257),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_421),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_430),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_409),
.B(n_349),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_411),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_337),
.B1(n_362),
.B2(n_387),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_411),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_362),
.B1(n_384),
.B2(n_382),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_341),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_403),
.B(n_373),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_409),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_374),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_430),
.B(n_383),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_430),
.B(n_403),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_385),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_431),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_441),
.Y(n_488)
);

BUFx4_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_345),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_413),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_375),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

NOR2x1p5_ASAP7_75t_L g497 ( 
.A(n_429),
.B(n_340),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_447),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_423),
.A2(n_351),
.B1(n_437),
.B2(n_425),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_446),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_402),
.B(n_419),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_423),
.A2(n_261),
.B1(n_289),
.B2(n_296),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_408),
.B(n_223),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_423),
.A2(n_261),
.B1(n_289),
.B2(n_312),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_420),
.B(n_269),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_425),
.B(n_356),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_420),
.B(n_179),
.Y(n_509)
);

AND2x2_ASAP7_75t_SL g510 ( 
.A(n_415),
.B(n_202),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_432),
.B(n_318),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_425),
.B(n_202),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_448),
.Y(n_516)
);

INVx4_ASAP7_75t_SL g517 ( 
.A(n_414),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_357),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_426),
.B(n_167),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_437),
.B(n_357),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_437),
.B(n_378),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_426),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_458),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_460),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_432),
.B(n_202),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_400),
.B(n_178),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_457),
.B(n_202),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_462),
.A2(n_381),
.B1(n_390),
.B2(n_388),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_457),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_436),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_400),
.B(n_189),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_378),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_394),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_436),
.B(n_444),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_397),
.B(n_379),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_397),
.B(n_379),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_460),
.B(n_263),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_462),
.A2(n_392),
.B1(n_390),
.B2(n_388),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_395),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_395),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_434),
.Y(n_552)
);

OAI21xp33_ASAP7_75t_SL g553 ( 
.A1(n_444),
.A2(n_392),
.B(n_386),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_443),
.B(n_367),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_396),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_414),
.B(n_381),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_460),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_416),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_396),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_416),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_462),
.A2(n_386),
.B1(n_263),
.B2(n_310),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_429),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_462),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_451),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_416),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_429),
.B(n_198),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_460),
.B(n_263),
.Y(n_571)
);

AND3x1_ASAP7_75t_L g572 ( 
.A(n_463),
.B(n_197),
.C(n_315),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_400),
.B(n_200),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_400),
.B(n_227),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_454),
.B(n_456),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_399),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_406),
.Y(n_578)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_439),
.B(n_230),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_463),
.A2(n_292),
.B1(n_203),
.B2(n_207),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_404),
.B(n_209),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_416),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_406),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_459),
.B(n_171),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_404),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_407),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_460),
.B(n_263),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_464),
.B(n_171),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_406),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_439),
.A2(n_263),
.B1(n_210),
.B2(n_254),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_439),
.B(n_449),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_407),
.B(n_219),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_460),
.B(n_229),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_449),
.A2(n_232),
.B1(n_252),
.B2(n_246),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_410),
.B(n_176),
.Y(n_595)
);

AOI21x1_ASAP7_75t_L g596 ( 
.A1(n_401),
.A2(n_240),
.B(n_237),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_416),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_449),
.A2(n_277),
.B1(n_259),
.B2(n_279),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_410),
.B(n_176),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_412),
.B(n_177),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_412),
.B(n_177),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_417),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_417),
.B(n_181),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_401),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_424),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_424),
.B(n_181),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_453),
.B(n_183),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_424),
.B(n_183),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_435),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_453),
.B(n_270),
.C(n_260),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_424),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_453),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_435),
.B(n_184),
.Y(n_613)
);

AO22x2_ASAP7_75t_L g614 ( 
.A1(n_455),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_406),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_455),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_SL g617 ( 
.A(n_530),
.B(n_184),
.Y(n_617)
);

AND2x6_ASAP7_75t_SL g618 ( 
.A(n_480),
.B(n_220),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_543),
.A2(n_304),
.B1(n_286),
.B2(n_225),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_578),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_543),
.B(n_435),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_481),
.B(n_435),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_578),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_485),
.A2(n_455),
.B(n_405),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_481),
.B(n_435),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_475),
.A2(n_175),
.B1(n_174),
.B2(n_173),
.C(n_313),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_536),
.B(n_435),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_467),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_583),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_502),
.B(n_435),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_591),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_502),
.B(n_427),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_523),
.B(n_186),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_523),
.B(n_427),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_504),
.A2(n_305),
.B1(n_173),
.B2(n_174),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_466),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_485),
.A2(n_553),
.B(n_519),
.C(n_505),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_482),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_472),
.B(n_405),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_510),
.A2(n_365),
.B1(n_366),
.B2(n_239),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_495),
.B(n_427),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_477),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_507),
.B(n_186),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_482),
.B(n_428),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_510),
.B(n_187),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_499),
.A2(n_484),
.B1(n_486),
.B2(n_483),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_518),
.B(n_428),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_583),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_504),
.A2(n_175),
.B(n_313),
.C(n_307),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_472),
.B(n_509),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_499),
.B(n_616),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_530),
.A2(n_438),
.B(n_428),
.C(n_405),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_487),
.B(n_438),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_568),
.B(n_438),
.Y(n_655)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_584),
.B(n_187),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_591),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_L g658 ( 
.A(n_584),
.B(n_188),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_468),
.B(n_188),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_567),
.B(n_191),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_479),
.A2(n_182),
.B1(n_306),
.B2(n_303),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_506),
.A2(n_169),
.B1(n_182),
.B2(n_307),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_491),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_511),
.A2(n_572),
.B1(n_473),
.B2(n_580),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_567),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_589),
.Y(n_666)
);

NAND2x1p5_ASAP7_75t_L g667 ( 
.A(n_525),
.B(n_405),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_493),
.B(n_405),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_522),
.B(n_191),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_613),
.A2(n_309),
.B(n_192),
.C(n_194),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_580),
.A2(n_309),
.B1(n_192),
.B2(n_194),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_588),
.B(n_294),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_588),
.B(n_294),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_471),
.B(n_280),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_496),
.B(n_239),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_500),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_471),
.B(n_281),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_605),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_503),
.B(n_235),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_522),
.B(n_235),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_516),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_469),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_470),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_605),
.B(n_300),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_520),
.B(n_526),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_SL g686 ( 
.A1(n_575),
.A2(n_306),
.B1(n_303),
.B2(n_234),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_531),
.B(n_302),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_539),
.B(n_302),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_589),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_529),
.B(n_300),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_552),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_600),
.B(n_274),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_601),
.B(n_268),
.Y(n_693)
);

INVx8_ASAP7_75t_L g694 ( 
.A(n_480),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_538),
.B(n_205),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_610),
.B(n_92),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_558),
.B(n_278),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_81),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_579),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_534),
.B(n_264),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_558),
.B(n_282),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_540),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_542),
.B(n_253),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_525),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_506),
.A2(n_287),
.B1(n_258),
.B2(n_291),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_468),
.B(n_301),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_508),
.Y(n_707)
);

OAI221xp5_ASAP7_75t_L g708 ( 
.A1(n_594),
.A2(n_301),
.B1(n_299),
.B2(n_297),
.C(n_295),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_545),
.B(n_205),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_546),
.B(n_299),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_550),
.B(n_205),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_546),
.B(n_297),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_551),
.B(n_195),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_580),
.A2(n_295),
.B1(n_234),
.B2(n_190),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_614),
.A2(n_190),
.B1(n_195),
.B2(n_14),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_469),
.Y(n_716)
);

OAI221xp5_ASAP7_75t_L g717 ( 
.A1(n_594),
.A2(n_6),
.B1(n_13),
.B2(n_15),
.C(n_16),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_614),
.A2(n_13),
.B1(n_17),
.B2(n_19),
.C(n_23),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_540),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_474),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_556),
.B(n_152),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_582),
.A2(n_145),
.B(n_140),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_546),
.B(n_17),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_563),
.B(n_137),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_492),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_573),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_574),
.B(n_135),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_614),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_615),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_492),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_577),
.B(n_129),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_547),
.B(n_27),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_585),
.B(n_123),
.Y(n_733)
);

AOI221xp5_ASAP7_75t_L g734 ( 
.A1(n_598),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_33),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_SL g735 ( 
.A(n_501),
.B(n_29),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_508),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_521),
.B(n_107),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_547),
.B(n_33),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_586),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_602),
.B(n_99),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_480),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_607),
.B(n_604),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_607),
.B(n_94),
.Y(n_743)
);

INVx8_ASAP7_75t_L g744 ( 
.A(n_490),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_547),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_521),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_490),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_595),
.B(n_35),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_606),
.B(n_66),
.Y(n_749)
);

BUFx8_ASAP7_75t_L g750 ( 
.A(n_555),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_474),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_611),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_615),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_478),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_492),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_490),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_608),
.B(n_35),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_478),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_492),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_595),
.B(n_52),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_612),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_494),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_527),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_599),
.B(n_52),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_565),
.B(n_560),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_565),
.B(n_37),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_532),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_599),
.B(n_38),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_532),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_470),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_603),
.B(n_40),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_494),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_590),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_42),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_488),
.B(n_48),
.C(n_51),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_512),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_566),
.B(n_497),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_576),
.B(n_613),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_590),
.B(n_564),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_544),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_533),
.B(n_549),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_581),
.B(n_592),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_554),
.B(n_569),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_544),
.A2(n_557),
.B1(n_512),
.B2(n_513),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_533),
.A2(n_549),
.B(n_598),
.C(n_528),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_527),
.B(n_560),
.Y(n_786)
);

AO22x1_ASAP7_75t_L g787 ( 
.A1(n_468),
.A2(n_515),
.B1(n_557),
.B2(n_513),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_498),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_527),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_782),
.B(n_554),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_665),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_782),
.B(n_569),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_645),
.B(n_541),
.Y(n_793)
);

O2A1O1Ixp5_ASAP7_75t_L g794 ( 
.A1(n_748),
.A2(n_593),
.B(n_571),
.C(n_548),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_637),
.B(n_561),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_648),
.B(n_564),
.Y(n_796)
);

AND2x2_ASAP7_75t_SL g797 ( 
.A(n_735),
.B(n_489),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_622),
.A2(n_535),
.B(n_537),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_625),
.A2(n_535),
.B(n_537),
.Y(n_799)
);

NOR2x1_ASAP7_75t_L g800 ( 
.A(n_777),
.B(n_498),
.Y(n_800)
);

INVx11_ASAP7_75t_L g801 ( 
.A(n_750),
.Y(n_801)
);

AOI22x1_ASAP7_75t_L g802 ( 
.A1(n_628),
.A2(n_514),
.B1(n_560),
.B2(n_527),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_644),
.B(n_514),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_621),
.A2(n_562),
.B(n_560),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_651),
.A2(n_562),
.B(n_597),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_647),
.A2(n_593),
.B(n_571),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_748),
.A2(n_587),
.B(n_548),
.C(n_597),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_639),
.B(n_524),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_468),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_672),
.B(n_524),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_638),
.A2(n_652),
.B(n_785),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_715),
.A2(n_728),
.B1(n_781),
.B2(n_773),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_631),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_665),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_768),
.A2(n_587),
.B(n_597),
.C(n_468),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_630),
.B(n_515),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_715),
.A2(n_596),
.B1(n_597),
.B2(n_559),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_742),
.B(n_515),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_642),
.A2(n_559),
.B(n_609),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_665),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_672),
.B(n_673),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_765),
.A2(n_559),
.B(n_609),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_778),
.B(n_541),
.Y(n_823)
);

BUFx8_ASAP7_75t_L g824 ( 
.A(n_683),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_765),
.A2(n_559),
.B(n_517),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_785),
.A2(n_515),
.B(n_517),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_778),
.B(n_561),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_779),
.A2(n_517),
.B(n_515),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_745),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_674),
.B(n_677),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_783),
.A2(n_627),
.B(n_786),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_664),
.B(n_702),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_673),
.B(n_692),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_692),
.B(n_693),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_728),
.A2(n_773),
.B1(n_619),
.B2(n_768),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_786),
.A2(n_730),
.B(n_725),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_619),
.B(n_626),
.C(n_633),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_760),
.A2(n_771),
.B1(n_764),
.B2(n_774),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_743),
.A2(n_646),
.B(n_737),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_694),
.B(n_741),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_725),
.A2(n_730),
.B(n_640),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_640),
.A2(n_657),
.B(n_685),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_693),
.B(n_632),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_717),
.A2(n_650),
.B(n_766),
.C(n_737),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_700),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_641),
.B(n_699),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_691),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_650),
.A2(n_766),
.B(n_646),
.C(n_634),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_663),
.B(n_676),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_681),
.B(n_726),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_714),
.A2(n_718),
.B1(n_635),
.B2(n_671),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_688),
.A2(n_698),
.B(n_670),
.C(n_757),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_657),
.A2(n_736),
.B1(n_719),
.B2(n_746),
.Y(n_853)
);

OA22x2_ASAP7_75t_L g854 ( 
.A1(n_738),
.A2(n_747),
.B1(n_756),
.B2(n_695),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_755),
.A2(n_763),
.B(n_759),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_723),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_739),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_755),
.A2(n_763),
.B(n_759),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_755),
.A2(n_763),
.B(n_759),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_707),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_755),
.B(n_759),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_678),
.B(n_656),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_678),
.B(n_658),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_636),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_763),
.A2(n_729),
.B(n_753),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_729),
.A2(n_753),
.B(n_749),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_643),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_789),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_688),
.A2(n_752),
.B(n_710),
.C(n_712),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_710),
.A2(n_712),
.B(n_707),
.C(n_761),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_695),
.A2(n_697),
.B1(n_701),
.B2(n_690),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_624),
.A2(n_704),
.B(n_789),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_654),
.A2(n_723),
.B(n_732),
.C(n_703),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_669),
.B(n_680),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_635),
.B(n_714),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_732),
.A2(n_655),
.B(n_690),
.C(n_713),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_704),
.A2(n_667),
.B(n_727),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_744),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_667),
.A2(n_727),
.B(n_668),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_682),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_787),
.A2(n_784),
.B(n_724),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_767),
.A2(n_780),
.B(n_769),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_669),
.B(n_680),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_686),
.B(n_687),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_662),
.B(n_661),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_776),
.B(n_682),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_772),
.B(n_733),
.Y(n_887)
);

O2A1O1Ixp5_ASAP7_75t_L g888 ( 
.A1(n_617),
.A2(n_784),
.B(n_687),
.C(n_684),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_721),
.A2(n_731),
.B(n_740),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_620),
.A2(n_689),
.B(n_623),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_776),
.B(n_772),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_675),
.B(n_679),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_716),
.B(n_762),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_662),
.B(n_709),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_660),
.B(n_684),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_629),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_649),
.A2(n_666),
.B(n_751),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_720),
.B(n_758),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_744),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_770),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_754),
.A2(n_659),
.B(n_660),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_744),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_711),
.B(n_788),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_694),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_653),
.A2(n_706),
.B(n_722),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_694),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_741),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_708),
.B(n_705),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_696),
.B(n_734),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_775),
.B(n_741),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_750),
.B(n_618),
.Y(n_911)
);

BUFx2_ASAP7_75t_R g912 ( 
.A(n_691),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_631),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_665),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_715),
.A2(n_728),
.B1(n_781),
.B2(n_773),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_787),
.A2(n_485),
.B(n_786),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_652),
.A2(n_646),
.B1(n_647),
.B2(n_621),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_622),
.A2(n_472),
.B(n_625),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_748),
.A2(n_768),
.B(n_543),
.C(n_638),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_647),
.A2(n_621),
.B(n_638),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_715),
.A2(n_728),
.B1(n_781),
.B2(n_773),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_635),
.A2(n_442),
.B(n_339),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_631),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_748),
.A2(n_768),
.B(n_652),
.C(n_764),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_782),
.B(n_543),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_707),
.B(n_736),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_622),
.A2(n_472),
.B(n_625),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_624),
.A2(n_640),
.B(n_783),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_622),
.A2(n_472),
.B(n_625),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_674),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_665),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_748),
.A2(n_768),
.B(n_652),
.C(n_764),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_631),
.Y(n_933)
);

BUFx10_ASAP7_75t_L g934 ( 
.A(n_691),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_622),
.A2(n_472),
.B(n_625),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_778),
.A2(n_543),
.B1(n_782),
.B2(n_481),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_631),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_631),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_782),
.B(n_543),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_SL g940 ( 
.A1(n_743),
.A2(n_785),
.B(n_766),
.C(n_737),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_782),
.B(n_543),
.Y(n_941)
);

CKINVDCx10_ASAP7_75t_R g942 ( 
.A(n_770),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_778),
.A2(n_543),
.B1(n_782),
.B2(n_481),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_778),
.B(n_510),
.Y(n_944)
);

INVx11_ASAP7_75t_L g945 ( 
.A(n_750),
.Y(n_945)
);

NOR2xp67_ASAP7_75t_L g946 ( 
.A(n_691),
.B(n_568),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_637),
.B(n_360),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_744),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_715),
.A2(n_728),
.B1(n_781),
.B2(n_773),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_782),
.B(n_543),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_782),
.B(n_543),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_637),
.B(n_360),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_782),
.B(n_543),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_672),
.B(n_673),
.C(n_619),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_782),
.B(n_543),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_631),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_782),
.B(n_543),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_647),
.A2(n_621),
.B(n_638),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_647),
.A2(n_621),
.B(n_638),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_637),
.B(n_360),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_622),
.A2(n_472),
.B(n_625),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_631),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_652),
.A2(n_646),
.B1(n_647),
.B2(n_621),
.Y(n_963)
);

AOI22x1_ASAP7_75t_L g964 ( 
.A1(n_628),
.A2(n_523),
.B1(n_502),
.B2(n_636),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_637),
.B(n_360),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_782),
.B(n_543),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_665),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_782),
.B(n_543),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_645),
.B(n_518),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_652),
.A2(n_646),
.B1(n_647),
.B2(n_621),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_635),
.A2(n_442),
.B(n_339),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_782),
.B(n_543),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_782),
.B(n_543),
.Y(n_973)
);

AOI21xp33_ASAP7_75t_L g974 ( 
.A1(n_672),
.A2(n_673),
.B(n_646),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_L g975 ( 
.A1(n_748),
.A2(n_485),
.B(n_768),
.C(n_543),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_631),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_631),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_748),
.A2(n_768),
.B1(n_764),
.B2(n_760),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_814),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_974),
.A2(n_833),
.B(n_954),
.C(n_834),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_821),
.A2(n_835),
.B1(n_936),
.B2(n_943),
.Y(n_981)
);

OA21x2_ASAP7_75t_L g982 ( 
.A1(n_811),
.A2(n_958),
.B(n_920),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_SL g983 ( 
.A(n_812),
.B(n_915),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_793),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_829),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_925),
.B(n_939),
.Y(n_986)
);

OR2x6_ASAP7_75t_L g987 ( 
.A(n_840),
.B(n_878),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_918),
.A2(n_929),
.B(n_927),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_941),
.B(n_950),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_935),
.A2(n_961),
.B(n_803),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_835),
.A2(n_812),
.B1(n_915),
.B2(n_921),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_824),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_798),
.A2(n_799),
.B(n_877),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_866),
.A2(n_872),
.B(n_879),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_824),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_951),
.A2(n_968),
.B1(n_973),
.B2(n_972),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_953),
.B(n_955),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_805),
.A2(n_822),
.B(n_842),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_814),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_861),
.A2(n_889),
.B(n_940),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_904),
.B(n_906),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_790),
.A2(n_792),
.B(n_957),
.Y(n_1003)
);

AO31x2_ASAP7_75t_L g1004 ( 
.A1(n_919),
.A2(n_839),
.A3(n_963),
.B(n_970),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_966),
.A2(n_841),
.B(n_796),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_908),
.A2(n_837),
.B1(n_949),
.B2(n_921),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_811),
.A2(n_958),
.B(n_920),
.Y(n_1007)
);

AOI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_924),
.A2(n_932),
.B(n_949),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_826),
.A2(n_802),
.B(n_836),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_826),
.A2(n_901),
.B(n_881),
.Y(n_1010)
);

NAND3x1_ASAP7_75t_L g1011 ( 
.A(n_875),
.B(n_885),
.C(n_911),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_959),
.A2(n_917),
.B(n_975),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_813),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_843),
.B(n_969),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_SL g1015 ( 
.A1(n_844),
.A2(n_848),
.B(n_858),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_933),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_830),
.B(n_856),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_SL g1018 ( 
.A1(n_855),
.A2(n_859),
.B(n_862),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_865),
.A2(n_959),
.B(n_816),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_825),
.A2(n_905),
.B(n_890),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_863),
.A2(n_905),
.B(n_828),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_806),
.A2(n_892),
.B(n_819),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_937),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_806),
.A2(n_794),
.B(n_978),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_944),
.A2(n_873),
.B(n_888),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_874),
.A2(n_895),
.B(n_971),
.C(n_922),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_942),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_897),
.A2(n_868),
.B(n_891),
.Y(n_1028)
);

INVx6_ASAP7_75t_L g1029 ( 
.A(n_934),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_818),
.A2(n_852),
.B(n_815),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_869),
.A2(n_909),
.B(n_810),
.C(n_894),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_SL g1032 ( 
.A(n_814),
.B(n_820),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_947),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_838),
.A2(n_807),
.B(n_870),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_886),
.A2(n_849),
.B(n_850),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_952),
.B(n_960),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_880),
.A2(n_838),
.B(n_817),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_876),
.A2(n_893),
.B(n_898),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_965),
.B(n_930),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_817),
.A2(n_884),
.A3(n_851),
.B(n_976),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_SL g1041 ( 
.A1(n_851),
.A2(n_964),
.B(n_871),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_883),
.A2(n_846),
.B(n_853),
.C(n_845),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_931),
.A2(n_977),
.B(n_962),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_832),
.B(n_857),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_832),
.B(n_923),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_913),
.A2(n_956),
.B(n_938),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_864),
.A2(n_867),
.A3(n_903),
.B(n_791),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_912),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_832),
.B(n_896),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_820),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_854),
.A2(n_823),
.B(n_827),
.Y(n_1051)
);

OA21x2_ASAP7_75t_L g1052 ( 
.A1(n_910),
.A2(n_926),
.B(n_887),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_832),
.B(n_926),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_967),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_791),
.A2(n_967),
.B(n_914),
.Y(n_1055)
);

INVx4_ASAP7_75t_L g1056 ( 
.A(n_820),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_967),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_860),
.B(n_914),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_860),
.B(n_914),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_900),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_854),
.A2(n_887),
.B(n_800),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_887),
.B(n_860),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_904),
.A2(n_906),
.B(n_907),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_795),
.B(n_808),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_899),
.A2(n_948),
.B(n_840),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_847),
.B(n_840),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_899),
.A2(n_948),
.B(n_887),
.C(n_878),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_946),
.A2(n_902),
.B(n_934),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_797),
.B(n_902),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_801),
.B(n_945),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_936),
.B(n_943),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_SL g1072 ( 
.A1(n_821),
.A2(n_833),
.B(n_834),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_969),
.B(n_793),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_SL g1076 ( 
.A1(n_919),
.A2(n_958),
.B(n_920),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_925),
.B(n_939),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_882),
.A2(n_916),
.B(n_809),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_811),
.A2(n_919),
.B(n_920),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_925),
.B(n_939),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_793),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_947),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_904),
.B(n_906),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_1087)
);

BUFx2_ASAP7_75t_SL g1088 ( 
.A(n_946),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_925),
.B(n_939),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_925),
.B(n_939),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_SL g1091 ( 
.A1(n_821),
.A2(n_833),
.B(n_834),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_936),
.B(n_466),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_936),
.B(n_466),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_974),
.A2(n_833),
.B(n_954),
.C(n_834),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_814),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_925),
.B(n_939),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_814),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_925),
.B(n_939),
.Y(n_1098)
);

CKINVDCx8_ASAP7_75t_R g1099 ( 
.A(n_942),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_824),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_811),
.A2(n_919),
.B(n_920),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_918),
.A2(n_472),
.B(n_927),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_925),
.B(n_939),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_829),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_811),
.A2(n_919),
.B(n_920),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_925),
.B(n_939),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_925),
.B(n_939),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_974),
.A2(n_833),
.B(n_954),
.C(n_834),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_814),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_813),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_904),
.B(n_906),
.Y(n_1117)
);

AOI21x1_ASAP7_75t_L g1118 ( 
.A1(n_882),
.A2(n_916),
.B(n_809),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_814),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_813),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_925),
.B(n_939),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_861),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_814),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_925),
.B(n_939),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_928),
.A2(n_831),
.B(n_804),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1075),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_1110),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_989),
.B(n_998),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_998),
.B(n_1078),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1016),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1078),
.B(n_1082),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1006),
.A2(n_992),
.B1(n_981),
.B2(n_1109),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1023),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_985),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1060),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_979),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_980),
.A2(n_1114),
.B(n_1094),
.C(n_1026),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1099),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1036),
.B(n_1033),
.Y(n_1139)
);

CKINVDCx8_ASAP7_75t_R g1140 ( 
.A(n_1088),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1007),
.A2(n_1008),
.B(n_1031),
.C(n_1103),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1084),
.B(n_1064),
.Y(n_1142)
);

INVx3_ASAP7_75t_SL g1143 ( 
.A(n_1029),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1082),
.A2(n_1112),
.B1(n_1113),
.B2(n_1109),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1001),
.A2(n_990),
.B(n_1076),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1017),
.B(n_984),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_987),
.B(n_1065),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1122),
.A2(n_1007),
.B(n_1071),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1116),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1120),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_988),
.A2(n_1022),
.B(n_1005),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1081),
.A2(n_1103),
.B(n_1111),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_987),
.B(n_1002),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_979),
.Y(n_1155)
);

CKINVDCx8_ASAP7_75t_R g1156 ( 
.A(n_993),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_984),
.B(n_1083),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1029),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1083),
.B(n_1014),
.Y(n_1159)
);

NOR2x1_ASAP7_75t_SL g1160 ( 
.A(n_987),
.B(n_1062),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1039),
.B(n_1069),
.Y(n_1161)
);

OR2x2_ASAP7_75t_SL g1162 ( 
.A(n_1066),
.B(n_1053),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1086),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1073),
.A2(n_1077),
.B(n_1074),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_1060),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1089),
.B(n_1112),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1089),
.A2(n_1113),
.B1(n_1098),
.B2(n_1124),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1080),
.A2(n_1102),
.B(n_1106),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1056),
.B(n_1097),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_986),
.B(n_1090),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1086),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_983),
.A2(n_1008),
.B1(n_1041),
.B2(n_1081),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1117),
.B(n_1068),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1107),
.A2(n_1108),
.B(n_994),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1096),
.B(n_1121),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1003),
.A2(n_1030),
.B(n_1038),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_1011),
.B(n_1044),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1012),
.A2(n_1021),
.B(n_1111),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1012),
.A2(n_1019),
.B(n_1024),
.Y(n_1179)
);

CKINVDCx8_ASAP7_75t_R g1180 ( 
.A(n_1100),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_996),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_983),
.B(n_1034),
.C(n_1024),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1025),
.A2(n_1010),
.B(n_1034),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1027),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1025),
.A2(n_1020),
.B(n_1009),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1042),
.B(n_1044),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_997),
.A2(n_1061),
.B(n_1049),
.C(n_1045),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1000),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_991),
.A2(n_1125),
.B(n_1085),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1117),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1045),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_997),
.B(n_1049),
.Y(n_1192)
);

O2A1O1Ixp5_ASAP7_75t_L g1193 ( 
.A1(n_1051),
.A2(n_1061),
.B(n_1037),
.C(n_1079),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1000),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1048),
.B(n_1040),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1056),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1000),
.Y(n_1198)
);

BUFx4_ASAP7_75t_SL g1199 ( 
.A(n_1054),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1040),
.B(n_1047),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_982),
.A2(n_1015),
.B1(n_1035),
.B2(n_1062),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1097),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_995),
.A2(n_999),
.B(n_982),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1115),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1115),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1070),
.B(n_1057),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_SL g1207 ( 
.A(n_1048),
.B(n_1119),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1052),
.B(n_1050),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1087),
.A2(n_1104),
.B(n_1101),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1040),
.B(n_1047),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1095),
.B(n_1123),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1050),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1095),
.B(n_1123),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1119),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1095),
.B(n_1123),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1067),
.Y(n_1216)
);

AO22x2_ASAP7_75t_L g1217 ( 
.A1(n_1004),
.A2(n_1018),
.B1(n_1043),
.B2(n_1046),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1047),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1052),
.B(n_1032),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1055),
.B(n_1118),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1063),
.A2(n_1028),
.B(n_1105),
.C(n_1072),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1091),
.B(n_1004),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1002),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1013),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1110),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1006),
.A2(n_939),
.B1(n_941),
.B2(n_925),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1002),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_989),
.B(n_925),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_987),
.B(n_1065),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_987),
.B(n_1065),
.Y(n_1230)
);

NAND2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1056),
.B(n_791),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1006),
.A2(n_939),
.B1(n_941),
.B2(n_925),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1001),
.A2(n_1005),
.B(n_990),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_980),
.A2(n_974),
.B(n_821),
.C(n_833),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1036),
.A2(n_810),
.B(n_797),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_983),
.A2(n_954),
.B1(n_974),
.B2(n_833),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_989),
.B(n_925),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1039),
.B(n_847),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1036),
.B(n_1033),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_L g1240 ( 
.A(n_1029),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1013),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_989),
.B(n_925),
.Y(n_1242)
);

OR2x2_ASAP7_75t_SL g1243 ( 
.A(n_1066),
.B(n_837),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1013),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_987),
.B(n_1065),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1002),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_987),
.B(n_1065),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1056),
.B(n_791),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1036),
.B(n_1033),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1075),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_987),
.B(n_1065),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1036),
.A2(n_954),
.B1(n_834),
.B2(n_833),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1075),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1060),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_987),
.B(n_1065),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_989),
.B(n_925),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1007),
.A2(n_954),
.B(n_919),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_989),
.B(n_925),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1200),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1236),
.A2(n_1235),
.B(n_1252),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1132),
.A2(n_1182),
.B1(n_1153),
.B2(n_1257),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1130),
.Y(n_1262)
);

CKINVDCx14_ASAP7_75t_R g1263 ( 
.A(n_1138),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1177),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1132),
.A2(n_1182),
.B1(n_1153),
.B2(n_1257),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1151),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1136),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1210),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1177),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1224),
.Y(n_1272)
);

INVx4_ASAP7_75t_SL g1273 ( 
.A(n_1216),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1186),
.A2(n_1172),
.B1(n_1149),
.B2(n_1226),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1147),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1166),
.B(n_1192),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1136),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

NAND2x1p5_ASAP7_75t_L g1279 ( 
.A(n_1147),
.B(n_1229),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1166),
.B(n_1144),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1226),
.A2(n_1232),
.B1(n_1177),
.B2(n_1195),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1136),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1196),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1240),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1232),
.A2(n_1126),
.B1(n_1253),
.B2(n_1250),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1184),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1240),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1209),
.A2(n_1203),
.B(n_1179),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1133),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1222),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1225),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_SL g1292 ( 
.A1(n_1160),
.A2(n_1187),
.B(n_1137),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1126),
.A2(n_1250),
.B1(n_1253),
.B2(n_1239),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1143),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1161),
.B(n_1249),
.Y(n_1295)
);

AO21x1_ASAP7_75t_SL g1296 ( 
.A1(n_1201),
.A2(n_1191),
.B(n_1128),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1229),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1139),
.A2(n_1142),
.B1(n_1167),
.B2(n_1159),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1167),
.A2(n_1170),
.B1(n_1175),
.B2(n_1256),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1144),
.B(n_1196),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1150),
.Y(n_1301)
);

NAND2x1p5_ASAP7_75t_L g1302 ( 
.A(n_1230),
.B(n_1245),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1228),
.A2(n_1258),
.B1(n_1242),
.B2(n_1256),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1228),
.A2(n_1258),
.B1(n_1242),
.B2(n_1237),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1237),
.A2(n_1255),
.B1(n_1230),
.B2(n_1245),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1238),
.A2(n_1207),
.B1(n_1255),
.B2(n_1251),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1241),
.Y(n_1307)
);

BUFx2_ASAP7_75t_SL g1308 ( 
.A(n_1140),
.Y(n_1308)
);

NAND2x1_ASAP7_75t_L g1309 ( 
.A(n_1148),
.B(n_1247),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1207),
.A2(n_1128),
.B1(n_1247),
.B2(n_1251),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1244),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1165),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1254),
.A2(n_1135),
.B1(n_1146),
.B2(n_1154),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1183),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1212),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1157),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1183),
.B(n_1173),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1127),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1145),
.A2(n_1209),
.B(n_1174),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1193),
.A2(n_1233),
.B(n_1152),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1234),
.B(n_1141),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1178),
.A2(n_1179),
.B1(n_1173),
.B2(n_1154),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1215),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1208),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1185),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1134),
.B(n_1190),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1199),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1198),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1178),
.A2(n_1176),
.B(n_1145),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1174),
.A2(n_1152),
.B(n_1203),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1231),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1198),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1189),
.A2(n_1168),
.B(n_1164),
.Y(n_1333)
);

INVx6_ASAP7_75t_L g1334 ( 
.A(n_1206),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1156),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1221),
.A2(n_1220),
.B(n_1219),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1163),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1217),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1211),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1162),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1243),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1211),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1206),
.A2(n_1180),
.B1(n_1246),
.B2(n_1190),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1223),
.A2(n_1246),
.B1(n_1227),
.B2(n_1171),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1223),
.B(n_1227),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1181),
.A2(n_1202),
.B1(n_1214),
.B2(n_1205),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1213),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1158),
.A2(n_1169),
.B1(n_1214),
.B2(n_1202),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1213),
.Y(n_1349)
);

AO21x1_ASAP7_75t_L g1350 ( 
.A1(n_1248),
.A2(n_1169),
.B(n_1213),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1155),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1197),
.A2(n_1204),
.B1(n_1205),
.B2(n_1194),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1248),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1188),
.A2(n_1209),
.B(n_1189),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1188),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_SL g1356 ( 
.A(n_1188),
.B(n_1194),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1194),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1225),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1225),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1236),
.A2(n_954),
.B(n_619),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1132),
.A2(n_954),
.B1(n_974),
.B2(n_833),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1218),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1129),
.B(n_1131),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1128),
.B(n_1036),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1252),
.A2(n_735),
.B1(n_833),
.B2(n_834),
.Y(n_1366)
);

AO21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1172),
.A2(n_1008),
.B(n_992),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1225),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1329),
.A2(n_1338),
.B(n_1288),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1314),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1283),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1283),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1329),
.A2(n_1338),
.B(n_1333),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1309),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1269),
.B(n_1276),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1269),
.B(n_1259),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1314),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1363),
.Y(n_1378)
);

NAND2xp33_ASAP7_75t_R g1379 ( 
.A(n_1335),
.B(n_1264),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1324),
.B(n_1290),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1317),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1358),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1291),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1276),
.B(n_1300),
.Y(n_1384)
);

INVxp33_ASAP7_75t_SL g1385 ( 
.A(n_1335),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1325),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1290),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1354),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1300),
.B(n_1280),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1334),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1362),
.A2(n_1366),
.B(n_1361),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1319),
.A2(n_1330),
.B(n_1292),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1309),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1395)
);

CKINVDCx6p67_ASAP7_75t_R g1396 ( 
.A(n_1286),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1397)
);

OAI21xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1280),
.A2(n_1265),
.B(n_1261),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1286),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1360),
.B(n_1364),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1281),
.B(n_1367),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1321),
.B(n_1336),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1367),
.B(n_1301),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1350),
.A2(n_1341),
.B(n_1320),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1292),
.A2(n_1322),
.B(n_1260),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1330),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1330),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1340),
.A2(n_1274),
.B1(n_1310),
.B2(n_1305),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1368),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1303),
.B(n_1304),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1319),
.A2(n_1336),
.B(n_1340),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1336),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1365),
.B(n_1299),
.Y(n_1413)
);

AOI21xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1287),
.A2(n_1306),
.B(n_1295),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1298),
.A2(n_1316),
.B(n_1285),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1289),
.A2(n_1307),
.B(n_1311),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1312),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1293),
.B(n_1318),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1270),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1345),
.A2(n_1331),
.B(n_1343),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1275),
.B(n_1297),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1328),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1332),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1262),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1266),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1296),
.B(n_1302),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1272),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1402),
.B(n_1297),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1370),
.B(n_1302),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1370),
.B(n_1302),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1389),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1402),
.B(n_1279),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1411),
.B(n_1349),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1377),
.B(n_1315),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1386),
.B(n_1337),
.Y(n_1435)
);

AO31x2_ASAP7_75t_L g1436 ( 
.A1(n_1378),
.A2(n_1353),
.A3(n_1342),
.B(n_1347),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1412),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1411),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1376),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1411),
.B(n_1369),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1376),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1390),
.B(n_1337),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1390),
.B(n_1273),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1373),
.B(n_1273),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1398),
.B(n_1353),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1373),
.B(n_1406),
.Y(n_1446)
);

OAI221xp5_ASAP7_75t_L g1447 ( 
.A1(n_1392),
.A2(n_1313),
.B1(n_1344),
.B2(n_1359),
.C(n_1346),
.Y(n_1447)
);

OAI321xp33_ASAP7_75t_L g1448 ( 
.A1(n_1410),
.A2(n_1348),
.A3(n_1326),
.B1(n_1352),
.B2(n_1287),
.C(n_1323),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1381),
.B(n_1273),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1373),
.B(n_1406),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1373),
.B(n_1273),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1407),
.B(n_1339),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1393),
.B(n_1351),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1447),
.A2(n_1408),
.B(n_1401),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1439),
.B(n_1383),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1447),
.A2(n_1413),
.B1(n_1414),
.B2(n_1418),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1441),
.B(n_1400),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1441),
.B(n_1400),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1447),
.A2(n_1415),
.B1(n_1398),
.B2(n_1414),
.C(n_1420),
.Y(n_1460)
);

AOI211xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1448),
.A2(n_1444),
.B(n_1451),
.C(n_1445),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1442),
.B(n_1422),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1442),
.B(n_1423),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1442),
.B(n_1384),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1448),
.B(n_1417),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1445),
.B(n_1405),
.C(n_1401),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1428),
.B(n_1384),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1428),
.B(n_1387),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1429),
.B(n_1375),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1445),
.B(n_1395),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1448),
.A2(n_1405),
.B(n_1379),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1443),
.A2(n_1396),
.B1(n_1419),
.B2(n_1405),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1443),
.A2(n_1426),
.B(n_1403),
.Y(n_1473)
);

NAND4xp25_ASAP7_75t_SL g1474 ( 
.A(n_1443),
.B(n_1327),
.C(n_1419),
.D(n_1426),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1449),
.B(n_1374),
.Y(n_1475)
);

NAND3xp33_ASAP7_75t_L g1476 ( 
.A(n_1433),
.B(n_1405),
.C(n_1380),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1434),
.B(n_1397),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1449),
.B(n_1374),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1429),
.B(n_1375),
.Y(n_1479)
);

NOR3xp33_ASAP7_75t_L g1480 ( 
.A(n_1444),
.B(n_1284),
.C(n_1404),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1380),
.C(n_1427),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1429),
.B(n_1404),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1449),
.B(n_1374),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1430),
.B(n_1412),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1434),
.B(n_1371),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1430),
.B(n_1412),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1434),
.B(n_1372),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1434),
.B(n_1403),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1449),
.B(n_1374),
.Y(n_1489)
);

OAI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1433),
.A2(n_1382),
.B1(n_1284),
.B2(n_1308),
.C(n_1391),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1435),
.B(n_1416),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1430),
.B(n_1393),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1431),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1449),
.B(n_1374),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1435),
.B(n_1416),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1443),
.A2(n_1374),
.B(n_1394),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1433),
.B(n_1427),
.C(n_1424),
.Y(n_1497)
);

OAI21xp33_ASAP7_75t_L g1498 ( 
.A1(n_1432),
.A2(n_1440),
.B(n_1438),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1435),
.B(n_1416),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_L g1500 ( 
.A(n_1440),
.B(n_1424),
.C(n_1425),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1430),
.B(n_1393),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1449),
.A2(n_1385),
.B(n_1394),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1470),
.B(n_1453),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1491),
.B(n_1453),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1482),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1492),
.B(n_1446),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1460),
.B(n_1456),
.C(n_1465),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1495),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1499),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1482),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1471),
.B(n_1449),
.Y(n_1512)
);

OR2x6_ASAP7_75t_SL g1513 ( 
.A(n_1466),
.B(n_1476),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1453),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1497),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1497),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1501),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1501),
.B(n_1446),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1454),
.A2(n_1425),
.B1(n_1438),
.B2(n_1388),
.C(n_1308),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1500),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1469),
.B(n_1450),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1500),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1493),
.B(n_1484),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1486),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1458),
.B(n_1452),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_1450),
.Y(n_1527)
);

NAND2x1_ASAP7_75t_L g1528 ( 
.A(n_1481),
.B(n_1444),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1481),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1485),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1464),
.B(n_1453),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1487),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1455),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1488),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1457),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1459),
.B(n_1452),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1466),
.B(n_1437),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1480),
.B(n_1437),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1476),
.B(n_1440),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1498),
.B(n_1440),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1524),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1535),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1508),
.B(n_1396),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1535),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1510),
.B(n_1462),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1515),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_1444),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1538),
.B(n_1475),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1533),
.B(n_1463),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1519),
.B(n_1451),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1519),
.B(n_1451),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1510),
.B(n_1467),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1522),
.B(n_1451),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1503),
.B(n_1477),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1516),
.Y(n_1557)
);

NOR3xp33_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1490),
.C(n_1454),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1522),
.B(n_1478),
.Y(n_1559)
);

NAND4xp75_ASAP7_75t_L g1560 ( 
.A(n_1520),
.B(n_1483),
.C(n_1494),
.D(n_1489),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1522),
.B(n_1496),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1534),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1520),
.B(n_1472),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_L g1564 ( 
.A(n_1529),
.B(n_1461),
.C(n_1498),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1527),
.B(n_1473),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1512),
.A2(n_1474),
.B1(n_1502),
.B2(n_1421),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1526),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1538),
.B(n_1524),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1526),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1502),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1536),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1503),
.B(n_1505),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1436),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1524),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1505),
.B(n_1436),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1521),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1436),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1562),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1543),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1548),
.B(n_1529),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1571),
.B(n_1399),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1563),
.A2(n_1558),
.B(n_1564),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1551),
.B(n_1534),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1547),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1569),
.B(n_1549),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1538),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1577),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1550),
.B(n_1531),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1577),
.B(n_1568),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1537),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1542),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1544),
.B(n_1531),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1560),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1531),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1572),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1567),
.A2(n_1549),
.B1(n_1528),
.B2(n_1569),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1554),
.B(n_1532),
.Y(n_1605)
);

NAND2x1_ASAP7_75t_L g1606 ( 
.A(n_1549),
.B(n_1537),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1576),
.A2(n_1528),
.B(n_1513),
.C(n_1523),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1569),
.B(n_1537),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1554),
.B(n_1532),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1547),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1545),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1545),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1514),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1556),
.B(n_1514),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1559),
.B(n_1552),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1559),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1552),
.B(n_1509),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1574),
.B(n_1513),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1553),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1553),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1565),
.B(n_1521),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1592),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1523),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1603),
.A2(n_1600),
.B1(n_1580),
.B2(n_1604),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1621),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_L g1626 ( 
.A(n_1607),
.B(n_1565),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1615),
.B(n_1565),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1618),
.A2(n_1539),
.B1(n_1540),
.B2(n_1513),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1579),
.B(n_1509),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1578),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1583),
.B(n_1263),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1592),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1582),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1581),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1591),
.B(n_1575),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1584),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1591),
.B(n_1608),
.Y(n_1638)
);

INVx2_ASAP7_75t_SL g1639 ( 
.A(n_1621),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1588),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1621),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1575),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1594),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1597),
.B(n_1575),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1596),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1581),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1596),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1616),
.A2(n_1539),
.B1(n_1541),
.B2(n_1540),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1598),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1602),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1611),
.B(n_1294),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1612),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1587),
.Y(n_1653)
);

AO21x2_ASAP7_75t_L g1654 ( 
.A1(n_1607),
.A2(n_1539),
.B(n_1540),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1585),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1606),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1573),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1622),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1593),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1655),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1628),
.A2(n_1606),
.B1(n_1593),
.B2(n_1597),
.C(n_1589),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1638),
.B(n_1585),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1623),
.A2(n_1628),
.B(n_1626),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1655),
.B(n_1589),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1630),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1624),
.A2(n_1609),
.B(n_1599),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_1619),
.Y(n_1667)
);

OAI31xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1626),
.A2(n_1617),
.A3(n_1590),
.B(n_1610),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1653),
.A2(n_1614),
.B(n_1613),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1649),
.A2(n_1595),
.B(n_1601),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1617),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1656),
.A2(n_1610),
.B1(n_1590),
.B2(n_1620),
.Y(n_1672)
);

AOI32xp33_ASAP7_75t_L g1673 ( 
.A1(n_1630),
.A2(n_1541),
.A3(n_1555),
.B1(n_1576),
.B2(n_1573),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1638),
.B(n_1555),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1651),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1656),
.A2(n_1506),
.B1(n_1511),
.B2(n_1525),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1630),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1645),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1622),
.Y(n_1679)
);

AOI321xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1635),
.A2(n_1438),
.A3(n_1518),
.B1(n_1507),
.B2(n_1504),
.C(n_1506),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1634),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1656),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1663),
.B(n_1652),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1660),
.B(n_1652),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1662),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1675),
.B(n_1632),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1662),
.B(n_1636),
.Y(n_1687)
);

NAND2x1_ASAP7_75t_L g1688 ( 
.A(n_1682),
.B(n_1639),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1665),
.B(n_1649),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1682),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1682),
.Y(n_1691)
);

AOI222xp33_ASAP7_75t_L g1692 ( 
.A1(n_1661),
.A2(n_1650),
.B1(n_1648),
.B2(n_1646),
.C1(n_1635),
.C2(n_1645),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1671),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1658),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1664),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1681),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1677),
.B(n_1650),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1677),
.B(n_1646),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1681),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1671),
.B(n_1636),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1683),
.A2(n_1668),
.B(n_1659),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1696),
.A2(n_1678),
.B1(n_1666),
.B2(n_1654),
.C(n_1679),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1685),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_L g1705 ( 
.A(n_1686),
.B(n_1667),
.C(n_1672),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1692),
.A2(n_1654),
.B1(n_1636),
.B2(n_1674),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1687),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1700),
.Y(n_1708)
);

OAI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1700),
.A2(n_1689),
.B(n_1690),
.C(n_1684),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1697),
.A2(n_1654),
.B1(n_1694),
.B2(n_1699),
.C(n_1693),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1701),
.A2(n_1654),
.B1(n_1670),
.B2(n_1669),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1693),
.B(n_1674),
.Y(n_1712)
);

AOI211x1_ASAP7_75t_L g1713 ( 
.A1(n_1702),
.A2(n_1698),
.B(n_1701),
.C(n_1687),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1705),
.B(n_1695),
.C(n_1691),
.D(n_1673),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1708),
.B(n_1691),
.Y(n_1715)
);

NAND4xp25_ASAP7_75t_L g1716 ( 
.A(n_1706),
.B(n_1695),
.C(n_1647),
.D(n_1641),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1712),
.Y(n_1717)
);

OAI322xp33_ASAP7_75t_L g1718 ( 
.A1(n_1704),
.A2(n_1688),
.A3(n_1633),
.B1(n_1639),
.B2(n_1647),
.C1(n_1625),
.C2(n_1641),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1711),
.B(n_1639),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1709),
.B(n_1688),
.Y(n_1720)
);

NOR4xp75_ASAP7_75t_L g1721 ( 
.A(n_1707),
.B(n_1629),
.C(n_1631),
.D(n_1642),
.Y(n_1721)
);

NAND5xp2_ASAP7_75t_L g1722 ( 
.A(n_1703),
.B(n_1710),
.C(n_1680),
.D(n_1644),
.E(n_1642),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1716),
.A2(n_1633),
.B1(n_1641),
.B2(n_1625),
.C(n_1647),
.Y(n_1723)
);

NOR3x1_ASAP7_75t_L g1724 ( 
.A(n_1714),
.B(n_1719),
.C(n_1717),
.Y(n_1724)
);

NOR4xp25_ASAP7_75t_L g1725 ( 
.A(n_1718),
.B(n_1625),
.C(n_1640),
.D(n_1637),
.Y(n_1725)
);

NAND4xp75_ASAP7_75t_L g1726 ( 
.A(n_1720),
.B(n_1644),
.C(n_1642),
.D(n_1643),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_L g1727 ( 
.A(n_1713),
.B(n_1634),
.C(n_1637),
.Y(n_1727)
);

NAND4xp25_ASAP7_75t_L g1728 ( 
.A(n_1715),
.B(n_1294),
.C(n_1284),
.D(n_1629),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1722),
.A2(n_1643),
.B(n_1640),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1727),
.Y(n_1730)
);

INVxp67_ASAP7_75t_SL g1731 ( 
.A(n_1724),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1726),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1728),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1729),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1725),
.B(n_1721),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1732),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1732),
.Y(n_1737)
);

AOI21xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1735),
.A2(n_1723),
.B(n_1657),
.Y(n_1738)
);

NOR4xp25_ASAP7_75t_L g1739 ( 
.A(n_1731),
.B(n_1734),
.C(n_1735),
.D(n_1733),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1730),
.B(n_1644),
.Y(n_1740)
);

XNOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1739),
.B(n_1730),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1740),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1737),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1741),
.A2(n_1739),
.B(n_1736),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1744),
.B(n_1742),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1742),
.B1(n_1743),
.B2(n_1738),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1745),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1743),
.B1(n_1631),
.B2(n_1657),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_SL g1749 ( 
.A1(n_1746),
.A2(n_1676),
.B(n_1356),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1748),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1749),
.A2(n_1627),
.B(n_1277),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1750),
.A2(n_1627),
.B1(n_1355),
.B2(n_1511),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1751),
.B1(n_1627),
.B2(n_1355),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_R g1754 ( 
.A1(n_1753),
.A2(n_1282),
.B1(n_1268),
.B2(n_1357),
.C(n_1356),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1278),
.B(n_1277),
.C(n_1357),
.Y(n_1755)
);


endmodule