module fake_jpeg_12652_n_601 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_601);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_62),
.B(n_69),
.Y(n_168)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_18),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_70),
.B(n_72),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_75),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_76),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_77),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_31),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_78),
.B(n_79),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_31),
.B(n_16),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_80),
.B(n_82),
.Y(n_173)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_83),
.Y(n_157)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_84),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_85),
.B(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_86),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_32),
.B(n_16),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_88),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_89),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_15),
.C(n_11),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_90),
.B(n_91),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_34),
.B(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_92),
.B(n_96),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_11),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_40),
.B(n_11),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_104),
.B(n_55),
.Y(n_200)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_37),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_117),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_37),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_40),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_125),
.Y(n_189)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_33),
.Y(n_125)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_27),
.B(n_44),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_133),
.B(n_113),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_137),
.A2(n_138),
.B1(n_159),
.B2(n_98),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_74),
.A2(n_52),
.B1(n_50),
.B2(n_21),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g279 ( 
.A(n_144),
.Y(n_279)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_48),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_147),
.B(n_153),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_46),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_149),
.B(n_93),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_100),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_84),
.A2(n_21),
.B1(n_46),
.B2(n_33),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_161),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_167),
.B(n_180),
.Y(n_249)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_90),
.B(n_46),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_171),
.A2(n_200),
.B(n_64),
.Y(n_224)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_89),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_89),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_182),
.B(n_188),
.Y(n_256)
);

HAxp5_ASAP7_75t_SL g184 ( 
.A(n_89),
.B(n_44),
.CON(n_184),
.SN(n_184)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_64),
.Y(n_240)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_113),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_121),
.A2(n_25),
.B1(n_27),
.B2(n_39),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_190),
.A2(n_75),
.B1(n_68),
.B2(n_59),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_103),
.A2(n_33),
.B1(n_25),
.B2(n_39),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_41),
.B1(n_36),
.B2(n_194),
.Y(n_215)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_195),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_115),
.B(n_55),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_197),
.B(n_131),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_110),
.B(n_51),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_105),
.Y(n_235)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_88),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_113),
.C(n_64),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_212),
.B(n_250),
.C(n_160),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_214),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_215),
.A2(n_239),
.B1(n_243),
.B2(n_157),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_149),
.A2(n_111),
.B1(n_108),
.B2(n_71),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_216),
.A2(n_226),
.B1(n_230),
.B2(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_219),
.B(n_220),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_221),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_222),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_61),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_223),
.B(n_229),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_224),
.B(n_238),
.Y(n_304)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g313 ( 
.A(n_228),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_41),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_66),
.B1(n_76),
.B2(n_73),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_36),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_234),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_173),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_235),
.B(n_237),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_173),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_190),
.A2(n_65),
.B1(n_94),
.B2(n_119),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_171),
.B(n_0),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_253),
.Y(n_295)
);

INVx3_ASAP7_75t_SL g242 ( 
.A(n_158),
.Y(n_242)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_124),
.B1(n_97),
.B2(n_114),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_132),
.Y(n_244)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_244),
.Y(n_315)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_246),
.Y(n_337)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_139),
.B(n_123),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_134),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_83),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

BUFx2_ASAP7_75t_SL g252 ( 
.A(n_181),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_252),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_10),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_137),
.A2(n_107),
.B1(n_99),
.B2(n_10),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_159),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_255),
.A2(n_134),
.B1(n_166),
.B2(n_204),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_189),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_260),
.Y(n_301)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_193),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_4),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_264),
.Y(n_318)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_146),
.Y(n_263)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_168),
.B(n_4),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_168),
.B(n_5),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_268),
.Y(n_326)
);

CKINVDCx12_ASAP7_75t_R g267 ( 
.A(n_150),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_267),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_164),
.B(n_5),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_193),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_275),
.Y(n_335)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_150),
.Y(n_271)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

CKINVDCx12_ASAP7_75t_R g272 ( 
.A(n_144),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_272),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_205),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_273),
.A2(n_274),
.B1(n_282),
.B2(n_210),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_148),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_187),
.B(n_9),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_172),
.B(n_156),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_278),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_133),
.A2(n_128),
.B1(n_145),
.B2(n_196),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_138),
.B1(n_235),
.B2(n_212),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_172),
.B(n_136),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_280),
.B(n_284),
.Y(n_303)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_192),
.Y(n_281)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_162),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_169),
.B(n_142),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_249),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_287),
.B(n_316),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_288),
.A2(n_282),
.B1(n_258),
.B2(n_263),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_219),
.A2(n_154),
.B(n_183),
.C(n_157),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_291),
.B(n_320),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_198),
.B(n_141),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_296),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_203),
.B1(n_140),
.B2(n_135),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_298),
.A2(n_311),
.B1(n_321),
.B2(n_339),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_219),
.A2(n_148),
.B(n_199),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_300),
.B(n_305),
.Y(n_370)
);

AND2x2_ASAP7_75t_SL g307 ( 
.A(n_241),
.B(n_129),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_325),
.C(n_329),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_310),
.A2(n_324),
.B1(n_242),
.B2(n_225),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_206),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_152),
.B1(n_196),
.B2(n_163),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_250),
.A2(n_238),
.B1(n_248),
.B2(n_268),
.Y(n_321)
);

AOI22x1_ASAP7_75t_L g324 ( 
.A1(n_250),
.A2(n_238),
.B1(n_231),
.B2(n_275),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_283),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_232),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_248),
.B(n_186),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_213),
.B(n_209),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_331),
.B(n_333),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_215),
.B(n_162),
.Y(n_332)
);

INVx4_ASAP7_75t_SL g378 ( 
.A(n_332),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_245),
.B(n_132),
.Y(n_333)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_238),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_341),
.B(n_345),
.Y(n_387)
);

BUFx24_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_342),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_343),
.A2(n_380),
.B(n_382),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_270),
.B1(n_213),
.B2(n_217),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_346),
.Y(n_394)
);

CKINVDCx10_ASAP7_75t_R g347 ( 
.A(n_290),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_347),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_350),
.Y(n_412)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_293),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_279),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_351),
.B(n_352),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_279),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_299),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_361),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_286),
.B(n_279),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_355),
.B(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_293),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

BUFx12_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_357),
.Y(n_390)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_358),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_359),
.A2(n_236),
.B1(n_221),
.B2(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_363),
.Y(n_391)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_366),
.Y(n_415)
);

INVx8_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_289),
.A2(n_179),
.B1(n_217),
.B2(n_265),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_383),
.B1(n_374),
.B2(n_370),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_372),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_288),
.A2(n_265),
.B1(n_218),
.B2(n_261),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_313),
.B1(n_332),
.B2(n_261),
.Y(n_389)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_377),
.Y(n_405)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_294),
.B(n_218),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_331),
.B(n_227),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_214),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_303),
.B(n_227),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_379),
.A2(n_337),
.B1(n_338),
.B2(n_309),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_271),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_232),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_289),
.A2(n_321),
.B1(n_324),
.B2(n_296),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_360),
.A2(n_304),
.B(n_285),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_304),
.B(n_311),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_416),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_360),
.A2(n_300),
.B(n_325),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_389),
.A2(n_399),
.B1(n_409),
.B2(n_413),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_393),
.A2(n_398),
.B1(n_407),
.B2(n_410),
.Y(n_446)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_364),
.A2(n_329),
.B(n_310),
.Y(n_396)
);

AO21x1_ASAP7_75t_L g449 ( 
.A1(n_396),
.A2(n_380),
.B(n_347),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_343),
.A2(n_291),
.B(n_310),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_307),
.B1(n_320),
.B2(n_326),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_359),
.A2(n_320),
.B1(n_313),
.B2(n_251),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_307),
.C(n_295),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_419),
.C(n_369),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_320),
.B1(n_323),
.B2(n_228),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_370),
.A2(n_330),
.B1(n_302),
.B2(n_179),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_378),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_368),
.A2(n_247),
.B1(n_340),
.B2(n_246),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_345),
.A2(n_340),
.B1(n_337),
.B2(n_315),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_376),
.B(n_312),
.C(n_214),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_381),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_426),
.C(n_432),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_404),
.B(n_354),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_421),
.B(n_424),
.Y(n_462)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_377),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_422),
.B(n_429),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_404),
.B(n_373),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_375),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_391),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_433),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_353),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_391),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_342),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_435),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_401),
.B(n_342),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_406),
.B(n_378),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_442),
.Y(n_458)
);

INVx13_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_384),
.B(n_341),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_386),
.Y(n_442)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_344),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_452),
.Y(n_473)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_372),
.C(n_365),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_388),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_350),
.Y(n_451)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_408),
.B(n_363),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_396),
.B(n_405),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_454),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_432),
.C(n_450),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_431),
.A2(n_397),
.B(n_387),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_464),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_451),
.Y(n_464)
);

BUFx24_ASAP7_75t_SL g467 ( 
.A(n_435),
.Y(n_467)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_467),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_446),
.A2(n_385),
.B1(n_399),
.B2(n_394),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_468),
.A2(n_481),
.B1(n_427),
.B2(n_436),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_405),
.Y(n_470)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_470),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_412),
.Y(n_471)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_423),
.A2(n_394),
.B1(n_385),
.B2(n_393),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_472),
.A2(n_476),
.B1(n_407),
.B2(n_436),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_439),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_430),
.Y(n_478)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_412),
.Y(n_479)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_480),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_427),
.A2(n_385),
.B1(n_389),
.B2(n_409),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_437),
.C(n_424),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_483),
.B(n_487),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_420),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_493),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_496),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_488),
.C(n_504),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_482),
.A2(n_387),
.B(n_438),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_426),
.C(n_438),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_440),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_443),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_506),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_495),
.A2(n_502),
.B1(n_475),
.B2(n_464),
.Y(n_515)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_453),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_482),
.A2(n_422),
.B(n_449),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_473),
.Y(n_527)
);

XNOR2x1_ASAP7_75t_L g500 ( 
.A(n_456),
.B(n_411),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_500),
.B(n_474),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_461),
.A2(n_441),
.B1(n_425),
.B2(n_414),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_501),
.A2(n_481),
.B1(n_468),
.B2(n_465),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_472),
.A2(n_396),
.B1(n_398),
.B2(n_425),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_458),
.A2(n_410),
.B1(n_414),
.B2(n_416),
.Y(n_503)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_503),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_411),
.C(n_408),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_454),
.B(n_392),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_402),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_500),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_459),
.B(n_362),
.C(n_444),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_469),
.C(n_463),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_471),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_513),
.B(n_525),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_515),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_496),
.B(n_462),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_516),
.B(n_527),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_475),
.B1(n_478),
.B2(n_459),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_523),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_519),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_521),
.A2(n_502),
.B1(n_499),
.B2(n_489),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_490),
.A2(n_455),
.B(n_470),
.Y(n_523)
);

INVx11_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_479),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_526),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_486),
.B(n_480),
.C(n_474),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_488),
.C(n_506),
.Y(n_532)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_505),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_529),
.B(n_530),
.Y(n_542)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_507),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_532),
.B(n_541),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_517),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_537),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_504),
.C(n_491),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_538),
.A2(n_515),
.B1(n_510),
.B2(n_522),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_501),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_512),
.B(n_491),
.C(n_494),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_547),
.C(n_511),
.Y(n_560)
);

INVx13_ASAP7_75t_L g545 ( 
.A(n_524),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_545),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_514),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_465),
.C(n_461),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_513),
.C(n_511),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_554),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_540),
.A2(n_523),
.B(n_520),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_557),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_556),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_514),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_537),
.A2(n_518),
.B(n_522),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_539),
.B(n_509),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_558),
.B(n_559),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_540),
.A2(n_469),
.B1(n_463),
.B2(n_403),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_561),
.C(n_562),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_532),
.B(n_519),
.C(n_531),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_534),
.B(n_413),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_541),
.B(n_395),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_563),
.B(n_533),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_551),
.Y(n_566)
);

INVxp33_ASAP7_75t_SL g579 ( 
.A(n_566),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_547),
.C(n_544),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_567),
.B(n_571),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_574),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_549),
.A2(n_542),
.B1(n_548),
.B2(n_545),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_550),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_572),
.A2(n_379),
.B(n_356),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_552),
.A2(n_546),
.B1(n_403),
.B2(n_543),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_562),
.C(n_553),
.Y(n_575)
);

INVxp33_ASAP7_75t_L g582 ( 
.A(n_575),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_573),
.A2(n_567),
.B(n_564),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_578),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_573),
.A2(n_563),
.B1(n_417),
.B2(n_349),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_580),
.B(n_581),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_569),
.B(n_366),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_575),
.B(n_361),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_583),
.B(n_568),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_586),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_578),
.A2(n_565),
.B(n_568),
.Y(n_586)
);

AOI322xp5_ASAP7_75t_L g587 ( 
.A1(n_584),
.A2(n_371),
.A3(n_357),
.B1(n_358),
.B2(n_214),
.C1(n_281),
.C2(n_269),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_587),
.B(n_271),
.C(n_290),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_582),
.B(n_222),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_579),
.B(n_357),
.Y(n_591)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_591),
.Y(n_595)
);

AOI21x1_ASAP7_75t_L g593 ( 
.A1(n_588),
.A2(n_579),
.B(n_576),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_593),
.B(n_594),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_596),
.B(n_592),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_597),
.A2(n_595),
.B(n_589),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_598),
.B(n_586),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_259),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_244),
.B1(n_259),
.B2(n_210),
.Y(n_601)
);


endmodule