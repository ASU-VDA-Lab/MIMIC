module fake_jpeg_1624_n_670 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_670);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_670;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_9),
.Y(n_44)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_71),
.Y(n_145)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_75),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_76),
.B(n_79),
.Y(n_147)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_11),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_83),
.Y(n_222)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_11),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_92),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_28),
.B(n_8),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_94),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_25),
.B(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_95),
.B(n_104),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_12),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_106),
.B(n_14),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_113),
.Y(n_221)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_23),
.Y(n_120)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_127),
.Y(n_206)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_25),
.B(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_30),
.B(n_7),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_129),
.B(n_51),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_29),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_30),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_133),
.B(n_214),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_101),
.B1(n_130),
.B2(n_64),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_137),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_58),
.B1(n_60),
.B2(n_34),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_144),
.A2(n_151),
.B1(n_163),
.B2(n_167),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_38),
.B1(n_53),
.B2(n_60),
.Y(n_150)
);

OA22x2_ASAP7_75t_SL g238 ( 
.A1(n_150),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_53),
.B1(n_34),
.B2(n_59),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_71),
.B(n_46),
.C(n_57),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_161),
.B(n_200),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_58),
.B1(n_59),
.B2(n_48),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_67),
.A2(n_58),
.B1(n_59),
.B2(n_48),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_73),
.B(n_58),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_179),
.Y(n_274)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_68),
.A2(n_42),
.B1(n_24),
.B2(n_57),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_194),
.A2(n_196),
.B1(n_217),
.B2(n_218),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_87),
.A2(n_83),
.B1(n_63),
.B2(n_123),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_43),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_17),
.Y(n_232)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_65),
.Y(n_207)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_19),
.Y(n_241)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_66),
.Y(n_213)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_72),
.B(n_42),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_69),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_215),
.B(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_80),
.Y(n_216)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_123),
.A2(n_51),
.B1(n_43),
.B2(n_13),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_70),
.A2(n_43),
.B1(n_13),
.B2(n_14),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_75),
.A2(n_43),
.B1(n_13),
.B2(n_14),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_219),
.A2(n_163),
.B1(n_144),
.B2(n_194),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_137),
.A2(n_100),
.B1(n_88),
.B2(n_91),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g361 ( 
.A1(n_225),
.A2(n_238),
.B1(n_256),
.B2(n_275),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_229),
.Y(n_349)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_181),
.Y(n_230)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_232),
.B(n_281),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_124),
.B1(n_122),
.B2(n_94),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_233),
.A2(n_234),
.B1(n_243),
.B2(n_247),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_107),
.B1(n_81),
.B2(n_113),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_153),
.Y(n_235)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_237),
.Y(n_356)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_L g360 ( 
.A1(n_240),
.A2(n_273),
.B1(n_253),
.B2(n_302),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_241),
.B(n_244),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_156),
.B(n_19),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_242),
.B(n_251),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_206),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_156),
.B(n_17),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_245),
.Y(n_357)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_140),
.Y(n_246)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_246),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_148),
.A2(n_16),
.B1(n_7),
.B2(n_3),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_149),
.Y(n_248)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_249),
.Y(n_353)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_147),
.B(n_16),
.Y(n_251)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_141),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_138),
.Y(n_255)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_150),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_150),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_257),
.A2(n_217),
.B1(n_196),
.B2(n_159),
.Y(n_315)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_162),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_263),
.Y(n_305)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_162),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_264),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_145),
.Y(n_265)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_265),
.Y(n_365)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_266),
.B(n_267),
.Y(n_329)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_145),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_147),
.A2(n_180),
.B(n_158),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_179),
.Y(n_308)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_270),
.B(n_271),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_272),
.B(n_277),
.Y(n_341)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_273),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_180),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_276),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_146),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_280),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_168),
.B(n_4),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_221),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_282),
.B(n_283),
.Y(n_345)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_284),
.B(n_285),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_165),
.B(n_4),
.Y(n_285)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_190),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_286),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_287),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_169),
.A2(n_197),
.B1(n_164),
.B2(n_167),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_289),
.A2(n_290),
.B1(n_293),
.B2(n_297),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_176),
.A2(n_6),
.B1(n_178),
.B2(n_224),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_189),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_292),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_192),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_160),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_174),
.B(n_6),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_294),
.B(n_303),
.Y(n_364)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_134),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_177),
.B(n_182),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_166),
.Y(n_313)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_358)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_135),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_159),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_136),
.B(n_139),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_235),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_313),
.B(n_319),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_315),
.A2(n_320),
.B1(n_360),
.B2(n_299),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_323),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_153),
.B(n_184),
.C(n_193),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_257),
.A2(n_175),
.B1(n_210),
.B2(n_220),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_175),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_220),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_327),
.Y(n_376)
);

AO21x2_ASAP7_75t_L g325 ( 
.A1(n_268),
.A2(n_162),
.B(n_166),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_325),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_210),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_333),
.C(n_338),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_170),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_238),
.A2(n_170),
.B1(n_172),
.B2(n_154),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_340),
.B1(n_286),
.B2(n_272),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_226),
.B(n_172),
.C(n_193),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_246),
.B(n_166),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_336),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_248),
.B(n_193),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_236),
.B(n_190),
.C(n_202),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_238),
.A2(n_202),
.B1(n_279),
.B2(n_240),
.Y(n_340)
);

AOI22x1_ASAP7_75t_SL g347 ( 
.A1(n_229),
.A2(n_250),
.B1(n_283),
.B2(n_270),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_347),
.A2(n_325),
.B1(n_358),
.B2(n_304),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_231),
.B(n_252),
.C(n_254),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_354),
.C(n_271),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_249),
.B(n_239),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_259),
.B(n_228),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_228),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_317),
.B(n_291),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_366),
.B(n_380),
.C(n_405),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_367),
.Y(n_421)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_370),
.B(n_374),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_371),
.B(n_311),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_315),
.A2(n_357),
.B1(n_348),
.B2(n_309),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_372),
.A2(n_395),
.B1(n_404),
.B2(n_306),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_323),
.A2(n_265),
.B(n_267),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_373),
.A2(n_378),
.B(n_413),
.Y(n_424)
);

AO22x2_ASAP7_75t_L g374 ( 
.A1(n_320),
.A2(n_245),
.B1(n_282),
.B2(n_284),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_319),
.A2(n_292),
.B(n_277),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_332),
.Y(n_379)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_308),
.B(n_364),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_382),
.B(n_384),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_391),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_345),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_325),
.A2(n_260),
.B1(n_261),
.B2(n_295),
.Y(n_385)
);

AO22x1_ASAP7_75t_SL g446 ( 
.A1(n_385),
.A2(n_387),
.B1(n_401),
.B2(n_408),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_394),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_325),
.A2(n_237),
.B1(n_230),
.B2(n_293),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_388),
.A2(n_393),
.B1(n_408),
.B2(n_407),
.Y(n_439)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_389),
.Y(n_453)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_392),
.B(n_350),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_324),
.A2(n_263),
.B1(n_264),
.B2(n_325),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_329),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_357),
.A2(n_348),
.B1(n_309),
.B2(n_356),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_363),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_397),
.B(n_409),
.Y(n_448)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_399),
.A2(n_307),
.B1(n_356),
.B2(n_312),
.Y(n_425)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_322),
.A2(n_361),
.B1(n_331),
.B2(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_402),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_326),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_412),
.Y(n_431)
);

BUFx8_ASAP7_75t_L g404 ( 
.A(n_305),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_310),
.C(n_337),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_352),
.C(n_333),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_355),
.C(n_334),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_338),
.B(n_361),
.Y(n_407)
);

XNOR2x2_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_361),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_336),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_343),
.B(n_328),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_410),
.B(n_411),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_314),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_313),
.A2(n_350),
.B(n_346),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_414),
.A2(n_419),
.B(n_425),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_388),
.A2(n_361),
.B1(n_360),
.B2(n_335),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_415),
.A2(n_439),
.B1(n_445),
.B2(n_451),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_423),
.B(n_432),
.C(n_442),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_396),
.A2(n_328),
.B(n_334),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g433 ( 
.A1(n_376),
.A2(n_347),
.A3(n_312),
.B1(n_355),
.B2(n_342),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_435),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_342),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_344),
.Y(n_437)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_383),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_440),
.B(n_444),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_380),
.B(n_344),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_378),
.A2(n_349),
.B(n_316),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_369),
.B(n_316),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_376),
.A2(n_332),
.B1(n_349),
.B2(n_321),
.Y(n_445)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_306),
.B(n_321),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_374),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_353),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_398),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_381),
.B(n_353),
.Y(n_450)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_407),
.A2(n_311),
.B1(n_393),
.B2(n_375),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_406),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_407),
.A2(n_368),
.B1(n_375),
.B2(n_381),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_454),
.A2(n_407),
.B1(n_368),
.B2(n_392),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_456),
.B(n_472),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_457),
.B(n_437),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_366),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_432),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_439),
.A2(n_407),
.B1(n_384),
.B2(n_401),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_462),
.A2(n_464),
.B1(n_466),
.B2(n_473),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_440),
.A2(n_413),
.B1(n_394),
.B2(n_367),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_418),
.A2(n_374),
.B1(n_387),
.B2(n_373),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_424),
.A2(n_404),
.B(n_385),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_470),
.A2(n_443),
.B(n_447),
.Y(n_510)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_417),
.Y(n_471)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_418),
.A2(n_374),
.B1(n_412),
.B2(n_390),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_405),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_423),
.C(n_452),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_386),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_475),
.B(n_478),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_441),
.Y(n_476)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_421),
.B(n_400),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_444),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_481),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_426),
.Y(n_480)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_480),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_428),
.A2(n_374),
.B1(n_402),
.B2(n_379),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_483),
.Y(n_502)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_434),
.Y(n_484)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_484),
.Y(n_507)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_485),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_421),
.B(n_404),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_486),
.B(n_422),
.Y(n_504)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_436),
.Y(n_488)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_404),
.C(n_389),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_414),
.Y(n_495)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_436),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_491),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_448),
.Y(n_491)
);

AND2x4_ASAP7_75t_SL g492 ( 
.A(n_459),
.B(n_424),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_SL g559 ( 
.A1(n_492),
.A2(n_498),
.B(n_510),
.C(n_438),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_494),
.B(n_511),
.C(n_512),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_460),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_456),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_497),
.B(n_506),
.Y(n_537)
);

OAI22x1_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_425),
.B1(n_414),
.B2(n_438),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_465),
.A2(n_431),
.B1(n_428),
.B2(n_420),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_503),
.A2(n_467),
.B1(n_473),
.B2(n_466),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_504),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_463),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_509),
.B(n_515),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_449),
.C(n_442),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_431),
.C(n_420),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_479),
.B(n_450),
.Y(n_514)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_514),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_435),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_463),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_517),
.B(n_519),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_458),
.A2(n_430),
.B(n_451),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_459),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_455),
.B(n_467),
.Y(n_523)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_523),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_461),
.B(n_416),
.C(n_446),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_525),
.C(n_518),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_474),
.B(n_416),
.C(n_446),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_472),
.B(n_433),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_527),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_464),
.B(n_446),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_505),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_529),
.A2(n_539),
.B1(n_544),
.B2(n_545),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_556),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_480),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_532),
.B(n_548),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_521),
.A2(n_499),
.B1(n_468),
.B2(n_516),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_534),
.A2(n_498),
.B1(n_526),
.B2(n_524),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_550),
.Y(n_562)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_505),
.Y(n_538)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_538),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_523),
.Y(n_539)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_499),
.Y(n_541)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_455),
.Y(n_543)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_514),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_492),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_546),
.B(n_477),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_512),
.B(n_471),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_492),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_549),
.B(n_552),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_521),
.A2(n_468),
.B1(n_462),
.B2(n_487),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_554),
.B1(n_557),
.B2(n_558),
.Y(n_563)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_500),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_494),
.B(n_489),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_553),
.B(n_555),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_518),
.B(n_489),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_511),
.B(n_470),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_527),
.A2(n_469),
.B1(n_487),
.B2(n_415),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_516),
.A2(n_481),
.B1(n_438),
.B2(n_458),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_559),
.B(n_557),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_528),
.A2(n_510),
.B(n_519),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_560),
.A2(n_575),
.B(n_582),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_508),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_561),
.B(n_417),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_564),
.A2(n_574),
.B1(n_580),
.B2(n_559),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_533),
.A2(n_501),
.B1(n_525),
.B2(n_513),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_567),
.B(n_530),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_497),
.C(n_556),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_568),
.B(n_576),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_571),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_495),
.B1(n_501),
.B2(n_506),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_549),
.A2(n_520),
.B(n_513),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_542),
.B(n_520),
.C(n_507),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_554),
.A2(n_502),
.B1(n_507),
.B2(n_484),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_577),
.A2(n_536),
.B1(n_531),
.B2(n_552),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_550),
.B(n_547),
.C(n_537),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_578),
.B(n_535),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_547),
.B(n_502),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_553),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_541),
.A2(n_447),
.B1(n_445),
.B2(n_483),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_558),
.A2(n_485),
.B(n_490),
.Y(n_582)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_583),
.Y(n_592)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_584),
.Y(n_594)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_598),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_589),
.B(n_596),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_576),
.B(n_562),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_590),
.B(n_600),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_562),
.B(n_537),
.C(n_555),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_593),
.Y(n_610)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_570),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_563),
.A2(n_536),
.B1(n_531),
.B2(n_543),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_597),
.A2(n_582),
.B1(n_573),
.B2(n_566),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_545),
.C(n_488),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_602),
.C(n_565),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_578),
.B(n_559),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_601),
.B(n_607),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_579),
.B(n_496),
.C(n_559),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_569),
.B(n_496),
.Y(n_603)
);

CKINVDCx14_ASAP7_75t_R g619 ( 
.A(n_603),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_569),
.B(n_453),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_604),
.B(n_566),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_584),
.A2(n_559),
.B(n_570),
.C(n_573),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_605),
.A2(n_575),
.B(n_572),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_447),
.Y(n_607)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_608),
.Y(n_628)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_611),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_621),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_594),
.A2(n_585),
.B1(n_564),
.B2(n_560),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_613),
.B(n_614),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_587),
.B(n_574),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_615),
.B(n_623),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_599),
.B(n_565),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_620),
.B(n_592),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_585),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_596),
.A2(n_577),
.B(n_571),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_622),
.A2(n_624),
.B(n_605),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_590),
.B(n_581),
.C(n_580),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_595),
.B(n_453),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_625),
.B(n_598),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_631),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_629),
.B(n_632),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_625),
.B(n_600),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_R g632 ( 
.A(n_618),
.B(n_594),
.C(n_611),
.Y(n_632)
);

INVxp33_ASAP7_75t_L g645 ( 
.A(n_633),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_610),
.B(n_592),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_635),
.B(n_636),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_614),
.B(n_609),
.C(n_623),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_616),
.B(n_586),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_638),
.B(n_640),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_609),
.B(n_591),
.C(n_595),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_639),
.B(n_622),
.C(n_588),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_617),
.B(n_597),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_630),
.A2(n_619),
.B1(n_621),
.B2(n_613),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_641),
.B(n_646),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_639),
.B(n_602),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_636),
.B(n_618),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_647),
.B(n_648),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_608),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_649),
.B(n_626),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_634),
.A2(n_624),
.B(n_589),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_651),
.A2(n_633),
.B(n_645),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_650),
.B(n_630),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_654),
.B(n_656),
.Y(n_663)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_655),
.Y(n_660)
);

MAJx2_ASAP7_75t_L g656 ( 
.A(n_642),
.B(n_637),
.C(n_628),
.Y(n_656)
);

INVxp33_ASAP7_75t_L g662 ( 
.A(n_657),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_643),
.A2(n_632),
.B(n_631),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_658),
.A2(n_659),
.B(n_653),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_649),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_646),
.C(n_644),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_661),
.A2(n_664),
.B1(n_607),
.B2(n_453),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_662),
.A2(n_645),
.B(n_644),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_665),
.B(n_666),
.Y(n_667)
);

BUFx24_ASAP7_75t_SL g668 ( 
.A(n_667),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_668),
.B(n_660),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_669),
.B(n_663),
.Y(n_670)
);


endmodule