module fake_jpeg_29512_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_49),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_50),
.Y(n_94)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_69),
.B1(n_63),
.B2(n_51),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_93),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_51),
.B1(n_48),
.B2(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_101),
.Y(n_111)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_48),
.B1(n_61),
.B2(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_57),
.B1(n_54),
.B2(n_53),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_19),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_2),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_45),
.B1(n_60),
.B2(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_1),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_20),
.A3(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_113),
.B(n_118),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_17),
.A3(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_109),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_4),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_16),
.C(n_30),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_105),
.C(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_7),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_9),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_10),
.Y(n_122)
);

NOR4xp25_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_15),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_133),
.C(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_135),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_142),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_114),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_145),
.B(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_134),
.B1(n_139),
.B2(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_140),
.B1(n_132),
.B2(n_125),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_106),
.B(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_138),
.Y(n_153)
);


endmodule