module real_aes_6964_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_756;
wire n_713;
wire n_598;
wire n_288;
wire n_404;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_0), .A2(n_70), .B1(n_503), .B2(n_591), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_1), .A2(n_40), .B1(n_465), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_2), .A2(n_207), .B1(n_348), .B2(n_626), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_3), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_4), .A2(n_265), .B1(n_403), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_5), .A2(n_98), .B1(n_368), .B2(n_413), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_6), .A2(n_24), .B1(n_126), .B2(n_312), .C1(n_495), .C2(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_7), .A2(n_125), .B1(n_504), .B2(n_509), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_8), .A2(n_99), .B1(n_668), .B2(n_777), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_9), .A2(n_232), .B1(n_463), .B2(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g786 ( .A(n_10), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_11), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_12), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_13), .A2(n_129), .B1(n_418), .B2(n_422), .C(n_424), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_14), .A2(n_31), .B1(n_353), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_15), .A2(n_146), .B1(n_774), .B2(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_16), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_17), .A2(n_151), .B1(n_428), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_18), .A2(n_134), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_19), .A2(n_38), .B1(n_645), .B2(n_704), .C(n_705), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_20), .A2(n_222), .B1(n_360), .B2(n_684), .C(n_686), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_21), .A2(n_133), .B1(n_559), .B2(n_651), .Y(n_843) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_22), .A2(n_88), .B1(n_294), .B2(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g822 ( .A(n_22), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_23), .A2(n_77), .B1(n_587), .B2(n_588), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_25), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_26), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_27), .A2(n_73), .B1(n_692), .B2(n_695), .C(n_698), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_28), .Y(n_287) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_29), .A2(n_214), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_30), .A2(n_259), .B1(n_368), .B2(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_32), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_33), .A2(n_191), .B1(n_352), .B2(n_591), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_34), .A2(n_137), .B1(n_522), .B2(n_656), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_35), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_36), .A2(n_42), .B1(n_366), .B2(n_556), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_37), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_39), .A2(n_161), .B1(n_354), .B2(n_376), .Y(n_676) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_41), .A2(n_91), .B1(n_294), .B2(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g823 ( .A(n_41), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_43), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_44), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_45), .A2(n_219), .B1(n_457), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_46), .A2(n_211), .B1(n_366), .B2(n_367), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_47), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_48), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_49), .A2(n_194), .B1(n_501), .B2(n_503), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_50), .A2(n_212), .B1(n_373), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_51), .A2(n_244), .B1(n_348), .B2(n_356), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_52), .A2(n_86), .B1(n_358), .B2(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_53), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_54), .A2(n_104), .B1(n_349), .B2(n_390), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_55), .A2(n_74), .B1(n_372), .B2(n_376), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_56), .A2(n_230), .B1(n_329), .B2(n_640), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_57), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_58), .A2(n_236), .B1(n_403), .B2(n_507), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_59), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_60), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_61), .A2(n_178), .B1(n_320), .B2(n_551), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_62), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_63), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_64), .A2(n_119), .B1(n_496), .B2(n_612), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_65), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_66), .A2(n_128), .B1(n_367), .B2(n_594), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_67), .A2(n_136), .B1(n_451), .B2(n_496), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_68), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_69), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_71), .A2(n_202), .B1(n_845), .B2(n_847), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_72), .A2(n_132), .B1(n_358), .B2(n_801), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_75), .B(n_328), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_76), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_78), .A2(n_93), .B1(n_403), .B2(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_79), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_80), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_81), .A2(n_116), .B1(n_356), .B2(n_360), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_82), .A2(n_225), .B1(n_329), .B2(n_544), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_83), .A2(n_187), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_84), .A2(n_141), .B1(n_614), .B2(n_615), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_85), .A2(n_154), .B1(n_531), .B2(n_533), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_87), .A2(n_156), .B1(n_354), .B2(n_590), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_89), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_90), .A2(n_169), .B1(n_591), .B2(n_882), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_92), .A2(n_682), .B1(n_712), .B2(n_713), .Y(n_681) );
INVx1_ASAP7_75t_L g712 ( .A(n_92), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_94), .Y(n_875) );
INVx1_ASAP7_75t_L g277 ( .A(n_95), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_96), .A2(n_192), .B1(n_690), .B2(n_729), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_97), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_100), .Y(n_608) );
INVx1_ASAP7_75t_L g274 ( .A(n_101), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_102), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_103), .A2(n_175), .B1(n_376), .B2(n_877), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_105), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_106), .A2(n_114), .B1(n_465), .B2(n_509), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_107), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_108), .A2(n_262), .B1(n_330), .B2(n_452), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_109), .A2(n_238), .B1(n_386), .B2(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_110), .A2(n_188), .B1(n_755), .B2(n_756), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_111), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_112), .A2(n_246), .B1(n_668), .B2(n_777), .Y(n_776) );
XOR2xp5_ASAP7_75t_L g825 ( .A(n_113), .B(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_115), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_117), .A2(n_120), .B1(n_452), .B2(n_551), .Y(n_550) );
OA22x2_ASAP7_75t_L g537 ( .A1(n_118), .A2(n_538), .B1(n_539), .B2(n_561), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_118), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_121), .B(n_580), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_122), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_123), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_124), .B(n_419), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_127), .Y(n_740) );
AOI22xp5_ASAP7_75t_SL g781 ( .A1(n_130), .A2(n_782), .B1(n_783), .B2(n_806), .Y(n_781) );
INVx1_ASAP7_75t_L g806 ( .A(n_130), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_131), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_135), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_138), .A2(n_170), .B1(n_756), .B2(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_139), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_140), .B(n_614), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_142), .Y(n_745) );
XNOR2x2_ASAP7_75t_L g750 ( .A(n_143), .B(n_751), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_144), .A2(n_162), .B1(n_348), .B2(n_352), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_145), .Y(n_395) );
INVx2_ASAP7_75t_L g278 ( .A(n_147), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_148), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_149), .A2(n_173), .B1(n_596), .B2(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_150), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_152), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_153), .B(n_547), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g427 ( .A1(n_155), .A2(n_218), .B1(n_252), .B2(n_312), .C1(n_328), .C2(n_428), .Y(n_427) );
AND2x6_ASAP7_75t_L g273 ( .A(n_157), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_157), .Y(n_816) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_158), .A2(n_223), .B1(n_294), .B2(n_298), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_159), .A2(n_198), .B1(n_367), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_160), .A2(n_229), .B1(n_618), .B2(n_620), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_163), .A2(n_240), .B1(n_772), .B2(n_774), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_164), .B(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_165), .Y(n_326) );
INVx1_ASAP7_75t_L g338 ( .A(n_166), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_167), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_168), .A2(n_263), .B1(n_397), .B2(n_622), .Y(n_621) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_171), .A2(n_271), .B(n_279), .C(n_824), .Y(n_270) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_172), .A2(n_227), .B1(n_453), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_174), .A2(n_242), .B1(n_372), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_176), .A2(n_241), .B1(n_520), .B2(n_525), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_177), .A2(n_256), .B1(n_354), .B2(n_504), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_179), .A2(n_186), .B1(n_531), .B2(n_544), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_180), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_181), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_182), .A2(n_206), .B1(n_366), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_183), .A2(n_250), .B1(n_520), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_184), .A2(n_269), .B1(n_650), .B2(n_651), .Y(n_649) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_185), .A2(n_248), .B1(n_294), .B2(n_295), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_189), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_189), .A2(n_857), .B1(n_859), .B2(n_884), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_190), .B(n_328), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_193), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_195), .A2(n_224), .B1(n_376), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_196), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_197), .A2(n_249), .B1(n_451), .B2(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_199), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_200), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_201), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_203), .A2(n_253), .B1(n_695), .B2(n_849), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_204), .A2(n_221), .B1(n_451), .B2(n_452), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_205), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_208), .A2(n_719), .B1(n_747), .B2(n_748), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_208), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_209), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_210), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_213), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_215), .B(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_216), .A2(n_381), .B1(n_430), .B2(n_431), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_216), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_217), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_220), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_223), .B(n_821), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_226), .Y(n_743) );
OA22x2_ASAP7_75t_L g602 ( .A1(n_228), .A2(n_603), .B1(n_604), .B2(n_628), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_228), .Y(n_603) );
INVx1_ASAP7_75t_L g516 ( .A(n_231), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_233), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_234), .Y(n_868) );
INVx1_ASAP7_75t_L g510 ( .A(n_235), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_237), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_239), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_243), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_245), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_247), .Y(n_866) );
INVx1_ASAP7_75t_L g819 ( .A(n_248), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_251), .Y(n_401) );
OA22x2_ASAP7_75t_SL g282 ( .A1(n_254), .A2(n_283), .B1(n_284), .B2(n_379), .Y(n_282) );
INVx1_ASAP7_75t_L g379 ( .A(n_254), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_255), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_257), .Y(n_576) );
INVx1_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_260), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_261), .Y(n_458) );
OA22x2_ASAP7_75t_L g437 ( .A1(n_264), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_264), .Y(n_438) );
AOI22x1_ASAP7_75t_L g567 ( .A1(n_266), .A2(n_568), .B1(n_597), .B2(n_598), .Y(n_567) );
INVx1_ASAP7_75t_L g597 ( .A(n_266), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_267), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_268), .Y(n_870) );
INVx2_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_274), .Y(n_815) );
OA21x2_ASAP7_75t_L g855 ( .A1(n_275), .A2(n_814), .B(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_600), .B1(n_809), .B2(n_810), .C(n_811), .Y(n_279) );
INVx1_ASAP7_75t_L g810 ( .A(n_280), .Y(n_810) );
XOR2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_434), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_380), .B1(n_432), .B2(n_433), .Y(n_281) );
INVx2_ASAP7_75t_L g432 ( .A(n_282), .Y(n_432) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_285), .B(n_345), .Y(n_284) );
NOR3xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_310), .C(n_332), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B1(n_304), .B2(n_305), .Y(n_286) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g443 ( .A(n_289), .Y(n_443) );
INVx1_ASAP7_75t_SL g744 ( .A(n_289), .Y(n_744) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx3_ASAP7_75t_L g485 ( .A(n_290), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_290), .A2(n_307), .B1(n_528), .B2(n_529), .C(n_530), .Y(n_527) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_290), .Y(n_832) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_299), .Y(n_290) );
INVx2_ASAP7_75t_L g359 ( .A(n_291), .Y(n_359) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_292), .B(n_297), .Y(n_309) );
AND2x2_ASAP7_75t_L g351 ( .A(n_292), .B(n_324), .Y(n_351) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g315 ( .A(n_293), .B(n_297), .Y(n_315) );
AND2x2_ASAP7_75t_L g325 ( .A(n_293), .B(n_303), .Y(n_325) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_296), .Y(n_298) );
INVx2_ASAP7_75t_L g324 ( .A(n_297), .Y(n_324) );
INVx1_ASAP7_75t_L g378 ( .A(n_297), .Y(n_378) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_300), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g354 ( .A(n_300), .B(n_351), .Y(n_354) );
AND2x4_ASAP7_75t_L g421 ( .A(n_300), .B(n_359), .Y(n_421) );
AND2x6_ASAP7_75t_L g423 ( .A(n_300), .B(n_309), .Y(n_423) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
INVx1_ASAP7_75t_L g323 ( .A(n_301), .Y(n_323) );
INVx1_ASAP7_75t_L g344 ( .A(n_301), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_301), .B(n_303), .Y(n_363) );
AND2x2_ASAP7_75t_L g316 ( .A(n_302), .B(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g370 ( .A(n_303), .B(n_344), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_305), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_305), .A2(n_832), .B1(n_862), .B2(n_863), .Y(n_861) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g746 ( .A(n_307), .Y(n_746) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g488 ( .A(n_308), .Y(n_488) );
AND2x4_ASAP7_75t_L g366 ( .A(n_309), .B(n_316), .Y(n_366) );
AND2x2_ASAP7_75t_L g375 ( .A(n_309), .B(n_370), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_309), .B(n_370), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_318), .B1(n_319), .B2(n_326), .C(n_327), .Y(n_310) );
OAI21xp5_ASAP7_75t_SL g785 ( .A1(n_311), .A2(n_786), .B(n_787), .Y(n_785) );
OAI21xp33_ASAP7_75t_SL g835 ( .A1(n_311), .A2(n_836), .B(n_837), .Y(n_835) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_313), .A2(n_490), .B(n_491), .Y(n_489) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g449 ( .A(n_314), .Y(n_449) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_314), .Y(n_575) );
INVx2_ASAP7_75t_L g607 ( .A(n_314), .Y(n_607) );
INVx2_ASAP7_75t_L g736 ( .A(n_314), .Y(n_736) );
AND2x6_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
AND2x4_ASAP7_75t_L g453 ( .A(n_315), .B(n_343), .Y(n_453) );
AND2x2_ASAP7_75t_L g350 ( .A(n_316), .B(n_351), .Y(n_350) );
AND2x6_ASAP7_75t_L g358 ( .A(n_316), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g429 ( .A(n_320), .Y(n_429) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_321), .Y(n_457) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_321), .Y(n_496) );
BUFx4f_ASAP7_75t_SL g544 ( .A(n_321), .Y(n_544) );
BUFx2_ASAP7_75t_L g739 ( .A(n_321), .Y(n_739) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g331 ( .A(n_323), .Y(n_331) );
INVx1_ASAP7_75t_L g337 ( .A(n_324), .Y(n_337) );
AND2x4_ASAP7_75t_L g330 ( .A(n_325), .B(n_331), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_325), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g531 ( .A(n_325), .B(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g839 ( .A(n_329), .Y(n_839) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx12f_ASAP7_75t_L g451 ( .A(n_330), .Y(n_451) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_330), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B1(n_338), .B2(n_339), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_334), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_334), .A2(n_708), .B1(n_870), .B2(n_871), .Y(n_869) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_SL g733 ( .A(n_335), .Y(n_733) );
INVx4_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_336), .A2(n_340), .B1(n_425), .B2(n_426), .Y(n_424) );
BUFx3_ASAP7_75t_L g459 ( .A(n_336), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_336), .A2(n_493), .B1(n_494), .B2(n_497), .Y(n_492) );
AND2x2_ASAP7_75t_L g522 ( .A(n_337), .B(n_362), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_339), .A2(n_459), .B1(n_582), .B2(n_583), .Y(n_581) );
OAI22xp5_ASAP7_75t_SL g838 ( .A1(n_339), .A2(n_839), .B1(n_840), .B2(n_841), .Y(n_838) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_340), .Y(n_709) );
OR2x6_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_364), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g346 ( .A(n_347), .B(n_355), .Y(n_346) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g587 ( .A(n_349), .Y(n_587) );
INVx3_ASAP7_75t_L g685 ( .A(n_349), .Y(n_685) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_349), .Y(n_755) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
BUFx2_ASAP7_75t_SL g469 ( .A(n_350), .Y(n_469) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_350), .Y(n_801) );
AND2x4_ASAP7_75t_L g361 ( .A(n_351), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g369 ( .A(n_351), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_351), .B(n_370), .Y(n_408) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g509 ( .A(n_354), .Y(n_509) );
INVx2_ASAP7_75t_L g657 ( .A(n_354), .Y(n_657) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_354), .Y(n_697) );
INVx4_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx4_ASAP7_75t_L g520 ( .A(n_357), .Y(n_520) );
INVx2_ASAP7_75t_SL g588 ( .A(n_357), .Y(n_588) );
INVx3_ASAP7_75t_L g797 ( .A(n_357), .Y(n_797) );
INVx11_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx11_ASAP7_75t_L g414 ( .A(n_358), .Y(n_414) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
BUFx2_ASAP7_75t_SL g472 ( .A(n_361), .Y(n_472) );
BUFx2_ASAP7_75t_L g504 ( .A(n_361), .Y(n_504) );
BUFx3_ASAP7_75t_L g591 ( .A(n_361), .Y(n_591) );
BUFx3_ASAP7_75t_L g620 ( .A(n_361), .Y(n_620) );
BUFx2_ASAP7_75t_SL g756 ( .A(n_361), .Y(n_756) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x6_ASAP7_75t_L g377 ( .A(n_363), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_371), .Y(n_364) );
INVx6_ASAP7_75t_L g404 ( .A(n_366), .Y(n_404) );
BUFx3_ASAP7_75t_L g525 ( .A(n_366), .Y(n_525) );
BUFx3_ASAP7_75t_L g594 ( .A(n_366), .Y(n_594) );
BUFx3_ASAP7_75t_L g701 ( .A(n_366), .Y(n_701) );
BUFx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g501 ( .A(n_369), .Y(n_501) );
BUFx3_ASAP7_75t_L g651 ( .A(n_369), .Y(n_651) );
BUFx3_ASAP7_75t_L g799 ( .A(n_369), .Y(n_799) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx5_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g463 ( .A(n_374), .Y(n_463) );
INVx3_ASAP7_75t_L g507 ( .A(n_374), .Y(n_507) );
INVx4_ASAP7_75t_L g556 ( .A(n_374), .Y(n_556) );
INVx2_ASAP7_75t_L g623 ( .A(n_374), .Y(n_623) );
BUFx3_ASAP7_75t_L g878 ( .A(n_374), .Y(n_878) );
INVx8_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx6_ASAP7_75t_SL g398 ( .A(n_377), .Y(n_398) );
INVx1_ASAP7_75t_L g532 ( .A(n_378), .Y(n_532) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
INVx1_ASAP7_75t_L g431 ( .A(n_381), .Y(n_431) );
AND4x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_399), .C(n_417), .D(n_427), .Y(n_381) );
NOR2xp33_ASAP7_75t_SL g382 ( .A(n_383), .B(n_391), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_388), .B2(n_389), .Y(n_383) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx3_ASAP7_75t_L g503 ( .A(n_387), .Y(n_503) );
INVx2_ASAP7_75t_L g849 ( .A(n_389), .Y(n_849) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_395), .B2(n_396), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_393), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
BUFx2_ASAP7_75t_R g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g465 ( .A(n_398), .Y(n_465) );
BUFx4f_ASAP7_75t_SL g596 ( .A(n_398), .Y(n_596) );
BUFx2_ASAP7_75t_L g690 ( .A(n_398), .Y(n_690) );
BUFx2_ASAP7_75t_L g847 ( .A(n_398), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_409), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_405), .B2(n_406), .Y(n_400) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g559 ( .A(n_404), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_404), .A2(n_478), .B1(n_763), .B2(n_764), .Y(n_762) );
INVx2_ASAP7_75t_L g804 ( .A(n_404), .Y(n_804) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g478 ( .A(n_407), .Y(n_478) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_415), .B2(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g760 ( .A(n_413), .Y(n_760) );
INVx5_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g475 ( .A(n_414), .Y(n_475) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_414), .Y(n_619) );
INVx4_ASAP7_75t_L g650 ( .A(n_414), .Y(n_650) );
INVx2_ASAP7_75t_SL g694 ( .A(n_414), .Y(n_694) );
INVx1_ASAP7_75t_L g626 ( .A(n_416), .Y(n_626) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx5_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g614 ( .A(n_420), .Y(n_614) );
INVx2_ASAP7_75t_L g643 ( .A(n_420), .Y(n_643) );
INVx2_ASAP7_75t_L g777 ( .A(n_420), .Y(n_777) );
INVx4_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g548 ( .A(n_423), .Y(n_548) );
BUFx4f_ASAP7_75t_L g645 ( .A(n_423), .Y(n_645) );
BUFx2_ASAP7_75t_L g668 ( .A(n_423), .Y(n_668) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
XOR2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_512), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_479), .B1(n_480), .B2(n_511), .Y(n_436) );
INVx2_ASAP7_75t_L g511 ( .A(n_437), .Y(n_511) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_460), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .C(n_454), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_443), .A2(n_487), .B1(n_571), .B2(n_572), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_450), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_448), .A2(n_535), .B(n_536), .Y(n_534) );
OAI21xp5_ASAP7_75t_SL g541 ( .A1(n_448), .A2(n_542), .B(n_543), .Y(n_541) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx4f_ASAP7_75t_SL g711 ( .A(n_451), .Y(n_711) );
INVx2_ASAP7_75t_L g789 ( .A(n_451), .Y(n_789) );
BUFx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_453), .Y(n_533) );
BUFx2_ASAP7_75t_SL g640 ( .A(n_453), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_458), .B2(n_459), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_466), .C(n_473), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_470), .B2(n_471), .Y(n_466) );
OAI221xp5_ASAP7_75t_SL g873 ( .A1(n_468), .A2(n_696), .B1(n_874), .B2(n_875), .C(n_876), .Y(n_873) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_476), .B1(n_477), .B2(n_478), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_478), .A2(n_699), .B1(n_700), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
XOR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_510), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_498), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .C(n_492), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_486), .B2(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g834 ( .A(n_488), .Y(n_834) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g727 ( .A(n_501), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_564), .B1(n_565), .B2(n_599), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g599 ( .A(n_514), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_537), .B1(n_562), .B2(n_563), .Y(n_514) );
INVx2_ASAP7_75t_SL g562 ( .A(n_515), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_515), .A2(n_562), .B1(n_566), .B2(n_567), .Y(n_565) );
XNOR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
NOR4xp75_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .C(n_527), .D(n_534), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_519), .B(n_521), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_524), .B(n_526), .Y(n_523) );
BUFx3_ASAP7_75t_L g551 ( .A(n_531), .Y(n_551) );
BUFx2_ASAP7_75t_L g612 ( .A(n_531), .Y(n_612) );
INVx1_ASAP7_75t_L g773 ( .A(n_531), .Y(n_773) );
BUFx2_ASAP7_75t_L g792 ( .A(n_531), .Y(n_792) );
INVx1_ASAP7_75t_SL g775 ( .A(n_533), .Y(n_775) );
INVx1_ASAP7_75t_L g563 ( .A(n_537), .Y(n_563) );
INVx1_ASAP7_75t_L g561 ( .A(n_539), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_552), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
INVx1_ASAP7_75t_L g577 ( .A(n_544), .Y(n_577) );
INVx1_ASAP7_75t_L g865 ( .A(n_544), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .C(n_550), .Y(n_545) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_SL g615 ( .A(n_548), .Y(n_615) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_556), .Y(n_729) );
INVx2_ASAP7_75t_L g846 ( .A(n_556), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_SL g598 ( .A(n_568), .Y(n_598) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_584), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .C(n_581), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_576), .B1(n_577), .B2(n_578), .C(n_579), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g638 ( .A(n_575), .Y(n_638) );
BUFx4f_ASAP7_75t_L g769 ( .A(n_580), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_592), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g809 ( .A(n_600), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_629), .B2(n_808), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g628 ( .A(n_604), .Y(n_628) );
NAND3x1_ASAP7_75t_L g604 ( .A(n_605), .B(n_616), .C(n_624), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_610), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B(n_609), .Y(n_606) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_607), .A2(n_663), .B(n_664), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g766 ( .A1(n_607), .A2(n_767), .B(n_768), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
BUFx2_ASAP7_75t_L g704 ( .A(n_614), .Y(n_704) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g808 ( .A(n_629), .Y(n_808) );
XNOR2xp5_ASAP7_75t_SL g629 ( .A(n_630), .B(n_679), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI22x1_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_659), .B2(n_678), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
XOR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_658), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_635), .B(n_647), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_641), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B(n_639), .Y(n_636) );
OAI222xp33_ASAP7_75t_L g864 ( .A1(n_638), .A2(n_839), .B1(n_865), .B2(n_866), .C1(n_867), .C2(n_868), .Y(n_864) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .C(n_646), .Y(n_641) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_648), .B(n_653), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx3_ASAP7_75t_L g678 ( .A(n_659), .Y(n_678) );
XOR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_677), .Y(n_659) );
NAND2x1_ASAP7_75t_SL g660 ( .A(n_661), .B(n_670), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .C(n_669), .Y(n_665) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B1(n_714), .B2(n_807), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g713 ( .A(n_682), .Y(n_713) );
AND4x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_691), .C(n_703), .D(n_710), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx4_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_696), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_758) );
INVx4_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_708), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g807 ( .A(n_714), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_778), .B2(n_779), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_749), .B2(n_750), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g748 ( .A(n_719), .Y(n_748) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_720), .B(n_730), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_728), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NOR3xp33_ASAP7_75t_SL g730 ( .A(n_731), .B(n_735), .C(n_742), .Y(n_730) );
OAI221xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_737), .B1(n_738), .B2(n_740), .C(n_741), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_742) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_752), .B(n_765), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_758), .C(n_762), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_757), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_770), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_776), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_784), .B(n_794), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_790), .Y(n_784) );
INVx3_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_802), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .Y(n_795) );
BUFx4f_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g883 ( .A(n_799), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
INVx1_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
NOR2x1_ASAP7_75t_L g812 ( .A(n_813), .B(n_817), .Y(n_812) );
OR2x2_ASAP7_75t_SL g887 ( .A(n_813), .B(n_818), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI322xp33_ASAP7_75t_L g824 ( .A1(n_815), .A2(n_825), .A3(n_851), .B1(n_855), .B2(n_857), .C1(n_858), .C2(n_885), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_815), .B(n_854), .Y(n_856) );
CKINVDCx16_ASAP7_75t_R g854 ( .A(n_816), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_842), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_835), .C(n_838), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B1(n_833), .B2(n_834), .Y(n_828) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
AND4x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .C(n_848), .D(n_850), .Y(n_842) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g884 ( .A(n_859), .Y(n_884) );
AND2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_872), .Y(n_859) );
NOR3xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_864), .C(n_869), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_879), .Y(n_872) );
INVx3_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NAND2xp5_ASAP7_75t_SL g879 ( .A(n_880), .B(n_881), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_887), .Y(n_886) );
endmodule