module real_jpeg_28628_n_17 (n_8, n_0, n_2, n_338, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_338;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_0),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_156),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_0),
.A2(n_99),
.B1(n_100),
.B2(n_156),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_0),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_302)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_62),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_62),
.B1(n_99),
.B2(n_100),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_2),
.A2(n_62),
.B1(n_159),
.B2(n_160),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_3),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_220),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_3),
.A2(n_99),
.B1(n_100),
.B2(n_220),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_3),
.A2(n_159),
.B1(n_160),
.B2(n_220),
.Y(n_333)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_5),
.A2(n_33),
.B1(n_35),
.B2(n_139),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_5),
.A2(n_99),
.B1(n_100),
.B2(n_139),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_5),
.A2(n_139),
.B1(n_159),
.B2(n_160),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_6),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_6),
.A2(n_33),
.B1(n_35),
.B2(n_116),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_6),
.A2(n_99),
.B1(n_100),
.B2(n_116),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_6),
.A2(n_116),
.B1(n_159),
.B2(n_160),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_8),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_201),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_8),
.A2(n_99),
.B1(n_100),
.B2(n_201),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_8),
.A2(n_159),
.B1(n_160),
.B2(n_201),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_34),
.B(n_35),
.C(n_38),
.D(n_42),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_59),
.B(n_63),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_99),
.B(n_101),
.C(n_102),
.D(n_106),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_10),
.B(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_10),
.A2(n_135),
.B(n_158),
.C(n_159),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_81),
.B1(n_159),
.B2(n_160),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_33),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_11),
.A2(n_44),
.B1(n_99),
.B2(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_44),
.B1(n_159),
.B2(n_160),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_55),
.B1(n_99),
.B2(n_100),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_55),
.B1(n_159),
.B2(n_160),
.Y(n_193)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_30),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_35),
.B(n_39),
.C(n_41),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_15),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_15),
.Y(n_105)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_329),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_316),
.B(n_328),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_280),
.A3(n_309),
.B1(n_314),
.B2(n_315),
.C(n_337),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_230),
.A3(n_269),
.B1(n_274),
.B2(n_279),
.C(n_338),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_180),
.C(n_226),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_147),
.B(n_179),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_122),
.B(n_146),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_94),
.B(n_121),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_68),
.B(n_93),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_27),
.B(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_37),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_37),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.A3(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_29),
.B(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_30),
.B(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_33),
.B(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_35),
.A2(n_100),
.A3(n_101),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_38),
.A2(n_41),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_38),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_38),
.A2(n_41),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_38),
.A2(n_41),
.B1(n_246),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_42),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_54),
.B(n_56),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_45),
.A2(n_56),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_45),
.A2(n_143),
.B1(n_178),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_45),
.A2(n_143),
.B1(n_203),
.B2(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_45),
.A2(n_143),
.B(n_255),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_58),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_53),
.C(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_50),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_50),
.A2(n_102),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_50),
.A2(n_102),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_50),
.A2(n_102),
.B1(n_258),
.B2(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_50),
.A2(n_102),
.B(n_321),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_51),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_54),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_67),
.B1(n_115),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_59),
.A2(n_67),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_59),
.A2(n_200),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_59),
.A2(n_76),
.B(n_219),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_84),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_66),
.A2(n_73),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx5_ASAP7_75t_SL g218 ( 
.A(n_66),
.Y(n_218)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_78),
.B(n_92),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_77),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_76),
.B(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_85),
.B(n_91),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_99),
.B(n_134),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_96),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_112),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_109),
.C(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_100),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_108),
.A2(n_128),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_108),
.A2(n_188),
.B1(n_215),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_108),
.A2(n_188),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_124),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_140),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_141),
.C(n_142),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_131),
.C(n_137),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_133),
.A2(n_165),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_133),
.A2(n_165),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_133),
.A2(n_165),
.B1(n_324),
.B2(n_333),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_135),
.B1(n_159),
.B2(n_160),
.Y(n_166)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_149),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_163),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_151),
.B(n_152),
.C(n_163),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_161),
.Y(n_184)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_173),
.C(n_176),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B(n_168),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_175),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_181),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_205),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_182),
.B(n_205),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_197),
.C(n_204),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_186),
.C(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_196),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B(n_190),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_191),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_194),
.B(n_195),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_194),
.A2(n_195),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_194),
.A2(n_237),
.B1(n_265),
.B2(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_194),
.A2(n_237),
.B1(n_292),
.B2(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_204),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_202),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_216),
.C(n_225),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_250),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_250),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_242),
.C(n_249),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_242),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_241),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_240),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_248),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_248),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_248),
.A2(n_263),
.B(n_266),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_268),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_260),
.B1(n_261),
.B2(n_267),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_256),
.B(n_259),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_259),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_259),
.A2(n_282),
.B1(n_283),
.B2(n_294),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_267),
.C(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_270),
.A2(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_297),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_297),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_294),
.C(n_295),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_291),
.B2(n_293),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_286),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_290),
.C(n_291),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_287),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_290),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_301),
.C(n_305),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_291),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_293),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_300),
.C(n_308),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_296),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_308),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_302),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_307),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_327),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_322),
.B1(n_325),
.B2(n_326),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_320),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_326),
.C(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_334),
.Y(n_335)
);


endmodule