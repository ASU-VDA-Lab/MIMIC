module fake_netlist_1_1053_n_877 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_115, n_97, n_80, n_107, n_60, n_114, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_113, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_877);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_113;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_877;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_769;
wire n_624;
wire n_725;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_771;
wire n_696;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_823;
wire n_822;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g116 ( .A(n_26), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_108), .Y(n_119) );
BUFx2_ASAP7_75t_SL g120 ( .A(n_56), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_92), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_43), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_24), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_42), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_22), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_8), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_12), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_21), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_18), .Y(n_131) );
NOR2xp67_ASAP7_75t_L g132 ( .A(n_91), .B(n_74), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_44), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_61), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_19), .Y(n_135) );
NOR2xp67_ASAP7_75t_L g136 ( .A(n_62), .B(n_97), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_81), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_75), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_18), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_28), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_20), .Y(n_143) );
INVxp33_ASAP7_75t_SL g144 ( .A(n_110), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_5), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_55), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_25), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_37), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_2), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_6), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_113), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_16), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_107), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_0), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_45), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_102), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_4), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_53), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_59), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_9), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_34), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_24), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_64), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_73), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_19), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_88), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_58), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_41), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_31), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_33), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_172), .Y(n_173) );
NAND2xp33_ASAP7_75t_R g174 ( .A(n_144), .B(n_27), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_146), .B(n_0), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_158), .B(n_1), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_146), .B(n_1), .Y(n_177) );
BUFx12f_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_121), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_158), .B(n_2), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_119), .B(n_122), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_118), .B(n_3), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_172), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_163), .B(n_169), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_124), .B(n_3), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_121), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_128), .Y(n_193) );
INVx6_ASAP7_75t_L g194 ( .A(n_120), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_128), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_118), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
BUFx8_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
NAND2xp33_ASAP7_75t_R g199 ( .A(n_144), .B(n_29), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_117), .B(n_4), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_194), .B(n_130), .Y(n_203) );
INVx4_ASAP7_75t_SL g204 ( .A(n_194), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_186), .B(n_139), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_198), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_193), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_186), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_186), .B(n_176), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_193), .Y(n_210) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_194), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_193), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_193), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_197), .B(n_143), .Y(n_214) );
INVxp33_ASAP7_75t_L g215 ( .A(n_197), .Y(n_215) );
NAND2xp33_ASAP7_75t_L g216 ( .A(n_181), .B(n_134), .Y(n_216) );
NAND2xp33_ASAP7_75t_L g217 ( .A(n_181), .B(n_138), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_186), .B(n_117), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_176), .B(n_153), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_179), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_193), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_194), .B(n_141), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_179), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_189), .B(n_153), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_194), .B(n_149), .Y(n_225) );
INVxp33_ASAP7_75t_SL g226 ( .A(n_189), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_193), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_198), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_178), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_178), .Y(n_230) );
AND2x6_ASAP7_75t_L g231 ( .A(n_177), .B(n_166), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_178), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_191), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_191), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_182), .B(n_129), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_177), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_185), .B(n_147), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_182), .B(n_138), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_183), .B(n_156), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_198), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_173), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_183), .B(n_152), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_184), .B(n_152), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_184), .B(n_156), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_199), .B1(n_174), .B2(n_200), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_244), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_208), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_244), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_234), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_206), .B(n_154), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_239), .B(n_187), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_241), .B(n_187), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_224), .B(n_180), .Y(n_260) );
AO21x1_ASAP7_75t_L g261 ( .A1(n_213), .A2(n_190), .B(n_192), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_215), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_233), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_234), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_244), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
INVxp67_ASAP7_75t_SL g267 ( .A(n_234), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_226), .B(n_180), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_209), .B(n_192), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_214), .B(n_175), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_219), .B(n_200), .Y(n_271) );
NOR2xp33_ASAP7_75t_R g272 ( .A(n_229), .B(n_133), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_246), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_235), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_247), .B(n_202), .Y(n_275) );
BUFx12f_ASAP7_75t_L g276 ( .A(n_230), .Y(n_276) );
INVx4_ASAP7_75t_L g277 ( .A(n_243), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_219), .B(n_202), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_209), .B(n_201), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_244), .Y(n_280) );
OR2x6_ASAP7_75t_L g281 ( .A(n_209), .B(n_201), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_230), .B(n_154), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_208), .A2(n_168), .B1(n_157), .B2(n_126), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_236), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_244), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_248), .B(n_165), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_232), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_236), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
BUFx8_ASAP7_75t_SL g292 ( .A(n_276), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_279), .B(n_231), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
OAI22xp5_ASAP7_75t_SL g295 ( .A1(n_287), .A2(n_151), .B1(n_123), .B2(n_131), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
AOI21x1_ASAP7_75t_L g297 ( .A1(n_261), .A2(n_213), .B(n_221), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_279), .B(n_231), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_268), .B(n_206), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_279), .A2(n_205), .B1(n_231), .B2(n_218), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_262), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_254), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_279), .B(n_231), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_264), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_263), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_259), .A2(n_228), .B(n_211), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_263), .Y(n_307) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_270), .B(n_250), .C(n_271), .Y(n_308) );
BUFx4f_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_269), .B(n_237), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_269), .B(n_231), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_256), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_269), .B(n_231), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_256), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_278), .A2(n_240), .B1(n_237), .B2(n_218), .C(n_242), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_274), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_269), .B(n_231), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_252), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_309), .B(n_264), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_323), .B(n_281), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_316), .B(n_260), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_297), .A2(n_261), .B(n_255), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_323), .B(n_281), .Y(n_333) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_297), .A2(n_250), .B(n_246), .Y(n_334) );
OAI21x1_ASAP7_75t_L g335 ( .A1(n_306), .A2(n_255), .B(n_251), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_308), .A2(n_205), .B1(n_275), .B2(n_218), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_302), .A2(n_255), .B(n_251), .Y(n_337) );
OAI21x1_ASAP7_75t_L g338 ( .A1(n_305), .A2(n_265), .B(n_251), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_301), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_309), .A2(n_283), .B1(n_289), .B2(n_282), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_305), .A2(n_280), .B(n_265), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_308), .A2(n_284), .B1(n_288), .B2(n_218), .Y(n_342) );
AO21x2_ASAP7_75t_L g343 ( .A1(n_307), .A2(n_246), .B(n_195), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_307), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_310), .Y(n_345) );
AOI21xp33_ASAP7_75t_SL g346 ( .A1(n_295), .A2(n_286), .B(n_257), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_311), .B(n_284), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_310), .A2(n_265), .B(n_280), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_311), .B(n_252), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_317), .A2(n_288), .B(n_252), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_317), .A2(n_290), .B(n_253), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_319), .A2(n_228), .B(n_267), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_319), .A2(n_285), .B(n_280), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_326), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_342), .A2(n_309), .B(n_322), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_340), .A2(n_309), .B1(n_295), .B2(n_299), .Y(n_357) );
OAI211xp5_ASAP7_75t_L g358 ( .A1(n_346), .A2(n_272), .B(n_318), .C(n_301), .Y(n_358) );
AOI221x1_ASAP7_75t_SL g359 ( .A1(n_330), .A2(n_148), .B1(n_129), .B2(n_162), .C(n_164), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_331), .A2(n_195), .B(n_221), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_342), .A2(n_289), .B(n_256), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_347), .B(n_320), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_333), .A2(n_205), .B1(n_298), .B2(n_303), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g364 ( .A1(n_339), .A2(n_291), .B1(n_293), .B2(n_298), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_335), .A2(n_256), .B(n_243), .Y(n_365) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_339), .A2(n_291), .B1(n_135), .B2(n_300), .C(n_164), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_329), .A2(n_303), .B1(n_293), .B2(n_321), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_333), .A2(n_205), .B1(n_312), .B2(n_321), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_336), .A2(n_314), .B1(n_312), .B2(n_325), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_354), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_327), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_347), .B(n_314), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_328), .A2(n_148), .B1(n_162), .B2(n_127), .C1(n_140), .C2(n_142), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_327), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_354), .B(n_296), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_333), .A2(n_205), .B1(n_217), .B2(n_216), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_346), .B(n_205), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_335), .A2(n_352), .B(n_334), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_333), .A2(n_205), .B1(n_120), .B2(n_304), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_328), .B(n_296), .Y(n_383) );
AO31x2_ASAP7_75t_L g384 ( .A1(n_332), .A2(n_249), .A3(n_225), .B(n_222), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_332), .B(n_296), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_327), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_335), .A2(n_256), .B(n_264), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_329), .A2(n_238), .B1(n_245), .B2(n_223), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_329), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_329), .A2(n_238), .B1(n_245), .B2(n_223), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_329), .A2(n_304), .B1(n_325), .B2(n_292), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_367), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_357), .A2(n_336), .B1(n_345), .B2(n_344), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_355), .B(n_344), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_377), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_359), .B(n_345), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
INVx5_ASAP7_75t_L g399 ( .A(n_373), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_359), .B(n_349), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_371), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_375), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_372), .B(n_334), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_377), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_334), .Y(n_406) );
INVx4_ASAP7_75t_L g407 ( .A(n_373), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_375), .B(n_334), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_389), .B(n_343), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_383), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_358), .A2(n_349), .B1(n_350), .B2(n_351), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_389), .B(n_350), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_343), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_378), .B(n_385), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_366), .B(n_349), .Y(n_417) );
INVx4_ASAP7_75t_R g418 ( .A(n_362), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_362), .B(n_343), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_360), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_386), .B(n_343), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_360), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_360), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_360), .Y(n_428) );
INVx4_ASAP7_75t_R g429 ( .A(n_391), .Y(n_429) );
BUFx3_ASAP7_75t_L g430 ( .A(n_386), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_376), .B(n_349), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_386), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_374), .B(n_220), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_388), .B(n_331), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_384), .B(n_351), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_388), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_384), .B(n_331), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_390), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_380), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_390), .B(n_220), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_384), .B(n_220), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_356), .B(n_353), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
OR2x6_ASAP7_75t_L g445 ( .A(n_368), .B(n_353), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_368), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_364), .A2(n_304), .B1(n_325), .B2(n_324), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_370), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_363), .B(n_220), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_387), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_382), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_381), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_361), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_365), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_369), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_379), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_398), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_416), .B(n_132), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_399), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_397), .B(n_136), .C(n_125), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_416), .B(n_353), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_412), .B(n_337), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_414), .B(n_337), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_407), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_392), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_392), .Y(n_466) );
AOI33xp33_ASAP7_75t_L g467 ( .A1(n_455), .A2(n_116), .A3(n_145), .B1(n_150), .B2(n_155), .B3(n_167), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_399), .Y(n_468) );
NOR2x1_ASAP7_75t_SL g469 ( .A(n_407), .B(n_315), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_425), .B(n_196), .Y(n_470) );
INVx5_ASAP7_75t_L g471 ( .A(n_407), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_410), .B(n_196), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_393), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_410), .B(n_196), .Y(n_475) );
OAI22xp5_ASAP7_75t_SL g476 ( .A1(n_429), .A2(n_165), .B1(n_170), .B2(n_171), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_395), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_395), .B(n_5), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_401), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_417), .A2(n_170), .B1(n_171), .B2(n_304), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_415), .B(n_196), .Y(n_481) );
OAI21x1_ASAP7_75t_L g482 ( .A1(n_452), .A2(n_450), .B(n_428), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_6), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_399), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_401), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_396), .B(n_7), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_400), .B(n_7), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_415), .B(n_8), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_414), .B(n_337), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_407), .Y(n_490) );
INVx5_ASAP7_75t_SL g491 ( .A(n_445), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_403), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_435), .B(n_348), .Y(n_493) );
OAI31xp33_ASAP7_75t_L g494 ( .A1(n_451), .A2(n_203), .A3(n_223), .B(n_245), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_435), .B(n_338), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_438), .B(n_338), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_421), .B(n_223), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_438), .B(n_348), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_421), .B(n_245), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_424), .Y(n_500) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_450), .A2(n_348), .B(n_341), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_451), .B(n_10), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_412), .B(n_338), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_403), .B(n_10), .Y(n_504) );
OAI33xp33_ASAP7_75t_L g505 ( .A1(n_455), .A2(n_227), .A3(n_210), .B1(n_212), .B2(n_15), .B3(n_16), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_412), .B(n_341), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_399), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_418), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_405), .B(n_11), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_436), .A2(n_325), .B1(n_313), .B2(n_324), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_399), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_405), .B(n_13), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_418), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_412), .B(n_341), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_393), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_399), .B(n_313), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_406), .B(n_13), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_402), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_402), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_419), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_430), .B(n_313), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_419), .B(n_14), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_436), .B(n_315), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_442), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_439), .B(n_14), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_406), .B(n_15), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_430), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_394), .B(n_17), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_430), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_442), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_436), .B(n_17), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_456), .A2(n_324), .B(n_227), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_409), .B(n_20), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_394), .B(n_21), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_441), .B(n_315), .Y(n_535) );
OAI21xp33_ASAP7_75t_SL g536 ( .A1(n_445), .A2(n_277), .B(n_23), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_428), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_449), .B(n_22), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_420), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_409), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_446), .B(n_23), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_449), .B(n_25), .Y(n_542) );
AOI33xp33_ASAP7_75t_L g543 ( .A1(n_446), .A2(n_26), .A3(n_212), .B1(n_210), .B2(n_273), .B3(n_285), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_422), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_432), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_441), .Y(n_546) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_423), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_437), .B(n_173), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_404), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_448), .B(n_173), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_448), .B(n_173), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_437), .A2(n_173), .B1(n_188), .B2(n_290), .C(n_253), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_444), .B(n_188), .Y(n_553) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_434), .B(n_315), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_447), .A2(n_188), .B1(n_290), .B2(n_253), .C(n_210), .Y(n_555) );
INVx5_ASAP7_75t_L g556 ( .A(n_432), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_404), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_448), .B(n_188), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_456), .A2(n_188), .B1(n_315), .B2(n_253), .Y(n_559) );
INVx2_ASAP7_75t_SL g560 ( .A(n_429), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_423), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_444), .B(n_188), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_411), .B(n_290), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_560), .A2(n_413), .B1(n_445), .B2(n_440), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_465), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_476), .B(n_433), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_466), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_479), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_517), .B(n_413), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_520), .B(n_408), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_536), .A2(n_453), .B(n_452), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_560), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_517), .B(n_413), .Y(n_573) );
AOI322xp5_ASAP7_75t_L g574 ( .A1(n_458), .A2(n_411), .A3(n_413), .B1(n_426), .B2(n_427), .C1(n_454), .C2(n_440), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_473), .Y(n_575) );
NOR2xp33_ASAP7_75t_R g576 ( .A(n_471), .B(n_426), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_526), .B(n_445), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_470), .A2(n_454), .B1(n_427), .B2(n_440), .C(n_408), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_458), .B(n_440), .Y(n_579) );
BUFx3_ASAP7_75t_L g580 ( .A(n_490), .Y(n_580) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_464), .B(n_434), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_549), .B(n_440), .Y(n_582) );
CKINVDCx8_ASAP7_75t_R g583 ( .A(n_471), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_546), .A2(n_445), .B1(n_443), .B2(n_315), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_473), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_485), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_502), .B(n_30), .Y(n_587) );
INVx5_ASAP7_75t_L g588 ( .A(n_471), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_515), .Y(n_589) );
AND3x1_ASAP7_75t_L g590 ( .A(n_502), .B(n_212), .C(n_35), .Y(n_590) );
INVx6_ASAP7_75t_L g591 ( .A(n_471), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_443), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_515), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_519), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_457), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_464), .B(n_277), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_557), .B(n_443), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_474), .B(n_443), .Y(n_598) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_460), .B(n_277), .C(n_273), .D(n_285), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_464), .B(n_277), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_540), .B(n_457), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_539), .Y(n_603) );
NAND4xp75_ASAP7_75t_SL g604 ( .A(n_494), .B(n_32), .C(n_36), .D(n_38), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_474), .B(n_443), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_477), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_500), .B(n_39), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_533), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_547), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_500), .B(n_244), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_525), .Y(n_611) );
INVx6_ASAP7_75t_L g612 ( .A(n_459), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_522), .B(n_40), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_478), .B(n_46), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_561), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_507), .B(n_47), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_531), .B(n_524), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_530), .B(n_48), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_461), .B(n_49), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_461), .B(n_50), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_507), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_463), .B(n_51), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_463), .B(n_52), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_489), .B(n_54), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_561), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_489), .B(n_57), .Y(n_626) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_459), .B(n_207), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_518), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_469), .A2(n_256), .B(n_211), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_511), .B(n_60), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_486), .B(n_63), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_519), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_468), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_493), .B(n_207), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_504), .Y(n_635) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_508), .B(n_211), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_539), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_468), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_484), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_544), .B(n_65), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_544), .B(n_538), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_493), .B(n_207), .Y(n_642) );
OAI33xp33_ASAP7_75t_L g643 ( .A1(n_528), .A2(n_66), .A3(n_67), .B1(n_68), .B2(n_69), .B3(n_70), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_488), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_542), .B(n_71), .Y(n_645) );
BUFx3_ASAP7_75t_L g646 ( .A(n_484), .Y(n_646) );
INVx4_ASAP7_75t_L g647 ( .A(n_511), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_537), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_495), .B(n_207), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_496), .B(n_72), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_496), .B(n_76), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_541), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_498), .B(n_77), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_495), .B(n_207), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_550), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_498), .B(n_79), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_472), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_475), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_487), .B(n_207), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_491), .A2(n_80), .B1(n_83), .B2(n_84), .Y(n_660) );
NAND4xp25_ASAP7_75t_SL g661 ( .A(n_467), .B(n_85), .C(n_86), .D(n_87), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_509), .B(n_89), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_512), .B(n_90), .Y(n_663) );
INVx3_ASAP7_75t_L g664 ( .A(n_462), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_487), .B(n_93), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_483), .B(n_94), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_516), .Y(n_667) );
INVx4_ASAP7_75t_L g668 ( .A(n_516), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_537), .B(n_96), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_467), .B(n_98), .Y(n_670) );
AND2x4_ASAP7_75t_SL g671 ( .A(n_513), .B(n_99), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_481), .B(n_100), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_534), .B(n_103), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_551), .B(n_104), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_558), .B(n_105), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_543), .B(n_109), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_527), .B(n_111), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_545), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_497), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_543), .B(n_112), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_529), .B(n_114), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_527), .B(n_115), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_545), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_641), .B(n_554), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_554), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_573), .B(n_523), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_565), .Y(n_688) );
OAI33xp33_ASAP7_75t_L g689 ( .A1(n_606), .A2(n_499), .A3(n_563), .B1(n_510), .B2(n_548), .B3(n_553), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_567), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_595), .B(n_523), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_595), .B(n_523), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_572), .B(n_480), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_602), .B(n_506), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_611), .B(n_529), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_592), .B(n_491), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_588), .B(n_514), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_580), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_602), .B(n_514), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_568), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_609), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_588), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_586), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_600), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_576), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_637), .B(n_491), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_643), .A2(n_505), .B(n_506), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_628), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_577), .B(n_514), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_570), .B(n_506), .Y(n_710) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_581), .B(n_462), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_655), .B(n_503), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_570), .B(n_462), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_617), .B(n_503), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_655), .B(n_503), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_615), .B(n_562), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_598), .B(n_535), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g718 ( .A(n_668), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_661), .A2(n_535), .B1(n_516), .B2(n_521), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_625), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_605), .B(n_556), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_574), .B(n_559), .C(n_552), .D(n_555), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_668), .B(n_556), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_583), .A2(n_559), .B1(n_556), .B2(n_532), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_652), .B(n_482), .Y(n_725) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_647), .B(n_646), .Y(n_726) );
OR2x6_ASAP7_75t_L g727 ( .A(n_591), .B(n_482), .Y(n_727) );
OR2x6_ASAP7_75t_L g728 ( .A(n_591), .B(n_521), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_608), .B(n_501), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_648), .B(n_501), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_588), .A2(n_556), .B1(n_521), .B2(n_211), .Y(n_731) );
NAND4xp25_ASAP7_75t_L g732 ( .A(n_566), .B(n_204), .C(n_579), .D(n_584), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_597), .B(n_204), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_647), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_575), .Y(n_735) );
AND2x2_ASAP7_75t_SL g736 ( .A(n_671), .B(n_204), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_585), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_582), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_582), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_661), .A2(n_204), .B1(n_599), .B2(n_670), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_635), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_597), .B(n_204), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_667), .B(n_678), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_679), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_683), .B(n_621), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_634), .B(n_642), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_591), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_644), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_578), .B(n_589), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_638), .B(n_639), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_657), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_593), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_638), .B(n_639), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_587), .A2(n_590), .B1(n_670), .B2(n_658), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_578), .B(n_632), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_594), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_634), .B(n_654), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_633), .B(n_664), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_610), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_664), .B(n_656), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_631), .B(n_612), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_642), .B(n_654), .Y(n_762) );
INVx2_ASAP7_75t_SL g763 ( .A(n_588), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_649), .B(n_610), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_623), .B(n_626), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_649), .B(n_564), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_612), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_627), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_571), .B(n_659), .Y(n_769) );
OR2x2_ASAP7_75t_L g770 ( .A(n_710), .B(n_650), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_688), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_754), .A2(n_665), .B1(n_660), .B2(n_571), .C(n_599), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_718), .A2(n_711), .B1(n_705), .B2(n_719), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_690), .Y(n_774) );
XOR2xp5_ASAP7_75t_L g775 ( .A(n_712), .B(n_651), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_700), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_703), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_732), .A2(n_612), .B1(n_653), .B2(n_622), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_704), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_729), .B(n_659), .Y(n_780) );
OAI21xp33_ASAP7_75t_L g781 ( .A1(n_729), .A2(n_660), .B(n_665), .Y(n_781) );
BUFx12f_ASAP7_75t_L g782 ( .A(n_736), .Y(n_782) );
OAI22xp33_ASAP7_75t_SL g783 ( .A1(n_726), .A2(n_640), .B1(n_630), .B2(n_616), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_711), .A2(n_643), .B1(n_666), .B2(n_645), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_698), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_701), .Y(n_786) );
AOI21xp33_ASAP7_75t_L g787 ( .A1(n_768), .A2(n_673), .B(n_676), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_708), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_769), .A2(n_680), .B1(n_676), .B2(n_673), .C(n_672), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_723), .Y(n_790) );
NOR5xp2_ASAP7_75t_SL g791 ( .A(n_724), .B(n_604), .C(n_636), .D(n_630), .E(n_616), .Y(n_791) );
O2A1O1Ixp33_ASAP7_75t_L g792 ( .A1(n_751), .A2(n_680), .B(n_614), .C(n_618), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_741), .B(n_613), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_685), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_748), .B(n_744), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_735), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_689), .A2(n_624), .B1(n_663), .B2(n_662), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_714), .B(n_619), .Y(n_798) );
NOR2x1_ASAP7_75t_L g799 ( .A(n_728), .B(n_604), .Y(n_799) );
INVx1_ASAP7_75t_SL g800 ( .A(n_750), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_738), .B(n_620), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_724), .A2(n_607), .B1(n_681), .B2(n_669), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_765), .A2(n_682), .B1(n_677), .B2(n_675), .Y(n_803) );
AOI32xp33_ASAP7_75t_SL g804 ( .A1(n_695), .A2(n_674), .A3(n_669), .B1(n_601), .B2(n_596), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_709), .B(n_674), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_725), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_725), .B(n_629), .C(n_596), .Y(n_807) );
INVx3_ASAP7_75t_L g808 ( .A(n_728), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_L g809 ( .A1(n_693), .A2(n_601), .B(n_629), .C(n_761), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_737), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_720), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_740), .A2(n_728), .B1(n_715), .B2(n_768), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_707), .A2(n_694), .B1(n_699), .B2(n_746), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_689), .A2(n_684), .B1(n_766), .B2(n_722), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_769), .A2(n_699), .B1(n_694), .B2(n_749), .C(n_755), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_766), .A2(n_713), .B1(n_710), .B2(n_759), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_814), .A2(n_782), .B1(n_813), .B2(n_773), .Y(n_817) );
AOI321xp33_ASAP7_75t_L g818 ( .A1(n_813), .A2(n_713), .A3(n_749), .B1(n_755), .B2(n_686), .C(n_707), .Y(n_818) );
OAI21xp33_ASAP7_75t_L g819 ( .A1(n_815), .A2(n_745), .B(n_758), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_773), .A2(n_734), .B1(n_763), .B2(n_702), .Y(n_820) );
XOR2x2_ASAP7_75t_L g821 ( .A(n_775), .B(n_736), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_816), .B(n_739), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_784), .B(n_767), .C(n_727), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_780), .B(n_794), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_802), .A2(n_747), .B1(n_727), .B2(n_697), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_785), .B(n_753), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_796), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_790), .B(n_721), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_786), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_812), .B(n_727), .C(n_691), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_780), .B(n_764), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_795), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_806), .B(n_764), .Y(n_833) );
INVx1_ASAP7_75t_SL g834 ( .A(n_800), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_771), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_803), .A2(n_762), .B1(n_757), .B2(n_731), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_799), .A2(n_731), .B(n_716), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_774), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_776), .B(n_743), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_789), .A2(n_772), .B1(n_781), .B2(n_812), .Y(n_840) );
XNOR2x1_ASAP7_75t_L g841 ( .A(n_802), .B(n_696), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_833), .Y(n_842) );
AOI322xp5_ASAP7_75t_L g843 ( .A1(n_817), .A2(n_778), .A3(n_793), .B1(n_797), .B2(n_809), .C1(n_787), .C2(n_808), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g844 ( .A1(n_817), .A2(n_792), .B(n_808), .C(n_798), .Y(n_844) );
OAI32xp33_ASAP7_75t_L g845 ( .A1(n_820), .A2(n_770), .A3(n_804), .B1(n_777), .B2(n_788), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_834), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g847 ( .A1(n_840), .A2(n_779), .B1(n_787), .B2(n_811), .C(n_783), .Y(n_847) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_821), .B(n_805), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_829), .Y(n_849) );
AO21x1_ASAP7_75t_L g850 ( .A1(n_825), .A2(n_791), .B(n_801), .Y(n_850) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_825), .B(n_807), .Y(n_851) );
CKINVDCx6p67_ASAP7_75t_R g852 ( .A(n_828), .Y(n_852) );
INVx2_ASAP7_75t_SL g853 ( .A(n_826), .Y(n_853) );
AOI21xp33_ASAP7_75t_L g854 ( .A1(n_840), .A2(n_733), .B(n_742), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_845), .A2(n_836), .B1(n_830), .B2(n_823), .C(n_819), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_846), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_L g857 ( .A1(n_850), .A2(n_837), .B(n_822), .C(n_824), .Y(n_857) );
O2A1O1Ixp33_ASAP7_75t_L g858 ( .A1(n_844), .A2(n_832), .B(n_838), .C(n_835), .Y(n_858) );
NOR2x2_ASAP7_75t_L g859 ( .A(n_848), .B(n_818), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_851), .A2(n_841), .B1(n_826), .B2(n_831), .Y(n_860) );
INVx2_ASAP7_75t_SL g861 ( .A(n_852), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_856), .B(n_843), .Y(n_862) );
NOR3xp33_ASAP7_75t_L g863 ( .A(n_855), .B(n_847), .C(n_854), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_861), .B(n_853), .Y(n_864) );
OAI31xp33_ASAP7_75t_L g865 ( .A1(n_857), .A2(n_854), .A3(n_843), .B(n_842), .Y(n_865) );
NAND4xp25_ASAP7_75t_L g866 ( .A(n_865), .B(n_860), .C(n_858), .D(n_859), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_864), .Y(n_867) );
O2A1O1Ixp33_ASAP7_75t_L g868 ( .A1(n_862), .A2(n_849), .B(n_839), .C(n_827), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_867), .B(n_863), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_868), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_869), .Y(n_871) );
NOR4xp75_ASAP7_75t_L g872 ( .A(n_869), .B(n_866), .C(n_742), .D(n_733), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_871), .A2(n_870), .B1(n_827), .B2(n_706), .Y(n_873) );
OAI22x1_ASAP7_75t_L g874 ( .A1(n_872), .A2(n_870), .B1(n_810), .B2(n_760), .Y(n_874) );
OAI21xp33_ASAP7_75t_SL g875 ( .A1(n_873), .A2(n_692), .B(n_730), .Y(n_875) );
AO221x1_ASAP7_75t_L g876 ( .A1(n_875), .A2(n_874), .B1(n_752), .B2(n_756), .C(n_687), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_876), .A2(n_717), .B1(n_730), .B2(n_716), .Y(n_877) );
endmodule