module fake_netlist_1_12503_n_715 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_715);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_715;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g106 ( .A(n_101), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_48), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_53), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
HB1xp67_ASAP7_75t_SL g112 ( .A(n_86), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_90), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_43), .B(n_37), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_23), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_61), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_10), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_35), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_41), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_105), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_11), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_24), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_51), .Y(n_133) );
INVxp33_ASAP7_75t_L g134 ( .A(n_10), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_7), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
INVx1_ASAP7_75t_SL g137 ( .A(n_42), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_12), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_63), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_32), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_1), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_4), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_102), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_9), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_39), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_70), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_5), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_20), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_138), .Y(n_152) );
AOI22xp33_ASAP7_75t_SL g153 ( .A1(n_123), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_107), .A2(n_52), .B(n_103), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_108), .B(n_2), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_129), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_138), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_138), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_108), .B(n_3), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_107), .A2(n_54), .B(n_100), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_134), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_145), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_145), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_117), .Y(n_167) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_117), .A2(n_56), .B(n_99), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
OR2x2_ASAP7_75t_L g171 ( .A(n_163), .B(n_164), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_156), .Y(n_175) );
XOR2xp5_ASAP7_75t_L g176 ( .A(n_153), .B(n_123), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g177 ( .A(n_162), .B(n_124), .C(n_130), .Y(n_177) );
OR2x6_ASAP7_75t_L g178 ( .A(n_155), .B(n_116), .Y(n_178) );
NOR2xp33_ASAP7_75t_SL g179 ( .A(n_167), .B(n_129), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_167), .B(n_140), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
INVxp67_ASAP7_75t_SL g185 ( .A(n_163), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_155), .A2(n_149), .B1(n_116), .B2(n_146), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_154), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_163), .B(n_139), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_164), .B(n_106), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_149), .B1(n_136), .B2(n_142), .Y(n_191) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_162), .B(n_144), .C(n_139), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_159), .B(n_148), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_154), .B(n_118), .C(n_119), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_194), .B(n_159), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_185), .B(n_159), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_181), .A2(n_166), .B(n_119), .C(n_118), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_176), .A2(n_153), .B1(n_150), .B2(n_148), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_178), .B(n_115), .Y(n_200) );
NOR2xp67_ASAP7_75t_L g201 ( .A(n_170), .B(n_115), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_178), .Y(n_202) );
NAND2x1p5_ASAP7_75t_L g203 ( .A(n_170), .B(n_154), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_185), .B(n_150), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_183), .B(n_137), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_179), .B(n_109), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_192), .A2(n_110), .B1(n_121), .B2(n_122), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_178), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_171), .B(n_112), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_175), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_183), .B(n_121), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_182), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_188), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_171), .B(n_111), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_178), .B(n_188), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_178), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_178), .B(n_122), .Y(n_219) );
AND2x6_ASAP7_75t_SL g220 ( .A(n_189), .B(n_113), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_179), .B(n_125), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_182), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_182), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_181), .A2(n_141), .B(n_133), .C(n_143), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_177), .B1(n_182), .B2(n_190), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_177), .A2(n_110), .B1(n_147), .B2(n_132), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_186), .B(n_110), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_184), .A2(n_110), .B1(n_126), .B2(n_128), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_191), .A2(n_131), .B(n_127), .C(n_120), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_202), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_200), .A2(n_187), .B1(n_176), .B2(n_184), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_197), .B(n_190), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_223), .A2(n_187), .B(n_195), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_217), .B(n_187), .Y(n_234) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_215), .A2(n_195), .B(n_114), .C(n_120), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_223), .A2(n_187), .B(n_161), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_219), .B(n_110), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_219), .B(n_114), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_210), .B(n_152), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_161), .B1(n_154), .B2(n_168), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_214), .Y(n_243) );
NOR3xp33_ASAP7_75t_L g244 ( .A(n_199), .B(n_157), .C(n_169), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_219), .B(n_154), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_204), .B(n_161), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_200), .A2(n_168), .B1(n_161), .B2(n_169), .Y(n_247) );
NOR2xp67_ASAP7_75t_L g248 ( .A(n_212), .B(n_6), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_202), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_204), .B(n_161), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_196), .B(n_7), .Y(n_253) );
INVx4_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_225), .B(n_168), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_218), .A2(n_168), .B1(n_157), .B2(n_169), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_206), .A2(n_168), .B(n_180), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_211), .A2(n_157), .B1(n_152), .B2(n_158), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_206), .A2(n_172), .B(n_180), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_207), .A2(n_172), .B(n_180), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_254), .B(n_227), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_203), .B(n_221), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_244), .A2(n_224), .B(n_198), .C(n_229), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_257), .A2(n_203), .B(n_208), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_243), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_207), .B(n_222), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_232), .B(n_227), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_249), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_254), .B(n_227), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_252), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_253), .B(n_216), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_203), .B(n_201), .Y(n_273) );
AO31x2_ASAP7_75t_L g274 ( .A1(n_255), .A2(n_213), .A3(n_222), .B(n_205), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_247), .A2(n_201), .B(n_214), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_235), .B(n_226), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_233), .A2(n_209), .B(n_226), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_241), .A2(n_228), .B(n_172), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_236), .A2(n_173), .B(n_152), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_231), .B(n_212), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_246), .A2(n_173), .B(n_193), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_251), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_259), .A2(n_173), .B(n_158), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_234), .B(n_220), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_281), .A2(n_235), .B(n_240), .Y(n_285) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_275), .A2(n_238), .B(n_239), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_275), .A2(n_240), .B(n_260), .Y(n_287) );
OAI21x1_ASAP7_75t_SL g288 ( .A1(n_282), .A2(n_258), .B(n_248), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_280), .A2(n_199), .B1(n_253), .B2(n_234), .Y(n_289) );
AOI21xp33_ASAP7_75t_SL g290 ( .A1(n_280), .A2(n_250), .B(n_9), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_272), .B(n_250), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_279), .A2(n_252), .B(n_160), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_282), .A2(n_230), .B(n_160), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_282), .A2(n_230), .B(n_193), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_279), .A2(n_158), .B(n_160), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_266), .A2(n_230), .B(n_160), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_273), .A2(n_160), .B(n_158), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_261), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_270), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_267), .B(n_230), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_265), .Y(n_302) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_273), .A2(n_160), .B(n_158), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_262), .A2(n_160), .B(n_158), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_284), .B(n_220), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_302), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_303), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_302), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_303), .Y(n_309) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_304), .A2(n_262), .B(n_264), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_304), .A2(n_264), .B(n_283), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_303), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_303), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_299), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_303), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_297), .Y(n_316) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_304), .A2(n_283), .B(n_278), .Y(n_317) );
AOI21xp33_ASAP7_75t_L g318 ( .A1(n_290), .A2(n_263), .B(n_284), .Y(n_318) );
BUFx2_ASAP7_75t_SL g319 ( .A(n_301), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_301), .Y(n_320) );
AO21x2_ASAP7_75t_L g321 ( .A1(n_288), .A2(n_277), .B(n_278), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_289), .A2(n_276), .B1(n_267), .B2(n_271), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_298), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_297), .Y(n_325) );
AO21x1_ASAP7_75t_SL g326 ( .A1(n_299), .A2(n_271), .B(n_274), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_286), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_298), .B(n_274), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_288), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_295), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_290), .B(n_158), .C(n_160), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_300), .B(n_274), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_332), .B(n_320), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_307), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_330), .Y(n_335) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_321), .A2(n_296), .B(n_292), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_330), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_332), .B(n_300), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_332), .B(n_274), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_307), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_320), .B(n_286), .Y(n_342) );
OR2x6_ASAP7_75t_L g343 ( .A(n_319), .B(n_286), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_307), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_307), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_328), .B(n_291), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_309), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_326), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_312), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_312), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_312), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_328), .B(n_291), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_306), .B(n_274), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_286), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_328), .B(n_306), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_313), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_328), .B(n_274), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_313), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_308), .B(n_286), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_308), .B(n_292), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_315), .B(n_292), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_326), .B(n_292), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_315), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_326), .B(n_295), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_315), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_327), .B(n_295), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_333), .B(n_319), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_361), .B(n_327), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_361), .B(n_327), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_360), .B(n_327), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_333), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_354), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_354), .B(n_329), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_334), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_360), .B(n_327), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_363), .B(n_316), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_316), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_366), .B(n_316), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_366), .B(n_323), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_348), .B(n_323), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_367), .B(n_325), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_348), .B(n_325), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_358), .B(n_321), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_367), .B(n_321), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_373), .B(n_329), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_339), .B(n_322), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_339), .B(n_322), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_340), .B(n_305), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_346), .B(n_321), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_346), .B(n_321), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_365), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_346), .B(n_329), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_334), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_341), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_346), .B(n_329), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_350), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_334), .B(n_310), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_334), .B(n_310), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_351), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_365), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_351), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_356), .B(n_310), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_340), .B(n_318), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_355), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_373), .B(n_324), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_356), .B(n_310), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_355), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_358), .B(n_318), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_356), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_359), .B(n_324), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_362), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_341), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_359), .B(n_324), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_362), .B(n_310), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_368), .B(n_310), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_368), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_372), .B(n_331), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_372), .B(n_331), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_374), .B(n_317), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_374), .B(n_317), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_370), .B(n_296), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_341), .Y(n_438) );
INVx4_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_370), .B(n_293), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_344), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_419), .B(n_344), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_439), .B(n_343), .Y(n_443) );
NOR2xp67_ASAP7_75t_L g444 ( .A(n_439), .B(n_385), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_387), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_383), .B(n_343), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_381), .B(n_342), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_410), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_380), .B(n_344), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_377), .B(n_342), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_383), .B(n_343), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_380), .B(n_352), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_377), .B(n_343), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_382), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_402), .A2(n_343), .B(n_375), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_382), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_386), .B(n_352), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_394), .B(n_396), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_386), .B(n_352), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_393), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_378), .B(n_375), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_393), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_424), .B(n_371), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_398), .B(n_353), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_384), .B(n_375), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_428), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_394), .B(n_353), .Y(n_470) );
INVx2_ASAP7_75t_SL g471 ( .A(n_376), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_378), .B(n_353), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_396), .B(n_357), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_379), .B(n_357), .Y(n_474) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_439), .B(n_369), .Y(n_475) );
AND3x2_ASAP7_75t_L g476 ( .A(n_384), .B(n_364), .C(n_357), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_426), .B(n_364), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_427), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_379), .B(n_364), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_405), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_405), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_388), .B(n_335), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_412), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_426), .B(n_335), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_376), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_388), .B(n_335), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_404), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_429), .B(n_337), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_391), .B(n_337), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_384), .B(n_369), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_391), .B(n_337), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_412), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_389), .B(n_338), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_429), .B(n_392), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_438), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_392), .B(n_338), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_395), .B(n_338), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_389), .B(n_369), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_390), .B(n_369), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_398), .B(n_336), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_400), .A2(n_276), .B1(n_371), .B2(n_336), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_390), .B(n_371), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_415), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_415), .B(n_336), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_401), .B(n_371), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_395), .B(n_371), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_421), .B(n_371), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_421), .B(n_336), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_407), .B(n_311), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_417), .B(n_317), .Y(n_512) );
NAND2x1_ASAP7_75t_L g513 ( .A(n_439), .B(n_311), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_417), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_420), .B(n_317), .Y(n_515) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_385), .B(n_311), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_420), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_421), .B(n_311), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_385), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_416), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_421), .B(n_311), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_437), .A2(n_276), .B1(n_261), .B2(n_269), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_385), .B(n_293), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_479), .B(n_430), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_445), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_445), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_503), .B(n_437), .C(n_440), .D(n_397), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_464), .B(n_399), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_496), .B(n_397), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_444), .B(n_409), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g531 ( .A1(n_506), .A2(n_433), .B(n_434), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_489), .Y(n_532) );
O2A1O1Ixp5_ASAP7_75t_L g533 ( .A1(n_513), .A2(n_409), .B(n_384), .C(n_399), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_489), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_451), .B(n_399), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_448), .B(n_399), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_442), .B(n_430), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_442), .B(n_431), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_447), .A2(n_409), .B1(n_425), .B2(n_414), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_460), .B(n_409), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_452), .B(n_413), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_443), .B(n_413), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_455), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_457), .Y(n_544) );
O2A1O1Ixp5_ASAP7_75t_R g545 ( .A1(n_502), .A2(n_437), .B(n_414), .C(n_13), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_500), .B(n_408), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_468), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_463), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_501), .B(n_408), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_520), .B(n_431), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_465), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_468), .B(n_411), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_516), .A2(n_432), .B(n_423), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_498), .B(n_423), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_481), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_454), .B(n_411), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_482), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_520), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_502), .B(n_435), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_499), .B(n_432), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_477), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_443), .B(n_437), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_467), .B(n_441), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_467), .B(n_441), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_495), .B(n_435), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_506), .B(n_436), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_484), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_494), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_505), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_517), .B(n_436), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_486), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_490), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_466), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_446), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_491), .B(n_403), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_450), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_485), .B(n_418), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_446), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_450), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_493), .B(n_403), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_466), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_449), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_453), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_449), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_507), .A2(n_406), .B1(n_418), .B2(n_422), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_485), .B(n_422), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_453), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_497), .B(n_406), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_459), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_459), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_487), .B(n_311), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_458), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_508), .B(n_317), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_461), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_504), .B(n_317), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_461), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_456), .A2(n_158), .B(n_285), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_497), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_526), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_532), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_545), .A2(n_471), .B(n_519), .C(n_511), .Y(n_602) );
OAI321xp33_ASAP7_75t_L g603 ( .A1(n_539), .A2(n_510), .A3(n_522), .B1(n_507), .B2(n_518), .C(n_521), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_540), .A2(n_452), .B1(n_492), .B2(n_443), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_562), .B(n_530), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_534), .B(n_483), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_577), .Y(n_607) );
AOI21xp33_ASAP7_75t_SL g608 ( .A1(n_539), .A2(n_492), .B(n_470), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_525), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_559), .B(n_488), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_547), .B(n_536), .Y(n_611) );
NOR2xp33_ASAP7_75t_SL g612 ( .A(n_530), .B(n_476), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_574), .B(n_473), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_580), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_584), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_533), .A2(n_475), .B(n_523), .Y(n_616) );
AOI211xp5_ASAP7_75t_SL g617 ( .A1(n_598), .A2(n_523), .B(n_509), .C(n_512), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_559), .B(n_474), .Y(n_618) );
OAI32xp33_ASAP7_75t_L g619 ( .A1(n_558), .A2(n_480), .A3(n_472), .B1(n_512), .B2(n_515), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_558), .B(n_523), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_588), .B(n_515), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_531), .A2(n_478), .B(n_458), .C(n_469), .Y(n_622) );
NAND2xp33_ASAP7_75t_SL g623 ( .A(n_541), .B(n_476), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_527), .A2(n_478), .B(n_469), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_561), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_590), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_527), .A2(n_462), .B1(n_295), .B2(n_294), .Y(n_627) );
OAI322xp33_ASAP7_75t_L g628 ( .A1(n_529), .A2(n_462), .A3(n_11), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_16), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_591), .B(n_8), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_553), .A2(n_269), .B1(n_261), .B2(n_265), .C1(n_268), .C2(n_18), .Y(n_630) );
OAI22xp5_ASAP7_75t_SL g631 ( .A1(n_542), .A2(n_295), .B1(n_269), .B2(n_261), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_595), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_597), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_550), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_571), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_531), .A2(n_8), .B(n_15), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_575), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_535), .B(n_287), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_566), .B(n_16), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_566), .B(n_17), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_553), .B(n_269), .C(n_265), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_528), .B(n_287), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_571), .B(n_17), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_542), .A2(n_268), .B1(n_19), .B2(n_20), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_552), .B(n_287), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_582), .A2(n_586), .B1(n_562), .B2(n_594), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_524), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_543), .Y(n_648) );
AOI221x1_ASAP7_75t_L g649 ( .A1(n_572), .A2(n_268), .B1(n_19), .B2(n_18), .C(n_193), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_623), .A2(n_596), .B1(n_573), .B2(n_537), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_608), .A2(n_592), .B(n_578), .Y(n_651) );
NOR2xp33_ASAP7_75t_SL g652 ( .A(n_612), .B(n_563), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_635), .B(n_544), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_607), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_625), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_603), .A2(n_538), .B1(n_555), .B2(n_557), .C(n_568), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_625), .B(n_589), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_630), .A2(n_578), .B(n_587), .C(n_589), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_646), .A2(n_587), .B1(n_556), .B2(n_567), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_612), .A2(n_565), .B1(n_560), .B2(n_554), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_613), .A2(n_569), .B1(n_548), .B2(n_570), .Y(n_661) );
OAI222xp33_ASAP7_75t_L g662 ( .A1(n_604), .A2(n_581), .B1(n_576), .B2(n_564), .C1(n_546), .C2(n_549), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_603), .A2(n_599), .B(n_551), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_634), .A2(n_593), .B1(n_585), .B2(n_583), .Y(n_664) );
BUFx3_ASAP7_75t_L g665 ( .A(n_605), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_602), .A2(n_579), .B(n_193), .C(n_174), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_605), .B(n_21), .Y(n_667) );
INVx2_ASAP7_75t_SL g668 ( .A(n_611), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_619), .A2(n_193), .B1(n_174), .B2(n_27), .C(n_28), .Y(n_669) );
XNOR2x1_ASAP7_75t_L g670 ( .A(n_639), .B(n_25), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_614), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_641), .A2(n_26), .B1(n_29), .B2(n_30), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_624), .A2(n_193), .B1(n_174), .B2(n_36), .C(n_38), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_615), .B(n_33), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_616), .A2(n_34), .B(n_40), .C(n_44), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_640), .A2(n_174), .B1(n_46), .B2(n_47), .C1(n_49), .C2(n_50), .Y(n_676) );
NOR4xp25_ASAP7_75t_L g677 ( .A(n_628), .B(n_45), .C(n_57), .D(n_58), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_617), .A2(n_59), .B(n_60), .C(n_62), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_631), .A2(n_174), .B1(n_65), .B2(n_66), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_647), .B(n_64), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_637), .Y(n_681) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_643), .A2(n_174), .B1(n_68), .B2(n_69), .C1(n_72), .C2(n_73), .Y(n_682) );
AOI221x1_ASAP7_75t_L g683 ( .A1(n_629), .A2(n_67), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_683) );
NAND3xp33_ASAP7_75t_SL g684 ( .A(n_622), .B(n_104), .C(n_79), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_627), .A2(n_77), .B(n_80), .Y(n_685) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_644), .B(n_82), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_636), .A2(n_83), .B(n_85), .C(n_87), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_626), .A2(n_89), .B1(n_94), .B2(n_95), .C(n_96), .Y(n_688) );
NOR3xp33_ASAP7_75t_SL g689 ( .A(n_600), .B(n_97), .C(n_601), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_610), .A2(n_618), .A3(n_642), .B1(n_638), .B2(n_645), .C1(n_606), .C2(n_632), .Y(n_690) );
AOI211xp5_ASAP7_75t_SL g691 ( .A1(n_609), .A2(n_633), .B(n_621), .C(n_648), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_666), .B(n_656), .C(n_691), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_655), .Y(n_693) );
NOR4xp25_ASAP7_75t_L g694 ( .A(n_662), .B(n_651), .C(n_650), .D(n_658), .Y(n_694) );
NAND4xp25_ASAP7_75t_SL g695 ( .A(n_690), .B(n_659), .C(n_663), .D(n_678), .Y(n_695) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_684), .B(n_686), .Y(n_696) );
NAND4xp25_ASAP7_75t_SL g697 ( .A(n_669), .B(n_675), .C(n_682), .D(n_676), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_660), .A2(n_677), .B1(n_652), .B2(n_664), .C(n_671), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_695), .B(n_687), .C(n_688), .Y(n_699) );
NAND4xp75_ASAP7_75t_L g700 ( .A(n_696), .B(n_667), .C(n_689), .D(n_683), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_694), .A2(n_670), .B(n_672), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_692), .B(n_688), .C(n_680), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_702), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_699), .B(n_698), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_701), .A2(n_693), .B1(n_665), .B2(n_668), .Y(n_705) );
OAI22x1_ASAP7_75t_L g706 ( .A1(n_704), .A2(n_697), .B1(n_700), .B2(n_661), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_703), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_705), .B1(n_657), .B2(n_654), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_706), .A2(n_653), .B1(n_681), .B2(n_673), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_708), .Y(n_710) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_709), .A2(n_672), .B1(n_679), .B2(n_674), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_710), .B(n_653), .Y(n_712) );
AOI21xp33_ASAP7_75t_SL g713 ( .A1(n_712), .A2(n_711), .B(n_674), .Y(n_713) );
OR2x6_ASAP7_75t_L g714 ( .A(n_713), .B(n_685), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_620), .B1(n_649), .B2(n_695), .Y(n_715) );
endmodule