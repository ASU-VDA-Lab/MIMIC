module fake_jpeg_6780_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_18),
.B1(n_13),
.B2(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_37),
.B1(n_23),
.B2(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_35),
.B1(n_10),
.B2(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_29),
.B1(n_36),
.B2(n_10),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_52),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_28),
.B1(n_21),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_46),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_56),
.B(n_45),
.C(n_54),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_66),
.B1(n_44),
.B2(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_55),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_57),
.A3(n_22),
.B1(n_41),
.B2(n_52),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_67),
.B(n_66),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_77),
.C(n_58),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_30),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_85),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_58),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_66),
.B(n_58),
.C(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_43),
.B1(n_39),
.B2(n_24),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_77),
.C(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_88),
.C(n_91),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_81),
.B(n_83),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_2),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_83),
.B(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_86),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_91),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_87),
.C(n_88),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_100),
.C(n_2),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_9),
.B(n_7),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.C(n_8),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_7),
.C(n_8),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_99),
.Y(n_109)
);


endmodule