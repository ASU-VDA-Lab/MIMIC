module real_jpeg_33144_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_57;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_58;
wire n_10;
wire n_31;
wire n_9;
wire n_49;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_56;
wire n_20;
wire n_48;
wire n_19;
wire n_32;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_2),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

AOI221xp5_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.C(n_58),
.Y(n_44)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx2_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2x1p5_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_15),
.Y(n_57)
);

AND2x4_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_4),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_7),
.B1(n_14),
.B2(n_15),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_31),
.Y(n_56)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_18),
.B1(n_36),
.B2(n_38),
.C(n_44),
.Y(n_8)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_37),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

OA21x2_ASAP7_75t_L g55 ( 
.A1(n_14),
.A2(n_56),
.B(n_57),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_24),
.B(n_32),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_23),
.B(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_30),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);


endmodule