module real_jpeg_12394_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_286;
wire n_215;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_3),
.B(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_3),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_3),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_3),
.B(n_49),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_52),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_5),
.B(n_43),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_49),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_5),
.B(n_62),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_7),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_7),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_7),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_7),
.B(n_60),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_7),
.B(n_29),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_8),
.B(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_8),
.B(n_29),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_8),
.B(n_49),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_8),
.B(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_8),
.B(n_52),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_31),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_29),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_9),
.B(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_9),
.B(n_49),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_43),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_10),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_10),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_10),
.B(n_31),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_10),
.B(n_60),
.Y(n_233)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_13),
.B(n_43),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_13),
.B(n_49),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_13),
.B(n_62),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_13),
.B(n_31),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_13),
.B(n_60),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_14),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_14),
.B(n_62),
.Y(n_129)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_157),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_156),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_20),
.B(n_121),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.C(n_99),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_21),
.B(n_84),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_54),
.C(n_71),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_46),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_23),
.B(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_28),
.C(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_28),
.B(n_153),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_28),
.A2(n_34),
.B1(n_152),
.B2(n_153),
.Y(n_234)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_32),
.B(n_45),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_32),
.B(n_66),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_36),
.A2(n_37),
.B1(n_46),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_37),
.A2(n_38),
.B(n_41),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_39),
.B(n_111),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_39),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_45),
.B(n_110),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_46),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.C(n_51),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_47),
.B(n_48),
.CI(n_51),
.CON(n_102),
.SN(n_102)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_71),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.C(n_69),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.C(n_64),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_59),
.B(n_66),
.Y(n_251)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_61),
.Y(n_171)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_64),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_75),
.C(n_77),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_75),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_78),
.B(n_81),
.C(n_82),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_80),
.A2(n_81),
.B1(n_104),
.B2(n_105),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_82),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_82),
.A2(n_83),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_82),
.B(n_221),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_93),
.C(n_98),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_89),
.C(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_97),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_113),
.C(n_116),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_100),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.C(n_106),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_101),
.A2(n_102),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_102),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_103),
.B(n_106),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_109),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_155),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_145),
.B2(n_146),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_135),
.B2(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_206),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_182),
.B(n_205),
.Y(n_159)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_160),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_180),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_168),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_165),
.B1(n_168),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_179),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_172),
.CI(n_179),
.CON(n_188),
.SN(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_173),
.A2(n_174),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_183),
.B(n_186),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_193),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_187),
.A2(n_188),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_188),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_285)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_195),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_198),
.B(n_199),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_287),
.C(n_288),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_281),
.B(n_286),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_266),
.B(n_280),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_236),
.B(n_265),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_223),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_211),
.B(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.C(n_220),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_262),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.CI(n_215),
.CON(n_212),
.SN(n_212)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_230),
.B2(n_235),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_229),
.C(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_233),
.C(n_234),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_259),
.B(n_264),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_249),
.B(n_258),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_244),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_247),
.C(n_248),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_253),
.B(n_257),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_261),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_268),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_274),
.C(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_278),
.B2(n_279),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);


endmodule