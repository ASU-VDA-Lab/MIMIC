module real_aes_10572_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1632;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1584;
wire n_1277;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_0), .A2(n_148), .B1(n_515), .B2(n_868), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_0), .A2(n_148), .B1(n_453), .B2(n_677), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_1), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_1), .A2(n_9), .B1(n_462), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_2), .A2(n_78), .B1(n_688), .B2(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g882 ( .A(n_2), .Y(n_882) );
INVx1_ASAP7_75t_L g1108 ( .A(n_3), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_4), .A2(n_210), .B1(n_543), .B2(n_544), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_4), .A2(n_210), .B1(n_495), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_5), .A2(n_17), .B1(n_491), .B2(n_913), .Y(n_912) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_5), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_6), .A2(n_160), .B1(n_479), .B2(n_562), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_6), .A2(n_160), .B1(n_651), .B2(n_657), .Y(n_1272) );
INVx1_ASAP7_75t_L g512 ( .A(n_7), .Y(n_512) );
INVx1_ASAP7_75t_L g852 ( .A(n_8), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_8), .A2(n_234), .B1(n_552), .B2(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g523 ( .A(n_9), .Y(n_523) );
INVxp33_ASAP7_75t_SL g902 ( .A(n_10), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_10), .A2(n_284), .B1(n_924), .B2(n_926), .Y(n_923) );
INVxp33_ASAP7_75t_SL g398 ( .A(n_11), .Y(n_398) );
AOI22xp5_ASAP7_75t_SL g490 ( .A1(n_11), .A2(n_257), .B1(n_491), .B2(n_495), .Y(n_490) );
INVx1_ASAP7_75t_L g801 ( .A(n_12), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_12), .A2(n_65), .B1(n_530), .B2(n_816), .Y(n_815) );
AO22x1_ASAP7_75t_L g339 ( .A1(n_13), .A2(n_340), .B1(n_341), .B2(n_503), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_13), .Y(n_340) );
AOI22xp33_ASAP7_75t_SL g1168 ( .A1(n_14), .A2(n_267), .B1(n_479), .B2(n_1169), .Y(n_1168) );
INVxp67_ASAP7_75t_L g1178 ( .A(n_14), .Y(n_1178) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_15), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_15), .A2(n_202), .B1(n_533), .B2(n_834), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_16), .A2(n_207), .B1(n_447), .B2(n_451), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_16), .A2(n_207), .B1(n_484), .B2(n_487), .Y(n_483) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_17), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_18), .A2(n_198), .B1(n_738), .B2(n_739), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_18), .A2(n_198), .B1(n_749), .B2(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g511 ( .A(n_19), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_19), .A2(n_60), .B1(n_530), .B2(n_546), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g1535 ( .A1(n_20), .A2(n_246), .B1(n_977), .B2(n_1536), .C(n_1538), .Y(n_1535) );
INVx1_ASAP7_75t_L g1599 ( .A(n_20), .Y(n_1599) );
INVx1_ASAP7_75t_L g726 ( .A(n_21), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_21), .A2(n_220), .B1(n_532), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_22), .A2(n_306), .B1(n_515), .B2(n_868), .Y(n_872) );
INVx1_ASAP7_75t_L g878 ( .A(n_22), .Y(n_878) );
XOR2x2_ASAP7_75t_L g889 ( .A(n_23), .B(n_890), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_23), .A2(n_116), .B1(n_1284), .B2(n_1292), .Y(n_1283) );
INVx1_ASAP7_75t_L g595 ( .A(n_24), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_25), .A2(n_73), .B1(n_455), .B2(n_1217), .Y(n_1216) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_25), .A2(n_73), .B1(n_1228), .B2(n_1229), .Y(n_1227) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_26), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_26), .A2(n_197), .B1(n_491), .B2(n_919), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_27), .A2(n_231), .B1(n_543), .B2(n_544), .Y(n_811) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_27), .A2(n_231), .B1(n_684), .B2(n_688), .Y(n_819) );
OAI211xp5_ASAP7_75t_L g1055 ( .A1(n_28), .A2(n_648), .B(n_1056), .C(n_1059), .Y(n_1055) );
INVx1_ASAP7_75t_L g1077 ( .A(n_28), .Y(n_1077) );
INVx1_ASAP7_75t_L g1200 ( .A(n_29), .Y(n_1200) );
INVx1_ASAP7_75t_L g1155 ( .A(n_30), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_30), .A2(n_33), .B1(n_532), .B2(n_768), .Y(n_1175) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_31), .A2(n_84), .B1(n_738), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_31), .A2(n_84), .B1(n_919), .B2(n_1042), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g1087 ( .A(n_32), .Y(n_1087) );
INVx1_ASAP7_75t_L g1156 ( .A(n_33), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1525 ( .A1(n_34), .A2(n_309), .B1(n_1526), .B2(n_1532), .Y(n_1525) );
INVx1_ASAP7_75t_L g1581 ( .A(n_34), .Y(n_1581) );
INVx1_ASAP7_75t_L g586 ( .A(n_35), .Y(n_586) );
INVx1_ASAP7_75t_L g787 ( .A(n_36), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_36), .A2(n_146), .B1(n_479), .B2(n_570), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_37), .A2(n_301), .B1(n_760), .B2(n_761), .Y(n_759) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_37), .Y(n_771) );
INVx1_ASAP7_75t_L g317 ( .A(n_38), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_39), .A2(n_108), .B1(n_1284), .B2(n_1292), .Y(n_1302) );
AOI221xp5_ASAP7_75t_L g1250 ( .A1(n_40), .A2(n_214), .B1(n_738), .B2(n_742), .C(n_1251), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_40), .A2(n_214), .B1(n_479), .B2(n_570), .Y(n_1262) );
INVx1_ASAP7_75t_L g1333 ( .A(n_41), .Y(n_1333) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_42), .A2(n_58), .B1(n_326), .B2(n_433), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_42), .A2(n_297), .B1(n_636), .B2(n_640), .Y(n_711) );
INVx1_ASAP7_75t_L g1547 ( .A(n_43), .Y(n_1547) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_43), .A2(n_282), .B1(n_734), .B2(n_879), .Y(n_1588) );
INVx1_ASAP7_75t_L g377 ( .A(n_44), .Y(n_377) );
INVx1_ASAP7_75t_L g1158 ( .A(n_45), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1622 ( .A(n_46), .Y(n_1622) );
AOI22xp33_ASAP7_75t_L g1638 ( .A1(n_46), .A2(n_173), .B1(n_552), .B2(n_1127), .Y(n_1638) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_47), .A2(n_170), .B1(n_465), .B2(n_734), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_47), .A2(n_170), .B1(n_374), .B2(n_753), .Y(n_752) );
INVxp33_ASAP7_75t_L g1020 ( .A(n_48), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_48), .A2(n_258), .B1(n_568), .B2(n_644), .Y(n_1045) );
INVxp33_ASAP7_75t_SL g430 ( .A(n_49), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_49), .A2(n_255), .B1(n_484), .B2(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_50), .A2(n_274), .B1(n_543), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_50), .A2(n_274), .B1(n_683), .B2(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g1563 ( .A(n_51), .Y(n_1563) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_51), .A2(n_286), .B1(n_972), .B2(n_1587), .Y(n_1586) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_52), .A2(n_71), .B1(n_1296), .B2(n_1300), .Y(n_1295) );
INVxp33_ASAP7_75t_SL g1109 ( .A(n_53), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_53), .A2(n_177), .B1(n_552), .B2(n_1127), .Y(n_1126) );
INVxp33_ASAP7_75t_SL g1123 ( .A(n_54), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_54), .A2(n_68), .B1(n_758), .B2(n_1140), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1626 ( .A1(n_55), .A2(n_76), .B1(n_651), .B2(n_657), .Y(n_1626) );
AOI22xp33_ASAP7_75t_L g1647 ( .A1(n_55), .A2(n_76), .B1(n_683), .B2(n_751), .Y(n_1647) );
INVxp67_ASAP7_75t_SL g1196 ( .A(n_56), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_56), .A2(n_67), .B1(n_570), .B2(n_1234), .Y(n_1233) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_57), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_57), .A2(n_194), .B1(n_742), .B2(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_58), .A2(n_165), .B1(n_690), .B2(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g1264 ( .A(n_59), .Y(n_1264) );
INVx1_ASAP7_75t_L g516 ( .A(n_60), .Y(n_516) );
INVx1_ASAP7_75t_L g528 ( .A(n_61), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_61), .A2(n_226), .B1(n_489), .B2(n_568), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g1243 ( .A1(n_62), .A2(n_648), .B(n_1244), .C(n_1245), .Y(n_1243) );
INVx1_ASAP7_75t_L g1258 ( .A(n_62), .Y(n_1258) );
INVx1_ASAP7_75t_L g790 ( .A(n_63), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_63), .A2(n_162), .B1(n_559), .B2(n_822), .Y(n_821) );
OAI211xp5_ASAP7_75t_L g829 ( .A1(n_63), .A2(n_434), .B(n_830), .C(n_832), .Y(n_829) );
XNOR2xp5_ASAP7_75t_L g844 ( .A(n_64), .B(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1319 ( .A1(n_64), .A2(n_182), .B1(n_1284), .B2(n_1292), .Y(n_1319) );
INVx1_ASAP7_75t_L g805 ( .A(n_65), .Y(n_805) );
OAI211xp5_ASAP7_75t_L g838 ( .A1(n_65), .A2(n_648), .B(n_839), .C(n_841), .Y(n_838) );
AO22x1_ASAP7_75t_SL g1358 ( .A1(n_66), .A2(n_117), .B1(n_1284), .B2(n_1292), .Y(n_1358) );
INVxp67_ASAP7_75t_SL g1203 ( .A(n_67), .Y(n_1203) );
INVxp67_ASAP7_75t_SL g1117 ( .A(n_68), .Y(n_1117) );
INVx1_ASAP7_75t_L g583 ( .A(n_69), .Y(n_583) );
INVx1_ASAP7_75t_L g802 ( .A(n_70), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_70), .A2(n_290), .B1(n_458), .B2(n_552), .Y(n_814) );
INVx1_ASAP7_75t_L g699 ( .A(n_72), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_74), .A2(n_196), .B1(n_1300), .B2(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g373 ( .A(n_75), .Y(n_373) );
AOI22xp33_ASAP7_75t_SL g464 ( .A1(n_75), .A2(n_112), .B1(n_447), .B2(n_465), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_77), .A2(n_235), .B1(n_1081), .B2(n_1082), .C(n_1084), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_77), .A2(n_235), .B1(n_570), .B2(n_604), .Y(n_1094) );
INVx1_ASAP7_75t_L g884 ( .A(n_78), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_79), .A2(n_90), .B1(n_1135), .B2(n_1137), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_79), .A2(n_90), .B1(n_758), .B2(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g363 ( .A(n_80), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_81), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g1324 ( .A1(n_82), .A2(n_103), .B1(n_1300), .B2(n_1321), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_83), .A2(n_222), .B1(n_651), .B2(n_657), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_83), .A2(n_222), .B1(n_562), .B2(n_604), .Y(n_1098) );
BUFx2_ASAP7_75t_L g395 ( .A(n_85), .Y(n_395) );
BUFx2_ASAP7_75t_L g439 ( .A(n_85), .Y(n_439) );
INVx1_ASAP7_75t_L g469 ( .A(n_85), .Y(n_469) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_85), .B(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g724 ( .A(n_86), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_86), .A2(n_174), .B1(n_734), .B2(n_744), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_87), .A2(n_224), .B1(n_907), .B2(n_910), .Y(n_906) );
INVxp67_ASAP7_75t_SL g941 ( .A(n_87), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_88), .A2(n_300), .B1(n_919), .B2(n_920), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_88), .A2(n_300), .B1(n_924), .B2(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g1111 ( .A(n_89), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_89), .A2(n_107), .B1(n_546), .B2(n_671), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_91), .A2(n_287), .B1(n_670), .B2(n_671), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_91), .A2(n_287), .B1(n_515), .B2(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g1335 ( .A(n_92), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_93), .A2(n_252), .B1(n_910), .B2(n_917), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_93), .A2(n_252), .B1(n_879), .B2(n_936), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_94), .A2(n_250), .B1(n_552), .B2(n_1131), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_94), .A2(n_250), .B1(n_482), .B2(n_1142), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_95), .A2(n_266), .B1(n_1284), .B2(n_1292), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_96), .A2(n_276), .B1(n_671), .B2(n_734), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_96), .A2(n_276), .B1(n_691), .B2(n_756), .Y(n_1226) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_97), .Y(n_1068) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_98), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g1167 ( .A1(n_99), .A2(n_304), .B1(n_680), .B2(n_691), .Y(n_1167) );
INVxp33_ASAP7_75t_L g1180 ( .A(n_99), .Y(n_1180) );
OAI22xp33_ASAP7_75t_L g1248 ( .A1(n_100), .A2(n_223), .B1(n_638), .B2(n_641), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_100), .A2(n_223), .B1(n_455), .B2(n_1222), .C(n_1256), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_101), .A2(n_238), .B1(n_1296), .B2(n_1300), .Y(n_1303) );
INVx1_ASAP7_75t_L g646 ( .A(n_102), .Y(n_646) );
INVx1_ASAP7_75t_L g384 ( .A(n_104), .Y(n_384) );
INVx1_ASAP7_75t_L g712 ( .A(n_105), .Y(n_712) );
INVx1_ASAP7_75t_L g1252 ( .A(n_106), .Y(n_1252) );
INVxp33_ASAP7_75t_SL g1105 ( .A(n_107), .Y(n_1105) );
INVx1_ASAP7_75t_L g633 ( .A(n_109), .Y(n_633) );
INVx1_ASAP7_75t_L g1361 ( .A(n_110), .Y(n_1361) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_111), .A2(n_139), .B1(n_548), .B2(n_677), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_111), .A2(n_139), .B1(n_489), .B2(n_568), .Y(n_818) );
INVxp33_ASAP7_75t_SL g344 ( .A(n_112), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_113), .Y(n_1085) );
INVx1_ASAP7_75t_L g600 ( .A(n_114), .Y(n_600) );
OAI22xp33_ASAP7_75t_SL g656 ( .A1(n_114), .A2(n_199), .B1(n_326), .B2(n_657), .Y(n_656) );
AO22x2_ASAP7_75t_L g1147 ( .A1(n_115), .A2(n_1148), .B1(n_1181), .B2(n_1182), .Y(n_1147) );
INVx1_ASAP7_75t_L g1181 ( .A(n_115), .Y(n_1181) );
INVx1_ASAP7_75t_L g1247 ( .A(n_118), .Y(n_1247) );
INVxp33_ASAP7_75t_SL g1017 ( .A(n_119), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_119), .A2(n_200), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_120), .A2(n_228), .B1(n_756), .B2(n_910), .Y(n_981) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_120), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_121), .A2(n_272), .B1(n_570), .B2(n_604), .Y(n_1162) );
AOI22xp33_ASAP7_75t_SL g1170 ( .A1(n_121), .A2(n_272), .B1(n_543), .B2(n_544), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g1548 ( .A1(n_122), .A2(n_279), .B1(n_1549), .B2(n_1551), .C(n_1553), .Y(n_1548) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_122), .A2(n_188), .B1(n_926), .B2(n_972), .Y(n_1585) );
INVx1_ASAP7_75t_L g851 ( .A(n_123), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_123), .A2(n_237), .B1(n_671), .B2(n_816), .Y(n_865) );
INVx1_ASAP7_75t_L g961 ( .A(n_124), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_124), .A2(n_268), .B1(n_532), .B2(n_768), .Y(n_988) );
INVxp33_ASAP7_75t_L g1206 ( .A(n_125), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_125), .A2(n_167), .B1(n_451), .B2(n_734), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_126), .A2(n_262), .B1(n_1028), .B2(n_1030), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_126), .A2(n_262), .B1(n_644), .B2(n_907), .Y(n_1040) );
INVxp33_ASAP7_75t_SL g1004 ( .A(n_127), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_127), .A2(n_296), .B1(n_1033), .B2(n_1035), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_128), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_128), .A2(n_193), .B1(n_453), .B2(n_670), .Y(n_1165) );
INVx1_ASAP7_75t_L g626 ( .A(n_129), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_129), .A2(n_131), .B1(n_636), .B2(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g1195 ( .A(n_130), .Y(n_1195) );
INVx1_ASAP7_75t_L g630 ( .A(n_131), .Y(n_630) );
INVxp33_ASAP7_75t_SL g1152 ( .A(n_132), .Y(n_1152) );
AOI22xp33_ASAP7_75t_SL g1164 ( .A1(n_132), .A2(n_281), .B1(n_543), .B2(n_544), .Y(n_1164) );
INVx1_ASAP7_75t_L g1288 ( .A(n_133), .Y(n_1288) );
OAI211xp5_ASAP7_75t_L g1627 ( .A1(n_134), .A2(n_434), .B(n_653), .C(n_1628), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g1646 ( .A1(n_134), .A2(n_233), .B1(n_868), .B2(n_1642), .Y(n_1646) );
INVxp33_ASAP7_75t_SL g953 ( .A(n_135), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_135), .A2(n_171), .B1(n_734), .B2(n_744), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_136), .A2(n_221), .B1(n_546), .B2(n_548), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_136), .A2(n_221), .B1(n_558), .B2(n_559), .Y(n_557) );
XOR2x2_ASAP7_75t_L g713 ( .A(n_137), .B(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_138), .A2(n_208), .B1(n_1633), .B2(n_1634), .Y(n_1632) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_138), .A2(n_208), .B1(n_683), .B2(n_751), .Y(n_1644) );
CKINVDCx20_ASAP7_75t_R g1198 ( .A(n_140), .Y(n_1198) );
INVx1_ASAP7_75t_L g1010 ( .A(n_141), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_141), .A2(n_254), .B1(n_768), .B2(n_793), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1329 ( .A1(n_142), .A2(n_216), .B1(n_1330), .B2(n_1331), .C(n_1332), .Y(n_1329) );
AO22x2_ASAP7_75t_SL g948 ( .A1(n_143), .A2(n_949), .B1(n_950), .B2(n_994), .Y(n_948) );
CKINVDCx16_ASAP7_75t_R g949 ( .A(n_143), .Y(n_949) );
INVxp33_ASAP7_75t_SL g893 ( .A(n_144), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_144), .A2(n_156), .B1(n_735), .B2(n_879), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_145), .A2(n_260), .B1(n_455), .B2(n_458), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_145), .A2(n_260), .B1(n_478), .B2(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g788 ( .A(n_146), .Y(n_788) );
INVx1_ASAP7_75t_L g1289 ( .A(n_147), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_147), .B(n_1287), .Y(n_1294) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_149), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_150), .A2(n_204), .B1(n_453), .B2(n_677), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_150), .A2(n_204), .B1(n_515), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1554 ( .A1(n_151), .A2(n_188), .B1(n_484), .B2(n_1555), .Y(n_1554) );
AOI22xp33_ASAP7_75t_SL g1584 ( .A1(n_151), .A2(n_279), .B1(n_415), .B2(n_448), .Y(n_1584) );
INVxp33_ASAP7_75t_SL g356 ( .A(n_152), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_152), .A2(n_217), .B1(n_455), .B2(n_462), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_153), .A2(n_163), .B1(n_636), .B2(n_638), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1072 ( .A1(n_153), .A2(n_269), .B1(n_455), .B2(n_969), .C(n_1073), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1540 ( .A1(n_154), .A2(n_757), .B(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1597 ( .A(n_154), .Y(n_1597) );
INVx2_ASAP7_75t_L g329 ( .A(n_155), .Y(n_329) );
INVxp67_ASAP7_75t_SL g896 ( .A(n_156), .Y(n_896) );
AO221x2_ASAP7_75t_L g1306 ( .A1(n_157), .A2(n_186), .B1(n_1296), .B2(n_1307), .C(n_1309), .Y(n_1306) );
INVxp33_ASAP7_75t_L g1003 ( .A(n_158), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_158), .A2(n_292), .B1(n_453), .B2(n_1038), .Y(n_1037) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_159), .A2(n_271), .B1(n_756), .B2(n_758), .Y(n_755) );
INVxp33_ASAP7_75t_SL g773 ( .A(n_159), .Y(n_773) );
BUFx3_ASAP7_75t_L g353 ( .A(n_161), .Y(n_353) );
INVx1_ASAP7_75t_L g371 ( .A(n_161), .Y(n_371) );
INVx1_ASAP7_75t_L g797 ( .A(n_162), .Y(n_797) );
INVx1_ASAP7_75t_L g1074 ( .A(n_163), .Y(n_1074) );
INVxp33_ASAP7_75t_L g1202 ( .A(n_164), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_164), .A2(n_219), .B1(n_756), .B2(n_1237), .Y(n_1236) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_165), .A2(n_434), .B(n_695), .C(n_698), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_166), .A2(n_211), .B1(n_455), .B2(n_969), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_166), .A2(n_211), .B1(n_976), .B2(n_977), .Y(n_975) );
INVx1_ASAP7_75t_L g1211 ( .A(n_167), .Y(n_1211) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_168), .A2(n_305), .B1(n_465), .B2(n_734), .Y(n_967) );
AOI22xp33_ASAP7_75t_SL g979 ( .A1(n_168), .A2(n_305), .B1(n_758), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_169), .A2(n_297), .B1(n_671), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g705 ( .A(n_169), .Y(n_705) );
INVx1_ASAP7_75t_L g959 ( .A(n_171), .Y(n_959) );
INVx1_ASAP7_75t_L g1620 ( .A(n_172), .Y(n_1620) );
INVx1_ASAP7_75t_L g1623 ( .A(n_173), .Y(n_1623) );
INVxp33_ASAP7_75t_SL g717 ( .A(n_174), .Y(n_717) );
XNOR2xp5_ASAP7_75t_L g1050 ( .A(n_175), .B(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g601 ( .A(n_176), .Y(n_601) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_176), .A2(n_434), .B(n_653), .C(n_655), .Y(n_652) );
INVxp33_ASAP7_75t_SL g1106 ( .A(n_177), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_178), .A2(n_256), .B1(n_636), .B2(n_640), .Y(n_1242) );
INVx1_ASAP7_75t_L g1271 ( .A(n_178), .Y(n_1271) );
INVx1_ASAP7_75t_L g393 ( .A(n_179), .Y(n_393) );
INVx1_ASAP7_75t_L g1524 ( .A(n_179), .Y(n_1524) );
INVx1_ASAP7_75t_L g700 ( .A(n_180), .Y(n_700) );
INVxp67_ASAP7_75t_L g538 ( .A(n_181), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_181), .A2(n_259), .B1(n_479), .B2(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g857 ( .A(n_183), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g880 ( .A1(n_183), .A2(n_288), .B1(n_768), .B2(n_793), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g1609 ( .A1(n_184), .A2(n_1610), .B1(n_1611), .B2(n_1612), .Y(n_1609) );
CKINVDCx5p33_ASAP7_75t_R g1610 ( .A(n_184), .Y(n_1610) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_185), .A2(n_302), .B1(n_543), .B2(n_544), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_185), .A2(n_302), .B1(n_482), .B2(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_187), .A2(n_245), .B1(n_1284), .B2(n_1292), .Y(n_1323) );
AOI22xp5_ASAP7_75t_L g1346 ( .A1(n_189), .A2(n_265), .B1(n_1300), .B2(n_1321), .Y(n_1346) );
INVx1_ASAP7_75t_L g1601 ( .A(n_189), .Y(n_1601) );
AOI22xp33_ASAP7_75t_L g1607 ( .A1(n_189), .A2(n_1608), .B1(n_1648), .B2(n_1652), .Y(n_1607) );
CKINVDCx14_ASAP7_75t_R g1239 ( .A(n_190), .Y(n_1239) );
INVx1_ASAP7_75t_L g721 ( .A(n_191), .Y(n_721) );
INVx1_ASAP7_75t_L g1246 ( .A(n_192), .Y(n_1246) );
INVxp33_ASAP7_75t_SL g1151 ( .A(n_193), .Y(n_1151) );
INVxp33_ASAP7_75t_SL g954 ( .A(n_194), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_195), .A2(n_264), .B1(n_482), .B2(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_195), .A2(n_264), .B1(n_651), .B2(n_657), .Y(n_693) );
INVxp33_ASAP7_75t_L g1120 ( .A(n_197), .Y(n_1120) );
INVx1_ASAP7_75t_L g605 ( .A(n_199), .Y(n_605) );
INVxp67_ASAP7_75t_SL g1018 ( .A(n_200), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_201), .A2(n_269), .B1(n_640), .B2(n_641), .Y(n_1054) );
INVx1_ASAP7_75t_L g1069 ( .A(n_201), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g899 ( .A(n_202), .Y(n_899) );
INVx1_ASAP7_75t_L g956 ( .A(n_203), .Y(n_956) );
INVx1_ASAP7_75t_L g901 ( .A(n_205), .Y(n_901) );
INVx1_ASAP7_75t_L g1619 ( .A(n_206), .Y(n_1619) );
INVx1_ASAP7_75t_L g1362 ( .A(n_209), .Y(n_1362) );
CKINVDCx20_ASAP7_75t_R g1310 ( .A(n_212), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1636 ( .A1(n_213), .A2(n_241), .B1(n_671), .B2(n_677), .Y(n_1636) );
AOI22xp33_ASAP7_75t_L g1641 ( .A1(n_213), .A2(n_241), .B1(n_568), .B2(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1254 ( .A(n_215), .Y(n_1254) );
INVxp33_ASAP7_75t_SL g367 ( .A(n_217), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_218), .A2(n_247), .B1(n_543), .B2(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g710 ( .A(n_218), .Y(n_710) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_219), .Y(n_1199) );
INVx1_ASAP7_75t_L g728 ( .A(n_220), .Y(n_728) );
INVxp67_ASAP7_75t_SL g944 ( .A(n_224), .Y(n_944) );
INVx1_ASAP7_75t_L g607 ( .A(n_225), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_225), .A2(n_236), .B1(n_433), .B2(n_651), .Y(n_650) );
INVxp33_ASAP7_75t_L g535 ( .A(n_226), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_227), .Y(n_1065) );
INVxp33_ASAP7_75t_L g993 ( .A(n_228), .Y(n_993) );
BUFx3_ASAP7_75t_L g355 ( .A(n_229), .Y(n_355) );
INVx1_ASAP7_75t_L g361 ( .A(n_229), .Y(n_361) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_230), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_230), .A2(n_240), .B1(n_455), .B2(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g1265 ( .A(n_232), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1629 ( .A1(n_233), .A2(n_289), .B1(n_326), .B2(n_433), .Y(n_1629) );
INVx1_ASAP7_75t_L g849 ( .A(n_234), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_236), .A2(n_242), .B1(n_640), .B2(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g854 ( .A(n_237), .Y(n_854) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_239), .Y(n_325) );
INVx1_ASAP7_75t_L g471 ( .A(n_239), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_239), .B(n_294), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_239), .B(n_402), .Y(n_1594) );
INVxp33_ASAP7_75t_SL g719 ( .A(n_240), .Y(n_719) );
INVx1_ASAP7_75t_L g627 ( .A(n_242), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g577 ( .A(n_243), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g348 ( .A(n_244), .Y(n_348) );
OR2x2_ASAP7_75t_L g1523 ( .A(n_244), .B(n_1524), .Y(n_1523) );
INVx1_ASAP7_75t_L g507 ( .A(n_245), .Y(n_507) );
INVx1_ASAP7_75t_L g1590 ( .A(n_246), .Y(n_1590) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_247), .Y(n_709) );
INVx1_ASAP7_75t_L g1006 ( .A(n_248), .Y(n_1006) );
INVx1_ASAP7_75t_L g1113 ( .A(n_249), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_249), .A2(n_278), .B1(n_532), .B2(n_533), .Y(n_1118) );
INVx1_ASAP7_75t_L g647 ( .A(n_251), .Y(n_647) );
INVx1_ASAP7_75t_L g1565 ( .A(n_253), .Y(n_1565) );
INVx1_ASAP7_75t_L g1011 ( .A(n_254), .Y(n_1011) );
INVx1_ASAP7_75t_L g414 ( .A(n_255), .Y(n_414) );
INVx1_ASAP7_75t_L g1257 ( .A(n_256), .Y(n_1257) );
INVxp33_ASAP7_75t_SL g407 ( .A(n_257), .Y(n_407) );
INVxp67_ASAP7_75t_SL g1014 ( .A(n_258), .Y(n_1014) );
INVx1_ASAP7_75t_L g536 ( .A(n_259), .Y(n_536) );
AO22x2_ASAP7_75t_L g783 ( .A1(n_261), .A2(n_784), .B1(n_825), .B2(n_826), .Y(n_783) );
INVxp67_ASAP7_75t_L g825 ( .A(n_261), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_263), .A2(n_293), .B1(n_518), .B2(n_521), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_263), .A2(n_293), .B1(n_532), .B2(n_533), .Y(n_531) );
INVxp33_ASAP7_75t_L g1177 ( .A(n_267), .Y(n_1177) );
INVx1_ASAP7_75t_L g962 ( .A(n_268), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_270), .Y(n_798) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_271), .Y(n_766) );
INVx1_ASAP7_75t_L g1191 ( .A(n_273), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g1624 ( .A1(n_275), .A2(n_289), .B1(n_636), .B2(n_640), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g1639 ( .A1(n_275), .A2(n_298), .B1(n_816), .B2(n_1137), .Y(n_1639) );
INVx1_ASAP7_75t_L g589 ( .A(n_277), .Y(n_589) );
INVx1_ASAP7_75t_L g1112 ( .A(n_278), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1207 ( .A(n_280), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_280), .A2(n_295), .B1(n_972), .B2(n_1222), .Y(n_1221) );
INVxp33_ASAP7_75t_SL g1159 ( .A(n_281), .Y(n_1159) );
INVx1_ASAP7_75t_L g1560 ( .A(n_282), .Y(n_1560) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_283), .B(n_317), .Y(n_1291) );
AND3x2_ASAP7_75t_L g1299 ( .A(n_283), .B(n_317), .C(n_1288), .Y(n_1299) );
INVxp33_ASAP7_75t_SL g894 ( .A(n_284), .Y(n_894) );
INVx2_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
INVx1_ASAP7_75t_L g1520 ( .A(n_286), .Y(n_1520) );
INVx1_ASAP7_75t_L g855 ( .A(n_288), .Y(n_855) );
INVx1_ASAP7_75t_L g807 ( .A(n_290), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_291), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1009 ( .A(n_292), .Y(n_1009) );
INVx1_ASAP7_75t_L g332 ( .A(n_294), .Y(n_332) );
INVx2_ASAP7_75t_L g402 ( .A(n_294), .Y(n_402) );
INVxp67_ASAP7_75t_SL g1209 ( .A(n_295), .Y(n_1209) );
INVxp33_ASAP7_75t_L g1007 ( .A(n_296), .Y(n_1007) );
INVx1_ASAP7_75t_L g1617 ( .A(n_298), .Y(n_1617) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_299), .Y(n_1061) );
INVxp33_ASAP7_75t_SL g770 ( .A(n_301), .Y(n_770) );
XOR2x2_ASAP7_75t_L g1101 ( .A(n_303), .B(n_1102), .Y(n_1101) );
INVxp67_ASAP7_75t_SL g1174 ( .A(n_304), .Y(n_1174) );
INVx1_ASAP7_75t_L g886 ( .A(n_306), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_307), .A2(n_310), .B1(n_983), .B2(n_984), .Y(n_982) );
INVxp33_ASAP7_75t_L g990 ( .A(n_307), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g1539 ( .A(n_308), .Y(n_1539) );
INVx1_ASAP7_75t_L g1579 ( .A(n_309), .Y(n_1579) );
INVxp67_ASAP7_75t_SL g991 ( .A(n_310), .Y(n_991) );
AO22x1_ASAP7_75t_L g998 ( .A1(n_311), .A2(n_999), .B1(n_1000), .B2(n_1049), .Y(n_998) );
INVxp67_ASAP7_75t_L g999 ( .A(n_311), .Y(n_999) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_333), .B(n_1273), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_320), .Y(n_314) );
AND2x4_ASAP7_75t_L g1606 ( .A(n_315), .B(n_321), .Y(n_1606) );
NOR2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_SL g1651 ( .A(n_316), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_316), .B(n_318), .Y(n_1657) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_318), .B(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x6_ASAP7_75t_L g438 ( .A(n_323), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g539 ( .A(n_323), .B(n_439), .Y(n_539) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g445 ( .A(n_324), .B(n_332), .Y(n_445) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g617 ( .A(n_325), .B(n_401), .Y(n_617) );
INVx8_ASAP7_75t_L g431 ( .A(n_326), .Y(n_431) );
OR2x6_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
OR2x6_ASAP7_75t_L g433 ( .A(n_327), .B(n_400), .Y(n_433) );
INVx2_ASAP7_75t_SL g612 ( .A(n_327), .Y(n_612) );
INVx2_ASAP7_75t_SL g1076 ( .A(n_327), .Y(n_1076) );
BUFx6f_ASAP7_75t_L g1086 ( .A(n_327), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_327), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1568 ( .A(n_327), .B(n_1569), .Y(n_1568) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
AND2x4_ASAP7_75t_L g411 ( .A(n_329), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_329), .Y(n_419) );
INVx1_ASAP7_75t_L g425 ( .A(n_329), .Y(n_425) );
AND2x2_ASAP7_75t_L g450 ( .A(n_329), .B(n_330), .Y(n_450) );
INVx1_ASAP7_75t_L g406 ( .A(n_330), .Y(n_406) );
INVx2_ASAP7_75t_L g412 ( .A(n_330), .Y(n_412) );
INVx1_ASAP7_75t_L g421 ( .A(n_330), .Y(n_421) );
INVx1_ASAP7_75t_L g615 ( .A(n_330), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_330), .B(n_404), .Y(n_621) );
AND2x4_ASAP7_75t_L g420 ( .A(n_331), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g533 ( .A(n_332), .B(n_424), .Y(n_533) );
OR2x2_ASAP7_75t_L g768 ( .A(n_332), .B(n_424), .Y(n_768) );
XNOR2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_777), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_573), .B1(n_574), .B2(n_776), .Y(n_334) );
INVx1_ASAP7_75t_L g776 ( .A(n_335), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_504), .B2(n_572), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g1309 ( .A1(n_340), .A2(n_1310), .B1(n_1311), .B2(n_1313), .Y(n_1309) );
INVx1_ASAP7_75t_L g503 ( .A(n_341), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_391), .B1(n_396), .B2(n_437), .C(n_440), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_362), .C(n_372), .D(n_387), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B1(n_356), .B2(n_357), .Y(n_343) );
AOI22xp5_ASAP7_75t_SL g510 ( .A1(n_345), .A2(n_364), .B1(n_511), .B2(n_512), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_345), .A2(n_357), .B1(n_851), .B2(n_852), .Y(n_850) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_345), .A2(n_357), .B1(n_388), .B2(n_893), .C(n_894), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_345), .A2(n_357), .B1(n_953), .B2(n_954), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_345), .A2(n_357), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_345), .A2(n_357), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_345), .A2(n_357), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
AND2x6_ASAP7_75t_L g368 ( .A(n_346), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g718 ( .A(n_346), .B(n_349), .Y(n_718) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g519 ( .A(n_347), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g359 ( .A(n_348), .Y(n_359) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_348), .Y(n_366) );
AND2x2_ASAP7_75t_L g476 ( .A(n_348), .B(n_393), .Y(n_476) );
INVx2_ASAP7_75t_L g502 ( .A(n_348), .Y(n_502) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g486 ( .A(n_350), .Y(n_486) );
INVx1_ASAP7_75t_L g558 ( .A(n_350), .Y(n_558) );
INVx1_ASAP7_75t_L g690 ( .A(n_350), .Y(n_690) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_350), .Y(n_754) );
INVx2_ASAP7_75t_L g757 ( .A(n_350), .Y(n_757) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_350), .Y(n_823) );
INVx2_ASAP7_75t_SL g909 ( .A(n_350), .Y(n_909) );
INVx6_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g364 ( .A(n_351), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g568 ( .A(n_351), .Y(n_568) );
INVx2_ASAP7_75t_L g681 ( .A(n_351), .Y(n_681) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_351), .B(n_1528), .Y(n_1573) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g386 ( .A(n_352), .Y(n_386) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g360 ( .A(n_353), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g376 ( .A(n_353), .B(n_355), .Y(n_376) );
INVx1_ASAP7_75t_L g383 ( .A(n_354), .Y(n_383) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g370 ( .A(n_355), .B(n_371), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_357), .A2(n_368), .B1(n_523), .B2(n_524), .Y(n_522) );
CKINVDCx6p67_ASAP7_75t_R g638 ( .A(n_357), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_357), .A2(n_368), .B1(n_709), .B2(n_710), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_357), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
AOI22xp5_ASAP7_75t_SL g800 ( .A1(n_357), .A2(n_718), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_357), .A2(n_718), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1621 ( .A1(n_357), .A2(n_368), .B1(n_1622), .B2(n_1623), .Y(n_1621) );
AND2x6_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
AND2x2_ASAP7_75t_L g514 ( .A(n_358), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g637 ( .A(n_358), .Y(n_637) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x6_ASAP7_75t_L g385 ( .A(n_359), .B(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g479 ( .A(n_360), .Y(n_479) );
INVx2_ASAP7_75t_SL g496 ( .A(n_360), .Y(n_496) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_360), .Y(n_585) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_360), .Y(n_604) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_360), .Y(n_683) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_360), .Y(n_688) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_360), .Y(n_976) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_360), .Y(n_1047) );
BUFx2_ASAP7_75t_L g1142 ( .A(n_360), .Y(n_1142) );
INVx1_ASAP7_75t_L g594 ( .A(n_361), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_367), .B2(n_368), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_363), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_429) );
INVx4_ASAP7_75t_L g640 ( .A(n_364), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_364), .A2(n_368), .B1(n_721), .B2(n_722), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_364), .A2(n_368), .B1(n_798), .B2(n_807), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_364), .A2(n_368), .B1(n_848), .B2(n_849), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_364), .A2(n_368), .B1(n_901), .B2(n_902), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_364), .A2(n_368), .B1(n_956), .B2(n_957), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_364), .A2(n_368), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_364), .A2(n_368), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_364), .A2(n_368), .B1(n_1158), .B2(n_1159), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_364), .A2(n_368), .B1(n_1195), .B2(n_1209), .Y(n_1208) );
AND2x4_ASAP7_75t_L g380 ( .A(n_365), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_SL g856 ( .A(n_365), .B(n_381), .Y(n_856) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx4_ASAP7_75t_L g641 ( .A(n_368), .Y(n_641) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_369), .Y(n_482) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_369), .Y(n_570) );
INVx2_ASAP7_75t_L g606 ( .A(n_369), .Y(n_606) );
INVx1_ASAP7_75t_L g875 ( .A(n_369), .Y(n_875) );
INVx1_ASAP7_75t_L g921 ( .A(n_369), .Y(n_921) );
INVx1_ASAP7_75t_L g1043 ( .A(n_369), .Y(n_1043) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g494 ( .A(n_370), .Y(n_494) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_370), .Y(n_562) );
INVx1_ASAP7_75t_L g685 ( .A(n_370), .Y(n_685) );
INVx1_ASAP7_75t_L g978 ( .A(n_370), .Y(n_978) );
INVx1_ASAP7_75t_L g593 ( .A(n_371), .Y(n_593) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_377), .B2(n_378), .C1(n_384), .C2(n_385), .Y(n_372) );
AOI222xp33_ASAP7_75t_L g853 ( .A1(n_374), .A2(n_385), .B1(n_854), .B2(n_855), .C1(n_856), .C2(n_857), .Y(n_853) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_375), .Y(n_489) );
INVx1_ASAP7_75t_L g499 ( .A(n_375), .Y(n_499) );
INVx1_ASAP7_75t_L g707 ( .A(n_375), .Y(n_707) );
BUFx4f_ASAP7_75t_L g758 ( .A(n_375), .Y(n_758) );
AND2x4_ASAP7_75t_L g1545 ( .A(n_375), .B(n_1546), .Y(n_1545) );
INVx2_ASAP7_75t_SL g1643 ( .A(n_375), .Y(n_1643) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_377), .A2(n_384), .B1(n_414), .B2(n_415), .C1(n_420), .C2(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx4f_ASAP7_75t_L g727 ( .A(n_380), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_380), .A2(n_385), .B1(n_791), .B2(n_794), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_380), .A2(n_385), .B1(n_1060), .B2(n_1061), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_380), .A2(n_385), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g520 ( .A(n_382), .Y(n_520) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g1531 ( .A(n_383), .Y(n_1531) );
INVx3_ASAP7_75t_L g521 ( .A(n_385), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g643 ( .A1(n_385), .A2(n_519), .B1(n_633), .B2(n_644), .C1(n_646), .C2(n_647), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g704 ( .A1(n_385), .A2(n_519), .B1(n_699), .B2(n_700), .C1(n_705), .C2(n_706), .Y(n_704) );
AOI222xp33_ASAP7_75t_L g723 ( .A1(n_385), .A2(n_724), .B1(n_725), .B2(n_726), .C1(n_727), .C2(n_728), .Y(n_723) );
AOI222xp33_ASAP7_75t_L g803 ( .A1(n_385), .A2(n_727), .B1(n_791), .B2(n_794), .C1(n_804), .C2(n_805), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_385), .A2(n_856), .B1(n_896), .B2(n_897), .C1(n_898), .C2(n_899), .Y(n_895) );
AOI222xp33_ASAP7_75t_L g958 ( .A1(n_385), .A2(n_727), .B1(n_959), .B2(n_960), .C1(n_961), .C2(n_962), .Y(n_958) );
AOI222xp33_ASAP7_75t_L g1008 ( .A1(n_385), .A2(n_489), .B1(n_856), .B2(n_1009), .C1(n_1010), .C2(n_1011), .Y(n_1008) );
AOI222xp33_ASAP7_75t_L g1110 ( .A1(n_385), .A2(n_856), .B1(n_910), .B2(n_1111), .C1(n_1112), .C2(n_1113), .Y(n_1110) );
AOI222xp33_ASAP7_75t_L g1153 ( .A1(n_385), .A2(n_498), .B1(n_856), .B2(n_1154), .C1(n_1155), .C2(n_1156), .Y(n_1153) );
AOI222xp33_ASAP7_75t_L g1210 ( .A1(n_385), .A2(n_727), .B1(n_1198), .B2(n_1200), .C1(n_1211), .C2(n_1212), .Y(n_1210) );
AOI222xp33_ASAP7_75t_L g1616 ( .A1(n_385), .A2(n_856), .B1(n_1617), .B2(n_1618), .C1(n_1619), .C2(n_1620), .Y(n_1616) );
BUFx3_ASAP7_75t_L g1534 ( .A(n_386), .Y(n_1534) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_387), .B(n_510), .C(n_513), .D(n_522), .Y(n_509) );
NAND4xp25_ASAP7_75t_SL g715 ( .A(n_387), .B(n_716), .C(n_720), .D(n_723), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g799 ( .A(n_387), .B(n_800), .C(n_803), .D(n_806), .Y(n_799) );
NAND4xp25_ASAP7_75t_L g846 ( .A(n_387), .B(n_847), .C(n_850), .D(n_853), .Y(n_846) );
NAND4xp25_ASAP7_75t_SL g951 ( .A(n_387), .B(n_952), .C(n_955), .D(n_958), .Y(n_951) );
NAND4xp25_ASAP7_75t_SL g1001 ( .A(n_387), .B(n_1002), .C(n_1005), .D(n_1008), .Y(n_1001) );
NAND4xp25_ASAP7_75t_L g1204 ( .A(n_387), .B(n_1205), .C(n_1208), .D(n_1210), .Y(n_1204) );
INVx5_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
CKINVDCx8_ASAP7_75t_R g648 ( .A(n_388), .Y(n_648) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_390), .Y(n_515) );
INVx1_ASAP7_75t_L g560 ( .A(n_390), .Y(n_560) );
INVx2_ASAP7_75t_L g645 ( .A(n_390), .Y(n_645) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_390), .Y(n_911) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_391), .Y(n_729) );
INVx1_ASAP7_75t_L g903 ( .A(n_391), .Y(n_903) );
AOI221xp5_ASAP7_75t_L g1102 ( .A1(n_391), .A2(n_437), .B1(n_1103), .B2(n_1114), .C(n_1124), .Y(n_1102) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
AND2x4_ASAP7_75t_L g525 ( .A(n_392), .B(n_394), .Y(n_525) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g501 ( .A(n_393), .B(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g1517 ( .A(n_394), .Y(n_1517) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g444 ( .A(n_395), .Y(n_444) );
OR2x6_ASAP7_75t_L g616 ( .A(n_395), .B(n_617), .Y(n_616) );
NAND4xp25_ASAP7_75t_SL g396 ( .A(n_397), .B(n_413), .C(n_429), .D(n_434), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_407), .B2(n_408), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_399), .A2(n_431), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_399), .A2(n_408), .B1(n_770), .B2(n_771), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_399), .A2(n_408), .B1(n_787), .B2(n_788), .Y(n_786) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_399), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
AOI22xp5_ASAP7_75t_SL g945 ( .A1(n_399), .A2(n_883), .B1(n_946), .B2(n_947), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_399), .A2(n_408), .B1(n_990), .B2(n_991), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_399), .A2(n_883), .B1(n_1017), .B2(n_1018), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_399), .A2(n_883), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g1176 ( .A1(n_399), .A2(n_883), .B1(n_1177), .B2(n_1178), .Y(n_1176) );
AOI22xp33_ASAP7_75t_SL g1194 ( .A1(n_399), .A2(n_774), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_403), .Y(n_399) );
AND2x4_ASAP7_75t_L g408 ( .A(n_400), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g658 ( .A(n_400), .Y(n_658) );
AND2x4_ASAP7_75t_L g883 ( .A(n_400), .B(n_409), .Y(n_883) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g428 ( .A(n_402), .Y(n_428) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_403), .Y(n_543) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_403), .Y(n_552) );
BUFx2_ASAP7_75t_L g738 ( .A(n_403), .Y(n_738) );
INVx1_ASAP7_75t_L g925 ( .A(n_403), .Y(n_925) );
BUFx2_ASAP7_75t_L g972 ( .A(n_403), .Y(n_972) );
INVx1_ASAP7_75t_L g1034 ( .A(n_403), .Y(n_1034) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_408), .A2(n_432), .B1(n_512), .B2(n_538), .Y(n_537) );
INVx5_ASAP7_75t_SL g651 ( .A(n_408), .Y(n_651) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g460 ( .A(n_411), .Y(n_460) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_411), .Y(n_544) );
INVx1_ASAP7_75t_L g934 ( .A(n_411), .Y(n_934) );
AND2x4_ASAP7_75t_L g418 ( .A(n_412), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g1137 ( .A(n_416), .Y(n_1137) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_417), .Y(n_1030) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g435 ( .A(n_418), .B(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
BUFx3_ASAP7_75t_L g530 ( .A(n_418), .Y(n_530) );
INVx1_ASAP7_75t_L g549 ( .A(n_418), .Y(n_549) );
BUFx3_ASAP7_75t_L g672 ( .A(n_418), .Y(n_672) );
BUFx2_ASAP7_75t_L g746 ( .A(n_418), .Y(n_746) );
INVx2_ASAP7_75t_L g532 ( .A(n_420), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_420), .A2(n_422), .B1(n_646), .B2(n_647), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_420), .A2(n_422), .B1(n_699), .B2(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g793 ( .A(n_420), .Y(n_793) );
INVx2_ASAP7_75t_L g834 ( .A(n_420), .Y(n_834) );
AOI222xp33_ASAP7_75t_SL g1064 ( .A1(n_420), .A2(n_795), .B1(n_1060), .B2(n_1061), .C1(n_1065), .C2(n_1066), .Y(n_1064) );
AOI222xp33_ASAP7_75t_L g1269 ( .A1(n_420), .A2(n_422), .B1(n_529), .B2(n_1246), .C1(n_1247), .C2(n_1265), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g1577 ( .A(n_421), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_422), .A2(n_791), .B1(n_794), .B2(n_833), .Y(n_832) );
AOI222xp33_ASAP7_75t_L g1197 ( .A1(n_422), .A2(n_792), .B1(n_879), .B2(n_1198), .C1(n_1199), .C2(n_1200), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1628 ( .A1(n_422), .A2(n_833), .B1(n_1619), .B2(n_1620), .Y(n_1628) );
AND2x4_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
AND2x4_ASAP7_75t_L g795 ( .A(n_423), .B(n_426), .Y(n_795) );
AND2x4_ASAP7_75t_L g1580 ( .A(n_423), .B(n_1578), .Y(n_1580) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_425), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g632 ( .A(n_425), .B(n_615), .Y(n_632) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g436 ( .A(n_427), .Y(n_436) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_428), .B(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_431), .A2(n_721), .B1(n_773), .B2(n_774), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_431), .A2(n_774), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_431), .A2(n_774), .B1(n_848), .B2(n_886), .Y(n_885) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_431), .A2(n_774), .B1(n_901), .B2(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_431), .A2(n_432), .B1(n_956), .B2(n_993), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_431), .A2(n_432), .B1(n_1006), .B2(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_431), .A2(n_774), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_431), .A2(n_432), .B1(n_1108), .B2(n_1123), .Y(n_1122) );
AOI22xp33_ASAP7_75t_SL g1179 ( .A1(n_431), .A2(n_432), .B1(n_1158), .B2(n_1180), .Y(n_1179) );
AOI22xp33_ASAP7_75t_SL g1201 ( .A1(n_431), .A2(n_883), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_431), .A2(n_774), .B1(n_1264), .B2(n_1271), .Y(n_1270) );
INVx5_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx4_ASAP7_75t_L g774 ( .A(n_433), .Y(n_774) );
NAND4xp25_ASAP7_75t_L g785 ( .A(n_434), .B(n_786), .C(n_789), .D(n_796), .Y(n_785) );
NAND3xp33_ASAP7_75t_SL g1063 ( .A(n_434), .B(n_1064), .C(n_1067), .Y(n_1063) );
NAND4xp25_ASAP7_75t_L g1193 ( .A(n_434), .B(n_1194), .C(n_1197), .D(n_1201), .Y(n_1193) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_434), .B(n_1269), .C(n_1270), .Y(n_1268) );
CKINVDCx11_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
AOI211xp5_ASAP7_75t_L g527 ( .A1(n_435), .A2(n_528), .B(n_529), .C(n_531), .Y(n_527) );
AOI211xp5_ASAP7_75t_SL g765 ( .A1(n_435), .A2(n_548), .B(n_766), .C(n_767), .Y(n_765) );
AOI211xp5_ASAP7_75t_L g877 ( .A1(n_435), .A2(n_878), .B(n_879), .C(n_880), .Y(n_877) );
AOI211xp5_ASAP7_75t_L g940 ( .A1(n_435), .A2(n_671), .B(n_941), .C(n_942), .Y(n_940) );
AOI211xp5_ASAP7_75t_L g986 ( .A1(n_435), .A2(n_671), .B(n_987), .C(n_988), .Y(n_986) );
AOI211xp5_ASAP7_75t_L g1013 ( .A1(n_435), .A2(n_879), .B(n_1014), .C(n_1015), .Y(n_1013) );
AOI211xp5_ASAP7_75t_L g1115 ( .A1(n_435), .A2(n_1116), .B(n_1117), .C(n_1118), .Y(n_1115) );
AOI211xp5_ASAP7_75t_L g1173 ( .A1(n_435), .A2(n_879), .B(n_1174), .C(n_1175), .Y(n_1173) );
OAI31xp33_ASAP7_75t_SL g649 ( .A1(n_437), .A2(n_650), .A3(n_652), .B(n_656), .Y(n_649) );
OAI31xp33_ASAP7_75t_SL g692 ( .A1(n_437), .A2(n_693), .A3(n_694), .B(n_701), .Y(n_692) );
AOI221x1_ASAP7_75t_L g784 ( .A1(n_437), .A2(n_729), .B1(n_785), .B2(n_799), .C(n_808), .Y(n_784) );
OAI31xp33_ASAP7_75t_L g827 ( .A1(n_437), .A2(n_828), .A3(n_829), .B(n_835), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g1062 ( .A1(n_437), .A2(n_1063), .B(n_1070), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1192 ( .A1(n_437), .A2(n_1193), .B1(n_1204), .B2(n_1213), .C(n_1214), .Y(n_1192) );
OAI21xp5_ASAP7_75t_L g1267 ( .A1(n_437), .A2(n_1268), .B(n_1272), .Y(n_1267) );
OAI31xp33_ASAP7_75t_L g1625 ( .A1(n_437), .A2(n_1626), .A3(n_1627), .B(n_1629), .Y(n_1625) );
CKINVDCx16_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
AOI31xp33_ASAP7_75t_L g764 ( .A1(n_438), .A2(n_765), .A3(n_769), .B(n_772), .Y(n_764) );
AOI31xp33_ASAP7_75t_L g876 ( .A1(n_438), .A2(n_877), .A3(n_881), .B(n_885), .Y(n_876) );
AOI31xp33_ASAP7_75t_SL g939 ( .A1(n_438), .A2(n_940), .A3(n_943), .B(n_945), .Y(n_939) );
AOI31xp33_ASAP7_75t_L g985 ( .A1(n_438), .A2(n_986), .A3(n_989), .B(n_992), .Y(n_985) );
AOI31xp33_ASAP7_75t_L g1012 ( .A1(n_438), .A2(n_1013), .A3(n_1016), .B(n_1019), .Y(n_1012) );
AND2x4_ASAP7_75t_L g500 ( .A(n_439), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g571 ( .A(n_439), .B(n_501), .Y(n_571) );
AND2x4_ASAP7_75t_L g1572 ( .A(n_439), .B(n_1573), .Y(n_1572) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_472), .Y(n_440) );
AOI33xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_446), .A3(n_454), .B1(n_461), .B2(n_464), .B3(n_466), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g1071 ( .A1(n_442), .A2(n_466), .B1(n_1072), .B2(n_1080), .C(n_1088), .Y(n_1071) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_442), .A2(n_466), .B1(n_1250), .B2(n_1255), .C(n_1259), .Y(n_1249) );
BUFx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_443), .B(n_542), .C(n_545), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_443), .B(n_667), .C(n_669), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_443), .B(n_811), .C(n_812), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g859 ( .A(n_443), .B(n_860), .C(n_861), .Y(n_859) );
INVx2_ASAP7_75t_L g966 ( .A(n_443), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g1022 ( .A(n_443), .B(n_1023), .C(n_1027), .Y(n_1022) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_443), .B(n_1130), .C(n_1134), .Y(n_1129) );
AOI33xp33_ASAP7_75t_L g1166 ( .A1(n_443), .A2(n_571), .A3(n_1167), .B1(n_1168), .B2(n_1170), .B3(n_1171), .Y(n_1166) );
NAND3xp33_ASAP7_75t_L g1631 ( .A(n_443), .B(n_1632), .C(n_1636), .Y(n_1631) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OR2x6_ASAP7_75t_L g474 ( .A(n_444), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g554 ( .A(n_444), .B(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g564 ( .A(n_444), .B(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g581 ( .A(n_444), .B(n_475), .Y(n_581) );
AND2x4_ASAP7_75t_L g732 ( .A(n_444), .B(n_445), .Y(n_732) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g547 ( .A(n_449), .Y(n_547) );
BUFx2_ASAP7_75t_L g816 ( .A(n_449), .Y(n_816) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g736 ( .A(n_450), .Y(n_736) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g465 ( .A(n_452), .Y(n_465) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_453), .Y(n_879) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_457), .B(n_1593), .Y(n_1600) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g668 ( .A(n_459), .Y(n_668) );
INVx2_ASAP7_75t_L g675 ( .A(n_459), .Y(n_675) );
INVx2_ASAP7_75t_SL g864 ( .A(n_459), .Y(n_864) );
INVx2_ASAP7_75t_L g1127 ( .A(n_459), .Y(n_1127) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g623 ( .A(n_460), .Y(n_623) );
INVx3_ASAP7_75t_L g1026 ( .A(n_460), .Y(n_1026) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_466), .B(n_674), .C(n_676), .Y(n_673) );
AOI33xp33_ASAP7_75t_L g731 ( .A1(n_466), .A2(n_732), .A3(n_733), .B1(n_737), .B2(n_741), .B3(n_743), .Y(n_731) );
AOI33xp33_ASAP7_75t_L g964 ( .A1(n_466), .A2(n_965), .A3(n_967), .B1(n_968), .B2(n_971), .B3(n_973), .Y(n_964) );
AOI33xp33_ASAP7_75t_L g1583 ( .A1(n_466), .A2(n_732), .A3(n_1584), .B1(n_1585), .B2(n_1586), .B3(n_1588), .Y(n_1583) );
INVx6_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx5_ASAP7_75t_L g928 ( .A(n_467), .Y(n_928) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g1593 ( .A(n_469), .B(n_1594), .Y(n_1593) );
INVx2_ASAP7_75t_L g555 ( .A(n_470), .Y(n_555) );
AOI33xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_477), .A3(n_483), .B1(n_490), .B2(n_497), .B3(n_500), .Y(n_472) );
AOI33xp33_ASAP7_75t_L g747 ( .A1(n_473), .A2(n_748), .A3(n_752), .B1(n_755), .B2(n_759), .B3(n_763), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g915 ( .A(n_473), .B(n_916), .C(n_918), .Y(n_915) );
AOI33xp33_ASAP7_75t_L g974 ( .A1(n_473), .A2(n_763), .A3(n_975), .B1(n_979), .B2(n_981), .B3(n_982), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_474), .Y(n_1230) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g565 ( .A(n_476), .Y(n_565) );
INVx2_ASAP7_75t_SL g1553 ( .A(n_476), .Y(n_1553) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_SL g1235 ( .A(n_479), .Y(n_1235) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g1237 ( .A(n_488), .Y(n_1237) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_SL g897 ( .A(n_489), .Y(n_897) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g1048 ( .A(n_492), .Y(n_1048) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g1169 ( .A(n_493), .Y(n_1169) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g984 ( .A(n_494), .Y(n_984) );
OR2x2_ASAP7_75t_L g1522 ( .A(n_494), .B(n_1523), .Y(n_1522) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g870 ( .A(n_496), .Y(n_870) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx4f_ASAP7_75t_L g763 ( .A(n_500), .Y(n_763) );
BUFx4f_ASAP7_75t_L g914 ( .A(n_500), .Y(n_914) );
INVx4_ASAP7_75t_L g1095 ( .A(n_500), .Y(n_1095) );
INVx2_ASAP7_75t_L g1541 ( .A(n_501), .Y(n_1541) );
AND2x4_ASAP7_75t_L g1528 ( .A(n_502), .B(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
XNOR2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AOI211xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_525), .B(n_526), .C(n_540), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_516), .B(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g1244 ( .A(n_514), .Y(n_1244) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_515), .Y(n_725) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_515), .Y(n_804) );
HB1xp67_ASAP7_75t_L g960 ( .A(n_515), .Y(n_960) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI31xp33_ASAP7_75t_L g634 ( .A1(n_525), .A2(n_635), .A3(n_639), .B(n_642), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_525), .A2(n_703), .B(n_711), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g845 ( .A1(n_525), .A2(n_846), .B(n_858), .C(n_876), .Y(n_845) );
OAI31xp33_ASAP7_75t_SL g1052 ( .A1(n_525), .A2(n_1053), .A3(n_1054), .B(n_1055), .Y(n_1052) );
AOI211x1_ASAP7_75t_L g1148 ( .A1(n_525), .A2(n_1149), .B(n_1160), .C(n_1172), .Y(n_1148) );
OAI31xp33_ASAP7_75t_L g1241 ( .A1(n_525), .A2(n_1242), .A3(n_1243), .B(n_1248), .Y(n_1241) );
OAI21xp5_ASAP7_75t_L g1614 ( .A1(n_525), .A2(n_1615), .B(n_1624), .Y(n_1614) );
AOI31xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_534), .A3(n_537), .B(n_539), .Y(n_526) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x6_ASAP7_75t_L g1595 ( .A(n_530), .B(n_1593), .Y(n_1595) );
AOI31xp33_ASAP7_75t_L g1172 ( .A1(n_539), .A2(n_1173), .A3(n_1176), .B(n_1179), .Y(n_1172) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_550), .C(n_556), .D(n_566), .Y(n_540) );
INVx2_ASAP7_75t_SL g740 ( .A(n_544), .Y(n_740) );
BUFx3_ASAP7_75t_L g742 ( .A(n_544), .Y(n_742) );
INVx2_ASAP7_75t_SL g970 ( .A(n_544), .Y(n_970) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_544), .Y(n_1223) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g670 ( .A(n_547), .Y(n_670) );
INVx2_ASAP7_75t_SL g677 ( .A(n_547), .Y(n_677) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .C(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g628 ( .A(n_554), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g813 ( .A(n_554), .B(n_814), .C(n_815), .Y(n_813) );
NAND3xp33_ASAP7_75t_L g862 ( .A(n_554), .B(n_863), .C(n_865), .Y(n_862) );
AOI33xp33_ASAP7_75t_L g1161 ( .A1(n_554), .A2(n_563), .A3(n_1162), .B1(n_1163), .B2(n_1164), .B3(n_1165), .Y(n_1161) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .C(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g587 ( .A(n_562), .Y(n_587) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_562), .Y(n_751) );
INVx1_ASAP7_75t_L g762 ( .A(n_562), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_563), .B(n_679), .C(n_682), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_563), .B(n_818), .C(n_819), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g866 ( .A(n_563), .B(n_867), .C(n_869), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g1039 ( .A(n_563), .B(n_1040), .C(n_1041), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1138 ( .A(n_563), .B(n_1139), .C(n_1141), .Y(n_1138) );
NAND3xp33_ASAP7_75t_L g1640 ( .A(n_563), .B(n_1641), .C(n_1644), .Y(n_1640) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .C(n_571), .Y(n_566) );
INVx1_ASAP7_75t_L g608 ( .A(n_571), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_571), .B(n_687), .C(n_689), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_571), .B(n_821), .C(n_824), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g871 ( .A(n_571), .B(n_872), .C(n_873), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_571), .B(n_1045), .C(n_1046), .Y(n_1044) );
NAND3xp33_ASAP7_75t_L g1143 ( .A(n_571), .B(n_1144), .C(n_1145), .Y(n_1143) );
NAND3xp33_ASAP7_75t_L g1645 ( .A(n_571), .B(n_1646), .C(n_1647), .Y(n_1645) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_660), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_634), .C(n_649), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_609), .Y(n_579) );
OAI33xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .A3(n_588), .B1(n_599), .B2(n_602), .B3(n_608), .Y(n_580) );
OAI22xp5_ASAP7_75t_SL g1088 ( .A1(n_581), .A2(n_1089), .B1(n_1095), .B2(n_1096), .Y(n_1088) );
OAI22xp5_ASAP7_75t_SL g1259 ( .A1(n_581), .A2(n_1095), .B1(n_1260), .B2(n_1263), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_586), .B2(n_587), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_583), .A2(n_586), .B1(n_619), .B2(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx4f_ASAP7_75t_L g919 ( .A(n_585), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_595), .B2(n_596), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_589), .A2(n_595), .B1(n_611), .B2(n_613), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_590), .A2(n_596), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g636 ( .A(n_592), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g1091 ( .A(n_592), .Y(n_1091) );
OR2x2_ASAP7_75t_L g1562 ( .A(n_592), .B(n_1523), .Y(n_1562) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_593), .B(n_594), .Y(n_598) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g1097 ( .A(n_597), .Y(n_1097) );
BUFx4f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g840 ( .A(n_598), .Y(n_840) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_598), .Y(n_1058) );
INVx2_ASAP7_75t_L g1093 ( .A(n_598), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g1228 ( .A(n_603), .Y(n_1228) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g1564 ( .A(n_604), .B(n_1546), .Y(n_1564) );
INVx1_ASAP7_75t_L g1555 ( .A(n_606), .Y(n_1555) );
OAI33xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_616), .A3(n_618), .B1(n_624), .B2(n_628), .B3(n_629), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_611), .A2(n_630), .B1(n_631), .B2(n_633), .Y(n_629) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g1079 ( .A(n_613), .Y(n_1079) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g625 ( .A(n_620), .Y(n_625) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g659 ( .A(n_621), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_622), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g926 ( .A(n_623), .Y(n_926) );
INVx1_ASAP7_75t_L g1218 ( .A(n_623), .Y(n_1218) );
AND2x4_ASAP7_75t_L g1592 ( .A(n_623), .B(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g831 ( .A(n_631), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_631), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_631), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1251) );
OAI22xp33_ASAP7_75t_SL g1256 ( .A1(n_631), .A2(n_1075), .B1(n_1257), .B2(n_1258), .Y(n_1256) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g654 ( .A(n_632), .Y(n_654) );
INVx2_ASAP7_75t_L g697 ( .A(n_632), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_643), .B(n_648), .Y(n_642) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g691 ( .A(n_645), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g703 ( .A(n_648), .B(n_704), .C(n_708), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g1103 ( .A(n_648), .B(n_1104), .C(n_1107), .D(n_1110), .Y(n_1103) );
NAND4xp25_ASAP7_75t_L g1149 ( .A(n_648), .B(n_1150), .C(n_1153), .D(n_1157), .Y(n_1149) );
NAND3xp33_ASAP7_75t_SL g1615 ( .A(n_648), .B(n_1616), .C(n_1621), .Y(n_1615) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_713), .B2(n_775), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
XOR2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_712), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_692), .C(n_702), .Y(n_664) );
AND4x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_673), .C(n_678), .D(n_686), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g789 ( .A1(n_671), .A2(n_790), .B1(n_791), .B2(n_792), .C1(n_794), .C2(n_795), .Y(n_789) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_671), .Y(n_1116) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g868 ( .A(n_681), .Y(n_868) );
INVx2_ASAP7_75t_L g750 ( .A(n_683), .Y(n_750) );
BUFx3_ASAP7_75t_L g913 ( .A(n_683), .Y(n_913) );
INVx2_ASAP7_75t_SL g1550 ( .A(n_683), .Y(n_1550) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
BUFx3_ASAP7_75t_L g983 ( .A(n_688), .Y(n_983) );
INVx2_ASAP7_75t_L g1537 ( .A(n_688), .Y(n_1537) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g1618 ( .A(n_707), .Y(n_1618) );
INVx2_ASAP7_75t_SL g775 ( .A(n_713), .Y(n_775) );
AOI211xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_729), .B(n_730), .C(n_764), .Y(n_714) );
OAI31xp33_ASAP7_75t_L g836 ( .A1(n_729), .A2(n_837), .A3(n_838), .B(n_842), .Y(n_836) );
AOI211x1_ASAP7_75t_SL g950 ( .A1(n_729), .A2(n_951), .B(n_963), .C(n_985), .Y(n_950) );
AOI211xp5_ASAP7_75t_L g1000 ( .A1(n_729), .A2(n_1001), .B(n_1012), .C(n_1021), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_747), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g929 ( .A(n_732), .B(n_930), .C(n_935), .Y(n_929) );
BUFx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_SL g938 ( .A(n_736), .Y(n_938) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_736), .Y(n_1029) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g1066 ( .A(n_745), .Y(n_1066) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_L g1582 ( .A(n_746), .B(n_1578), .Y(n_1582) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_SL g760 ( .A(n_750), .Y(n_760) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g917 ( .A(n_754), .Y(n_917) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g1212 ( .A(n_758), .Y(n_1212) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_1187), .B2(n_1188), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AO22x2_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_996), .B1(n_1185), .B2(n_1186), .Y(n_779) );
INVx1_ASAP7_75t_L g1185 ( .A(n_780), .Y(n_1185) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_887), .Y(n_780) );
AO22x2_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B1(n_843), .B2(n_844), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g835 ( .A(n_786), .Y(n_835) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g828 ( .A(n_796), .Y(n_828) );
INVxp67_ASAP7_75t_L g837 ( .A(n_800), .Y(n_837) );
INVxp67_ASAP7_75t_L g842 ( .A(n_806), .Y(n_842) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_809), .B(n_827), .C(n_836), .Y(n_826) );
AND4x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .C(n_817), .D(n_820), .Y(n_809) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx4_ASAP7_75t_L g980 ( .A(n_823), .Y(n_980) );
INVx2_ASAP7_75t_L g1140 ( .A(n_823), .Y(n_1140) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND4xp25_ASAP7_75t_L g858 ( .A(n_859), .B(n_862), .C(n_866), .D(n_871), .Y(n_858) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_948), .B2(n_995), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NOR3xp33_ASAP7_75t_L g890 ( .A(n_891), .B(n_904), .C(n_939), .Y(n_890) );
AOI31xp33_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_895), .A3(n_900), .B(n_903), .Y(n_891) );
INVx1_ASAP7_75t_L g1213 ( .A(n_903), .Y(n_1213) );
NAND4xp25_ASAP7_75t_L g904 ( .A(n_905), .B(n_915), .C(n_922), .D(n_929), .Y(n_904) );
NAND3xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_912), .C(n_914), .Y(n_905) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx6f_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g1552 ( .A(n_911), .Y(n_1552) );
AND2x4_ASAP7_75t_L g1556 ( .A(n_911), .B(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_927), .C(n_928), .Y(n_922) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g1081 ( .A(n_925), .Y(n_1081) );
INVx1_ASAP7_75t_L g1633 ( .A(n_925), .Y(n_1633) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_928), .B(n_1032), .C(n_1037), .Y(n_1031) );
NAND3xp33_ASAP7_75t_L g1125 ( .A(n_928), .B(n_1126), .C(n_1128), .Y(n_1125) );
NAND3xp33_ASAP7_75t_L g1220 ( .A(n_928), .B(n_1221), .C(n_1224), .Y(n_1220) );
NAND3xp33_ASAP7_75t_L g1637 ( .A(n_928), .B(n_1638), .C(n_1639), .Y(n_1637) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g1133 ( .A(n_934), .Y(n_1133) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_938), .Y(n_1038) );
INVx1_ASAP7_75t_L g1136 ( .A(n_938), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1598 ( .A(n_938), .B(n_1593), .Y(n_1598) );
INVx1_ASAP7_75t_L g995 ( .A(n_948), .Y(n_995) );
INVx1_ASAP7_75t_L g994 ( .A(n_950), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_974), .Y(n_963) );
NAND3xp33_ASAP7_75t_L g1215 ( .A(n_965), .B(n_1216), .C(n_1219), .Y(n_1215) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g1229 ( .A(n_978), .Y(n_1229) );
INVx1_ASAP7_75t_L g1186 ( .A(n_996), .Y(n_1186) );
AO22x2_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_1099), .B1(n_1100), .B2(n_1184), .Y(n_996) );
INVx1_ASAP7_75t_L g1184 ( .A(n_997), .Y(n_1184) );
XNOR2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_1050), .Y(n_997) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1000), .Y(n_1049) );
NAND4xp25_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1031), .C(n_1039), .D(n_1044), .Y(n_1021) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_1025), .Y(n_1024) );
INVx2_ASAP7_75t_L g1587 ( .A(n_1025), .Y(n_1587) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1026), .Y(n_1036) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1026), .Y(n_1083) );
INVx2_ASAP7_75t_L g1635 ( .A(n_1026), .Y(n_1635) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
NAND3x1_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1062), .C(n_1071), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
OAI21xp5_ASAP7_75t_SL g1538 ( .A1(n_1057), .A2(n_1539), .B(n_1540), .Y(n_1538) );
INVx2_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1096 ( .A1(n_1065), .A2(n_1068), .B1(n_1090), .B2(n_1097), .C(n_1098), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1074), .A2(n_1075), .B1(n_1077), .B2(n_1078), .Y(n_1073) );
INVx3_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1089 ( .A1(n_1085), .A2(n_1087), .B1(n_1090), .B2(n_1092), .C(n_1094), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1091), .Y(n_1261) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_1092), .A2(n_1252), .B1(n_1254), .B2(n_1261), .C(n_1262), .Y(n_1260) );
OAI221xp5_ASAP7_75t_L g1263 ( .A1(n_1092), .A2(n_1261), .B1(n_1264), .B2(n_1265), .C(n_1266), .Y(n_1263) );
BUFx3_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1095), .Y(n_1232) );
INVxp67_ASAP7_75t_SL g1099 ( .A(n_1100), .Y(n_1099) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1146), .B1(n_1147), .B2(n_1183), .Y(n_1100) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1101), .Y(n_1183) );
NAND3xp33_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1119), .C(n_1122), .Y(n_1114) );
NAND4xp25_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1129), .C(n_1138), .D(n_1143), .Y(n_1124) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1148), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1166), .Y(n_1160) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
XNOR2x2_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1238), .Y(n_1189) );
XNOR2xp5_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .Y(n_1190) );
NAND4xp25_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1220), .C(n_1225), .D(n_1231), .Y(n_1214) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
NAND3xp33_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1227), .C(n_1230), .Y(n_1225) );
NAND3xp33_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1233), .C(n_1236), .Y(n_1231) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
XNOR2xp5_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1240), .Y(n_1238) );
NAND3x1_ASAP7_75t_SL g1240 ( .A(n_1241), .B(n_1249), .C(n_1267), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1511), .B1(n_1512), .B2(n_1602), .C(n_1607), .Y(n_1273) );
AOI211xp5_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1422), .B(n_1464), .C(n_1490), .Y(n_1274) );
NAND5xp2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1384), .C(n_1409), .D(n_1414), .E(n_1419), .Y(n_1275) );
AOI21xp5_ASAP7_75t_L g1276 ( .A1(n_1277), .A2(n_1355), .B(n_1363), .Y(n_1276) );
OAI211xp5_ASAP7_75t_L g1277 ( .A1(n_1278), .A2(n_1315), .B(n_1325), .C(n_1349), .Y(n_1277) );
INVxp67_ASAP7_75t_SL g1278 ( .A(n_1279), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1304), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_1281), .A2(n_1340), .B1(n_1446), .B2(n_1447), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1301), .Y(n_1281) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1282), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1282), .B(n_1367), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1407 ( .A(n_1282), .B(n_1305), .Y(n_1407) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1282), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1282), .B(n_1356), .Y(n_1452) );
AOI221xp5_ASAP7_75t_L g1453 ( .A1(n_1282), .A2(n_1426), .B1(n_1454), .B2(n_1457), .C(n_1461), .Y(n_1453) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1282), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1295), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1290), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1286), .B(n_1291), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1289), .Y(n_1286) );
HB1xp67_ASAP7_75t_L g1656 ( .A(n_1287), .Y(n_1656) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1289), .Y(n_1298) );
AND2x4_ASAP7_75t_L g1292 ( .A(n_1290), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_1291), .B(n_1294), .Y(n_1314) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
BUFx3_ASAP7_75t_L g1330 ( .A(n_1296), .Y(n_1330) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1296), .Y(n_1360) );
AND2x4_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1299), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1297), .B(n_1299), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1654 ( .A(n_1297), .Y(n_1654) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
AND2x4_ASAP7_75t_L g1300 ( .A(n_1298), .B(n_1299), .Y(n_1300) );
INVx2_ASAP7_75t_L g1308 ( .A(n_1300), .Y(n_1308) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1301), .Y(n_1348) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1301), .Y(n_1367) );
BUFx6f_ASAP7_75t_L g1405 ( .A(n_1301), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1301), .B(n_1351), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1301), .B(n_1357), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1303), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1304), .B(n_1383), .Y(n_1434) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1304), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1304), .B(n_1394), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1304), .B(n_1366), .Y(n_1510) );
BUFx3_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_1305), .Y(n_1339) );
NOR2xp33_ASAP7_75t_L g1350 ( .A(n_1305), .B(n_1351), .Y(n_1350) );
BUFx2_ASAP7_75t_L g1391 ( .A(n_1305), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1305), .B(n_1322), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1305), .B(n_1426), .Y(n_1425) );
INVx2_ASAP7_75t_SL g1305 ( .A(n_1306), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1306), .B(n_1371), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1306), .B(n_1351), .Y(n_1504) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1308), .Y(n_1331) );
OAI22xp5_ASAP7_75t_SL g1359 ( .A1(n_1308), .A2(n_1360), .B1(n_1361), .B2(n_1362), .Y(n_1359) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_1311), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
HB1xp67_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1314), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1315), .B(n_1386), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1315), .B(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
AOI221xp5_ASAP7_75t_L g1424 ( .A1(n_1316), .A2(n_1373), .B1(n_1399), .B2(n_1425), .C(n_1427), .Y(n_1424) );
A2O1A1Ixp33_ASAP7_75t_SL g1441 ( .A1(n_1316), .A2(n_1380), .B(n_1442), .C(n_1443), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1322), .Y(n_1316) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1317), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1448 ( .A(n_1317), .B(n_1322), .Y(n_1448) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1318), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1318), .B(n_1343), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1318), .B(n_1344), .Y(n_1395) );
INVxp67_ASAP7_75t_SL g1401 ( .A(n_1318), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1318), .B(n_1322), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1320), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1322), .B(n_1341), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1322), .B(n_1353), .Y(n_1352) );
CKINVDCx5p33_ASAP7_75t_R g1371 ( .A(n_1322), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1322), .B(n_1400), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1322), .B(n_1395), .Y(n_1421) );
NOR2xp33_ASAP7_75t_L g1432 ( .A(n_1322), .B(n_1342), .Y(n_1432) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1322), .B(n_1375), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1322), .B(n_1378), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1322), .B(n_1342), .Y(n_1481) );
HB1xp67_ASAP7_75t_L g1493 ( .A(n_1322), .Y(n_1493) );
AND2x4_ASAP7_75t_SL g1322 ( .A(n_1323), .B(n_1324), .Y(n_1322) );
OAI21xp5_ASAP7_75t_SL g1325 ( .A1(n_1326), .A2(n_1338), .B(n_1347), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g1444 ( .A1(n_1326), .A2(n_1357), .B1(n_1445), .B2(n_1449), .C(n_1451), .Y(n_1444) );
INVx2_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1327), .B(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1327), .B(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1331), .Y(n_1511) );
OAI22xp33_ASAP7_75t_L g1332 ( .A1(n_1333), .A2(n_1334), .B1(n_1335), .B2(n_1336), .Y(n_1332) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
OAI31xp33_ASAP7_75t_L g1466 ( .A1(n_1338), .A2(n_1410), .A3(n_1467), .B(n_1469), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1339), .B(n_1378), .Y(n_1377) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1339), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1339), .B(n_1432), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1339), .B(n_1366), .Y(n_1463) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1343), .B(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1344), .B(n_1401), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1346), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1348), .B(n_1357), .Y(n_1388) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1348), .Y(n_1403) );
OAI32xp33_ASAP7_75t_L g1427 ( .A1(n_1348), .A2(n_1378), .A3(n_1405), .B1(n_1428), .B2(n_1430), .Y(n_1427) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1348), .B(n_1357), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1348), .B(n_1356), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1352), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1351), .B(n_1367), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1351), .B(n_1356), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1353), .B(n_1371), .Y(n_1383) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1353), .Y(n_1497) );
NAND2xp5_ASAP7_75t_SL g1365 ( .A(n_1356), .B(n_1366), .Y(n_1365) );
AOI32xp33_ASAP7_75t_L g1368 ( .A1(n_1356), .A2(n_1357), .A3(n_1369), .B1(n_1374), .B2(n_1376), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1356), .B(n_1413), .Y(n_1500) );
CKINVDCx6p67_ASAP7_75t_R g1356 ( .A(n_1357), .Y(n_1356) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1357), .B(n_1373), .Y(n_1418) );
CKINVDCx5p33_ASAP7_75t_R g1423 ( .A(n_1357), .Y(n_1423) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1357), .B(n_1504), .Y(n_1503) );
OR2x6_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1359), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1368), .B1(n_1379), .B2(n_1381), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1366), .Y(n_1396) );
AOI211xp5_ASAP7_75t_L g1433 ( .A1(n_1366), .A2(n_1434), .B(n_1435), .C(n_1444), .Y(n_1433) );
INVxp67_ASAP7_75t_SL g1369 ( .A(n_1370), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1372), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1371), .B(n_1378), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1371), .B(n_1395), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1371), .B(n_1400), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1460 ( .A(n_1371), .B(n_1377), .Y(n_1460) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_1371), .B(n_1455), .Y(n_1498) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
OAI21xp5_ASAP7_75t_SL g1409 ( .A1(n_1378), .A2(n_1410), .B(n_1411), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1378), .B(n_1402), .Y(n_1479) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1383), .Y(n_1381) );
AOI311xp33_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1388), .A3(n_1389), .B(n_1392), .C(n_1397), .Y(n_1384) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1388), .B(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1388), .Y(n_1482) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1390), .B(n_1421), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1390), .B(n_1439), .Y(n_1438) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1391), .B(n_1413), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1391), .B(n_1395), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_1391), .B(n_1403), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1391), .B(n_1456), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1391), .B(n_1439), .Y(n_1459) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1391), .B(n_1408), .Y(n_1468) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1396), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1508 ( .A1(n_1393), .A2(n_1405), .B1(n_1509), .B2(n_1510), .Y(n_1508) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
OAI21xp33_ASAP7_75t_L g1437 ( .A1(n_1394), .A2(n_1438), .B(n_1440), .Y(n_1437) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1395), .Y(n_1496) );
OAI21xp33_ASAP7_75t_SL g1397 ( .A1(n_1398), .A2(n_1403), .B(n_1404), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
NAND2xp67_ASAP7_75t_L g1489 ( .A(n_1399), .B(n_1426), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1399), .B(n_1471), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1402), .Y(n_1399) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1400), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1400), .B(n_1429), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1406), .Y(n_1404) );
CKINVDCx14_ASAP7_75t_R g1458 ( .A(n_1405), .Y(n_1458) );
NOR2xp33_ASAP7_75t_SL g1488 ( .A(n_1406), .B(n_1450), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1408), .Y(n_1406) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1410), .Y(n_1506) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1413), .Y(n_1436) );
INVxp67_ASAP7_75t_SL g1414 ( .A(n_1415), .Y(n_1414) );
NOR2xp33_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1418), .Y(n_1415) );
OAI211xp5_ASAP7_75t_L g1435 ( .A1(n_1416), .A2(n_1436), .B(n_1437), .C(n_1441), .Y(n_1435) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1418), .Y(n_1440) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1421), .Y(n_1507) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_1423), .A2(n_1424), .B(n_1433), .C(n_1453), .Y(n_1422) );
AOI221xp5_ASAP7_75t_L g1474 ( .A1(n_1423), .A2(n_1426), .B1(n_1475), .B2(n_1483), .C(n_1485), .Y(n_1474) );
OAI22xp33_ASAP7_75t_SL g1485 ( .A1(n_1423), .A2(n_1486), .B1(n_1488), .B2(n_1489), .Y(n_1485) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
OAI21xp33_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1459), .B(n_1460), .Y(n_1457) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
O2A1O1Ixp33_ASAP7_75t_L g1501 ( .A1(n_1463), .A2(n_1502), .B(n_1505), .C(n_1508), .Y(n_1501) );
A2O1A1Ixp33_ASAP7_75t_L g1464 ( .A1(n_1465), .A2(n_1466), .B(n_1473), .C(n_1474), .Y(n_1464) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1471), .B(n_1484), .Y(n_1483) );
INVx3_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_1476), .A2(n_1478), .B1(n_1480), .B2(n_1482), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
A2O1A1Ixp33_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1498), .B(n_1499), .C(n_1501), .Y(n_1490) );
INVxp67_ASAP7_75t_SL g1491 ( .A(n_1492), .Y(n_1491) );
NOR2xp33_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1494), .Y(n_1492) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1497), .Y(n_1495) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVxp67_ASAP7_75t_SL g1502 ( .A(n_1503), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1506), .B(n_1507), .Y(n_1505) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
HB1xp67_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
XNOR2xp5_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1601), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1574), .Y(n_1515) );
AOI22xp5_ASAP7_75t_L g1516 ( .A1(n_1517), .A2(n_1518), .B1(n_1565), .B2(n_1566), .Y(n_1516) );
NAND3xp33_ASAP7_75t_SL g1518 ( .A(n_1519), .B(n_1542), .C(n_1559), .Y(n_1518) );
AOI211xp5_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1521), .B(n_1525), .C(n_1535), .Y(n_1519) );
INVx4_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVx2_ASAP7_75t_L g1546 ( .A(n_1523), .Y(n_1546) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1524), .Y(n_1529) );
INVx2_ASAP7_75t_SL g1526 ( .A(n_1527), .Y(n_1526) );
AND2x4_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1530), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1528), .B(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1528), .Y(n_1558) );
INVx2_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
INVx2_ASAP7_75t_SL g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_1539), .A2(n_1590), .B1(n_1591), .B2(n_1595), .Y(n_1589) );
AOI221xp5_ASAP7_75t_L g1542 ( .A1(n_1543), .A2(n_1547), .B1(n_1548), .B2(n_1554), .C(n_1556), .Y(n_1542) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx2_ASAP7_75t_SL g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_SL g1557 ( .A(n_1558), .Y(n_1557) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_1560), .A2(n_1561), .B1(n_1563), .B2(n_1564), .Y(n_1559) );
INVx6_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx5_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1571), .Y(n_1567) );
INVx3_ASAP7_75t_L g1578 ( .A(n_1569), .Y(n_1578) );
INVx2_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
AND4x1_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1583), .C(n_1589), .D(n_1596), .Y(n_1574) );
AOI221xp5_ASAP7_75t_L g1575 ( .A1(n_1576), .A2(n_1579), .B1(n_1580), .B2(n_1581), .C(n_1582), .Y(n_1575) );
AND2x4_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1578), .Y(n_1576) );
BUFx2_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
AOI22xp33_ASAP7_75t_L g1596 ( .A1(n_1597), .A2(n_1598), .B1(n_1599), .B2(n_1600), .Y(n_1596) );
CKINVDCx5p33_ASAP7_75t_R g1602 ( .A(n_1603), .Y(n_1602) );
BUFx2_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVxp33_ASAP7_75t_SL g1608 ( .A(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
HB1xp67_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
NAND3x1_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1625), .C(n_1630), .Y(n_1613) );
AND4x1_ASAP7_75t_L g1630 ( .A(n_1631), .B(n_1637), .C(n_1640), .D(n_1645), .Y(n_1630) );
INVx2_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
CKINVDCx5p33_ASAP7_75t_R g1649 ( .A(n_1650), .Y(n_1649) );
A2O1A1Ixp33_ASAP7_75t_L g1652 ( .A1(n_1651), .A2(n_1653), .B(n_1655), .C(n_1657), .Y(n_1652) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
endmodule