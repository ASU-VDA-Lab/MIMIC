module fake_jpeg_4214_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_8),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_44),
.B1(n_25),
.B2(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_54),
.B1(n_57),
.B2(n_16),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_55),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_56),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_31),
.B(n_23),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_16),
.B(n_32),
.C(n_28),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_39),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_69),
.B1(n_83),
.B2(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_72),
.Y(n_110)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_78),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_77),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_35),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_106),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_58),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_103),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_58),
.C(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_108),
.C(n_63),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_59),
.B1(n_55),
.B2(n_37),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_105),
.B1(n_107),
.B2(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_63),
.B1(n_83),
.B2(n_84),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_59),
.B1(n_34),
.B2(n_33),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_80),
.B1(n_45),
.B2(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_67),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_34),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_33),
.B1(n_32),
.B2(n_18),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_37),
.B1(n_45),
.B2(n_18),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_37),
.C(n_45),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_26),
.B1(n_22),
.B2(n_21),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_115),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_R g113 ( 
.A(n_90),
.B(n_63),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_117),
.B(n_127),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_110),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_121),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_75),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_107),
.B(n_105),
.C(n_97),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_128),
.B(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_67),
.B1(n_73),
.B2(n_62),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_134),
.B1(n_102),
.B2(n_86),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_77),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_108),
.C(n_102),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_77),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_73),
.B(n_74),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_133),
.B1(n_135),
.B2(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_76),
.B1(n_19),
.B2(n_21),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_144),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_111),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_149),
.Y(n_167)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_91),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_135),
.B(n_115),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_24),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_24),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_28),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_172),
.B1(n_173),
.B2(n_138),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_132),
.B1(n_128),
.B2(n_116),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_149),
.B1(n_137),
.B2(n_155),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_179),
.B(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_82),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_22),
.B(n_19),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_182),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_93),
.B(n_82),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_93),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_174),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_191),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_197),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_138),
.B1(n_147),
.B2(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_196),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_141),
.C(n_138),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_201),
.C(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_143),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_158),
.B1(n_159),
.B2(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_199),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_161),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_176),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_136),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_88),
.B1(n_94),
.B2(n_87),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_87),
.C(n_31),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_163),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_166),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_192),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_175),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_208),
.C(n_213),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_165),
.B(n_170),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_186),
.B(n_196),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_180),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.C(n_179),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_188),
.B(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_165),
.C(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_195),
.C(n_186),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_202),
.B1(n_193),
.B2(n_169),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_217),
.A2(n_218),
.B(n_216),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_225),
.C(n_227),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_194),
.B1(n_198),
.B2(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_177),
.B1(n_168),
.B2(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_226),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_210),
.B(n_1),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_204),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_208),
.C(n_213),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_197),
.C(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_215),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_230),
.B(n_232),
.Y(n_240)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_6),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_233),
.A2(n_219),
.B1(n_222),
.B2(n_5),
.Y(n_237)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_7),
.CI(n_10),
.CON(n_247),
.SN(n_247)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_243),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_235),
.B1(n_232),
.B2(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_231),
.C(n_236),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_7),
.B(n_9),
.Y(n_243)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_SL g246 ( 
.A1(n_240),
.A2(n_7),
.A3(n_9),
.B(n_10),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_251),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_238),
.A3(n_248),
.B1(n_245),
.B2(n_244),
.C1(n_247),
.C2(n_13),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_11),
.B(n_15),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_15),
.Y(n_256)
);


endmodule