module fake_jpeg_26024_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_20),
.B1(n_18),
.B2(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_25),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_45),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_54),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_43),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_21),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_2),
.B(n_3),
.Y(n_68)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_30),
.B1(n_44),
.B2(n_26),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_69),
.B1(n_41),
.B2(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_73),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_54),
.B1(n_48),
.B2(n_46),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_19),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_59),
.C(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_58),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_88),
.B(n_41),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_84),
.B1(n_41),
.B2(n_42),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_83),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_76),
.B1(n_71),
.B2(n_70),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_11),
.A3(n_16),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_66),
.B(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_68),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_98),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_14),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_86),
.B(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_82),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_19),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_87),
.B1(n_90),
.B2(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_78),
.B1(n_77),
.B2(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_92),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_98),
.C(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_112),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_115),
.Y(n_118)
);

OA21x2_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_16),
.B(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_114),
.B(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_120),
.B(n_104),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_104),
.B1(n_109),
.B2(n_103),
.C(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_111),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_124),
.B1(n_15),
.B2(n_7),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_113),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_116),
.A3(n_15),
.B1(n_7),
.B2(n_6),
.C1(n_3),
.C2(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_127),
.C(n_13),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);


endmodule