module fake_jpeg_16661_n_358 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_22),
.A2(n_0),
.B(n_1),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_26),
.C(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_46),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_19),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_18),
.B1(n_35),
.B2(n_27),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_64),
.B1(n_68),
.B2(n_24),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_35),
.B1(n_25),
.B2(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_41),
.B1(n_46),
.B2(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_35),
.B1(n_25),
.B2(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_66),
.B(n_52),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_28),
.B1(n_24),
.B2(n_32),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_19),
.B1(n_23),
.B2(n_32),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_52),
.B1(n_58),
.B2(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_94),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_42),
.C(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_45),
.B1(n_53),
.B2(n_51),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_50),
.B1(n_53),
.B2(n_51),
.Y(n_91)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_50),
.B1(n_51),
.B2(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_40),
.B1(n_23),
.B2(n_29),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_104),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_13),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_26),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_57),
.B1(n_65),
.B2(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_76),
.B1(n_69),
.B2(n_74),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_60),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_61),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_67),
.B(n_78),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_38),
.B(n_37),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_87),
.B1(n_88),
.B2(n_97),
.Y(n_139)
);

AO21x2_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_42),
.B(n_61),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_88),
.B1(n_100),
.B2(n_106),
.Y(n_146)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_92),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_42),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_76),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_91),
.A2(n_29),
.B1(n_31),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_130),
.A2(n_85),
.B1(n_99),
.B2(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_15),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_105),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_30),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_48),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_37),
.C(n_38),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_146),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_85),
.B1(n_83),
.B2(n_82),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_85),
.B1(n_95),
.B2(n_106),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_153),
.B(n_163),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_106),
.B(n_38),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_31),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_92),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_113),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_10),
.B1(n_17),
.B2(n_15),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_160),
.A2(n_166),
.B1(n_120),
.B2(n_109),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_0),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_121),
.B(n_0),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_134),
.B1(n_124),
.B2(n_108),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_96),
.B(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_92),
.B1(n_30),
.B2(n_33),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_159),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_187),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_188),
.B1(n_190),
.B2(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_113),
.B1(n_125),
.B2(n_123),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_155),
.B1(n_166),
.B2(n_138),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_192),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_118),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_183),
.B(n_164),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_114),
.B(n_118),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_112),
.C(n_116),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_198),
.C(n_160),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_130),
.B(n_30),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_162),
.B(n_158),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_123),
.B1(n_132),
.B2(n_135),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_120),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_161),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_142),
.A2(n_155),
.B1(n_163),
.B2(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_33),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_216),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_221),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_222),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_213),
.C(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_225),
.B1(n_177),
.B2(n_186),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_226),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_196),
.B1(n_197),
.B2(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_143),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_178),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_229),
.A2(n_214),
.B1(n_207),
.B2(n_219),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_177),
.B1(n_179),
.B2(n_190),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_245),
.B1(n_248),
.B2(n_250),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_256),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_240),
.C(n_255),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_182),
.C(n_183),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_193),
.B1(n_173),
.B2(n_177),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_227),
.A2(n_182),
.B1(n_187),
.B2(n_180),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_9),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_209),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_145),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_224),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_217),
.C(n_202),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_145),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_229),
.B(n_236),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_257),
.A2(n_259),
.B(n_264),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_201),
.B(n_216),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_205),
.C(n_207),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_270),
.C(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_211),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_272),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_237),
.C(n_238),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_211),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_223),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_279),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_1),
.B(n_2),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_231),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_226),
.B1(n_96),
.B2(n_10),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_280),
.A2(n_250),
.B1(n_249),
.B2(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_291),
.C(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_288),
.Y(n_305)
);

BUFx12_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_260),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_236),
.B(n_245),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_257),
.B(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_256),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_290),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_238),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_9),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_258),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_4),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_311),
.B(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

OAI221xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_267),
.B1(n_279),
.B2(n_268),
.C(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_266),
.C(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_313),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_283),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_262),
.C(n_270),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_261),
.B(n_263),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_263),
.C(n_261),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_297),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_267),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_285),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_321),
.B(n_325),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_313),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_322),
.C(n_309),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_294),
.B1(n_285),
.B2(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_320),
.B(n_326),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_312),
.A2(n_281),
.B(n_283),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_311),
.A2(n_287),
.B1(n_281),
.B2(n_297),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_295),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_284),
.Y(n_330)
);

XNOR2x2_ASAP7_75t_SL g334 ( 
.A(n_329),
.B(n_287),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_330),
.B(n_331),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_328),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_286),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g346 ( 
.A1(n_332),
.A2(n_336),
.B(n_326),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_303),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_335),
.C(n_339),
.Y(n_342)
);

OAI321xp33_ASAP7_75t_L g347 ( 
.A1(n_334),
.A2(n_12),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C(n_17),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_5),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_10),
.C(n_6),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_332),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_341),
.B(n_346),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_325),
.B(n_329),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_343),
.A2(n_344),
.B(n_347),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_SL g344 ( 
.A(n_338),
.B(n_319),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_318),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_6),
.C(n_7),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_350),
.C(n_352),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_340),
.C(n_341),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_7),
.C(n_12),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_349),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_351),
.B(n_13),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_354),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_13),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_14),
.Y(n_358)
);


endmodule