module fake_jpeg_15632_n_344 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.C(n_1),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_48),
.B(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_21),
.B1(n_16),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_67),
.B1(n_35),
.B2(n_28),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_19),
.C(n_17),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_29),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_69),
.Y(n_92)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_36),
.Y(n_85)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_35),
.B1(n_41),
.B2(n_17),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_62),
.B1(n_41),
.B2(n_70),
.Y(n_103)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_62),
.B1(n_47),
.B2(n_11),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_15),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_90),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_14),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_14),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_94),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_112),
.B1(n_95),
.B2(n_98),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_106),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_108),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_62),
.B1(n_56),
.B2(n_19),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_78),
.B(n_26),
.Y(n_147)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_81),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_56),
.B1(n_36),
.B2(n_49),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_64),
.B1(n_80),
.B2(n_74),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

AO21x1_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_64),
.B(n_42),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_42),
.C(n_49),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_90),
.CI(n_88),
.CON(n_130),
.SN(n_130)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_18),
.B1(n_24),
.B2(n_30),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_80),
.B1(n_24),
.B2(n_30),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_128),
.B1(n_144),
.B2(n_147),
.Y(n_157)
);

AOI22x1_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_87),
.B1(n_64),
.B2(n_98),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_102),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_91),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_93),
.B1(n_81),
.B2(n_78),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_143),
.B1(n_150),
.B2(n_152),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_141),
.B(n_145),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_140),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_96),
.B(n_89),
.C(n_92),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_122),
.B1(n_109),
.B2(n_124),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_46),
.B(n_69),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_92),
.B(n_74),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_126),
.B(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_42),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_151),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_34),
.B1(n_42),
.B2(n_31),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_114),
.B(n_46),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_107),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_104),
.B1(n_108),
.B2(n_113),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_140),
.B1(n_152),
.B2(n_141),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_105),
.C(n_115),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_174),
.C(n_175),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_177),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_149),
.B(n_151),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_100),
.C(n_126),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_102),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_147),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_100),
.C(n_117),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_127),
.C(n_144),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_146),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_209),
.B(n_69),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_128),
.B1(n_136),
.B2(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_207),
.B1(n_208),
.B2(n_156),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_137),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_201),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_161),
.A2(n_128),
.B1(n_154),
.B2(n_140),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_200),
.B1(n_173),
.B2(n_155),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_206),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_167),
.B1(n_155),
.B2(n_165),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_129),
.B1(n_141),
.B2(n_150),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_34),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_178),
.B(n_170),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_139),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_99),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_119),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_135),
.B1(n_142),
.B2(n_111),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_135),
.B1(n_117),
.B2(n_99),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_22),
.B(n_92),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_187),
.B1(n_191),
.B2(n_193),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_183),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_219),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_232),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_208),
.A2(n_157),
.B1(n_162),
.B2(n_168),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_157),
.B1(n_186),
.B2(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_159),
.B1(n_160),
.B2(n_172),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_182),
.B1(n_200),
.B2(n_196),
.Y(n_243)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

NAND2x1p5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_178),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_231),
.B(n_235),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_176),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_210),
.C(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_184),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_198),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_191),
.B(n_209),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_230),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_224),
.A2(n_227),
.B1(n_214),
.B2(n_229),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_211),
.C(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_250),
.C(n_256),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_202),
.B1(n_195),
.B2(n_99),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_235),
.A2(n_92),
.B1(n_89),
.B2(n_86),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_61),
.C(n_69),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_220),
.B(n_30),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_34),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_259),
.A2(n_271),
.B1(n_255),
.B2(n_9),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_222),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_264),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_233),
.C(n_43),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_266),
.C(n_270),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_43),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_267),
.B(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_31),
.C(n_27),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_24),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_275),
.C(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_31),
.C(n_27),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_27),
.C(n_18),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_244),
.B(n_12),
.CI(n_10),
.CON(n_277),
.SN(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_10),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_0),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_239),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_261),
.C(n_275),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_240),
.C(n_256),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_271),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_284),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_238),
.B1(n_251),
.B2(n_253),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_285),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_270),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_274),
.A2(n_240),
.B(n_241),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_289),
.B(n_277),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_251),
.B(n_243),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_248),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_310),
.C(n_283),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_298),
.C(n_4),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_261),
.C(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_295),
.C(n_281),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_288),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_308),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_246),
.B(n_276),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_305),
.B(n_4),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_279),
.A2(n_2),
.B(n_4),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_2),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_5),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_22),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_4),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_281),
.B(n_280),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g328 ( 
.A1(n_313),
.A2(n_316),
.B(n_317),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_320),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_5),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_303),
.B(n_5),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_321),
.B(n_306),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_6),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_322),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_309),
.B1(n_302),
.B2(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_325),
.B(n_326),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_305),
.B1(n_310),
.B2(n_297),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

HB1xp67_ASAP7_75t_SL g333 ( 
.A(n_328),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_324),
.B1(n_7),
.B2(n_8),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_334),
.A2(n_335),
.B(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_315),
.C(n_318),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_314),
.B(n_317),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_329),
.B(n_331),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_340),
.C(n_336),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_339),
.B(n_6),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_8),
.C(n_332),
.Y(n_344)
);


endmodule