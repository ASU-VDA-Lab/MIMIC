module fake_aes_7310_n_19 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_19);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_19;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
BUFx2_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_7), .B(n_6), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
OAI22x1_ASAP7_75t_L g12 ( .A1(n_9), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_13), .B(n_11), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
NOR2x1_ASAP7_75t_L g16 ( .A(n_15), .B(n_10), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_16), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AOI22xp5_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_1), .B1(n_4), .B2(n_5), .Y(n_19) );
endmodule