module fake_netlist_5_1618_n_1228 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1228);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1228;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_268;
wire n_913;
wire n_451;
wire n_523;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_532;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_1222;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_1157;
wire n_998;
wire n_1099;
wire n_841;
wire n_1050;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_1227;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_1128;
wire n_725;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_1203;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_946;
wire n_417;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_933;
wire n_516;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_739;
wire n_508;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_936;
wire n_373;
wire n_820;
wire n_1090;
wire n_757;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_1107;
wire n_1063;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_1104;
wire n_792;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_943;
wire n_524;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_204;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_1214;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_1221;
wire n_654;
wire n_370;
wire n_1172;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_833;
wire n_267;
wire n_570;
wire n_457;
wire n_428;
wire n_514;
wire n_297;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_995;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_1149;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_1225;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_962;
wire n_1219;
wire n_1204;
wire n_1215;
wire n_1216;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_1218;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_1223;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1071;
wire n_1165;
wire n_496;
wire n_1043;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_922;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_974;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_928;
wire n_749;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_197;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_1197;
wire n_1211;
wire n_1226;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_736;
wire n_595;
wire n_502;
wire n_893;
wire n_892;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_630;
wire n_420;
wire n_1202;
wire n_489;
wire n_632;
wire n_699;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_1101;
wire n_1053;
wire n_273;
wire n_1106;
wire n_585;
wire n_349;
wire n_1190;
wire n_1224;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_1116;
wire n_954;
wire n_627;
wire n_1212;
wire n_767;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_1217;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_707;
wire n_795;
wire n_710;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1220;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1072;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_1027;
wire n_490;
wire n_805;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_233;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1207;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_870;
wire n_334;
wire n_599;
wire n_811;
wire n_766;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_868;
wire n_262;
wire n_803;
wire n_666;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_1213;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g179 ( 
.A(n_38),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_165),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_62),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_9),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_81),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_37),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_47),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_29),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_3),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_69),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_0),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_56),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_27),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_37),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_14),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_105),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_23),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_144),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_38),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_91),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_61),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_73),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_90),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_93),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_124),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_41),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_22),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_100),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_28),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_83),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_57),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_104),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_72),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_175),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_64),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_54),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_59),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_114),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_141),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_35),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_110),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_201),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_181),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_186),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_193),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_203),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_207),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_209),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_211),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_212),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_214),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_188),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_243),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_241),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_249),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_251),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_255),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_185),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_258),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_185),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_264),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_265),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_244),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_239),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_261),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_252),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_243),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_271),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_275),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_288),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_302),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_315),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_270),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_269),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_267),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_308),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_272),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_274),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_309),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_309),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_317),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_329),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_337),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_348),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_348),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_346),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_324),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_331),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_331),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_323),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_323),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_324),
.Y(n_380)
);

OAI21x1_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_223),
.B(n_187),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_338),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_338),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_325),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_328),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_328),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_300),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_345),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_358),
.B(n_316),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_292),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_352),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_352),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_318),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_343),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_344),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_347),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_368),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_361),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_390),
.A2(n_362),
.B1(n_360),
.B2(n_327),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_322),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_391),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_371),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_389),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_400),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_363),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_370),
.A2(n_267),
.B1(n_276),
.B2(n_227),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_401),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_401),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_393),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_334),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_399),
.B(n_335),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_370),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_387),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_376),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_392),
.A2(n_355),
.B(n_354),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_335),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_369),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_378),
.B(n_336),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

NOR2x1_ASAP7_75t_L g458 ( 
.A(n_374),
.B(n_276),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_376),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_377),
.B(n_336),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_380),
.B(n_339),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_380),
.B(n_279),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_390),
.A2(n_293),
.B1(n_273),
.B2(n_268),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_390),
.A2(n_293),
.B1(n_273),
.B2(n_292),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_390),
.B(n_281),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_390),
.B(n_285),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_390),
.A2(n_287),
.B1(n_295),
.B2(n_301),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_380),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_381),
.A2(n_356),
.B(n_354),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_370),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_380),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_380),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_380),
.B(n_217),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_373),
.B(n_312),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

BUFx12f_ASAP7_75t_L g493 ( 
.A(n_376),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_390),
.B(n_201),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_217),
.Y(n_497)
);

OA21x2_ASAP7_75t_L g498 ( 
.A1(n_481),
.A2(n_191),
.B(n_190),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_441),
.B(n_351),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_468),
.B(n_190),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_476),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_470),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_191),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_434),
.B(n_282),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_474),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_413),
.B(n_210),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_442),
.A2(n_229),
.B1(n_208),
.B2(n_225),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_421),
.B(n_353),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_413),
.B(n_210),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_480),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_480),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_421),
.B(n_224),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_472),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_208),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_482),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_422),
.B(n_357),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_229),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_481),
.A2(n_236),
.B(n_224),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_484),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_487),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_434),
.B(n_437),
.C(n_449),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_472),
.B(n_236),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_414),
.B(n_206),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_488),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_489),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_422),
.B(n_282),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_435),
.B(n_282),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_467),
.B(n_183),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_424),
.B(n_228),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_472),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_448),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_492),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_495),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_416),
.B(n_222),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_545),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_545),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_505),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_499),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_496),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_535),
.Y(n_554)
);

NOR2x1p5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_442),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_544),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_541),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_511),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_496),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_506),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_509),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_505),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_539),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_R g564 ( 
.A(n_538),
.B(n_448),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_R g565 ( 
.A(n_538),
.B(n_483),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_509),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_522),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_501),
.B(n_424),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_522),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_512),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_501),
.B(n_426),
.Y(n_571)
);

AND3x2_ASAP7_75t_L g572 ( 
.A(n_512),
.B(n_491),
.C(n_465),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_510),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_517),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_517),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_542),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_543),
.B(n_483),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_497),
.B(n_435),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_542),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_542),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_511),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_533),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_543),
.B(n_462),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_533),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_533),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_533),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_553),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_560),
.B(n_502),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_442),
.B1(n_438),
.B2(n_435),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_587),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_558),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_549),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_450),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_553),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_435),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_576),
.B(n_446),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_562),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_559),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_583),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_587),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_583),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_568),
.B(n_435),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_566),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_566),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_556),
.B(n_446),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_573),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_574),
.A2(n_527),
.B(n_498),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_438),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_571),
.B(n_521),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_557),
.B(n_438),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_552),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_574),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_571),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_587),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_581),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_554),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_521),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_555),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_567),
.B(n_438),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_551),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_551),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_572),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_584),
.B(n_543),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_569),
.B(n_438),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_589),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_586),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_564),
.B(n_473),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_550),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_565),
.B(n_447),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_580),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_563),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_585),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_553),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_579),
.B(n_469),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_562),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_562),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_562),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_570),
.A2(n_513),
.B1(n_425),
.B2(n_456),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_579),
.B(n_415),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_579),
.B(n_433),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_579),
.B(n_433),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_581),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_553),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_553),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_579),
.B(n_475),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_553),
.Y(n_662)
);

AO22x1_ASAP7_75t_L g663 ( 
.A1(n_560),
.A2(n_462),
.B1(n_425),
.B2(n_461),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_581),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_568),
.B(n_526),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

NOR2x1p5_ASAP7_75t_L g667 ( 
.A(n_549),
.B(n_493),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_552),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_553),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_562),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_578),
.B(n_502),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_620),
.B(n_419),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_597),
.B(n_490),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_668),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_668),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_613),
.B(n_419),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_664),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_646),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_664),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_590),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_646),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_596),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_629),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_656),
.B(n_425),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_625),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_646),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_657),
.B(n_425),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_631),
.B(n_423),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_596),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_598),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_631),
.B(n_423),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_602),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_633),
.B(n_425),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_600),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_606),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_607),
.Y(n_696)
);

AND2x6_ASAP7_75t_L g697 ( 
.A(n_628),
.B(n_504),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_665),
.B(n_490),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_655),
.A2(n_471),
.B1(n_479),
.B2(n_454),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_622),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_608),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_641),
.A2(n_461),
.B1(n_464),
.B2(n_460),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_608),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_614),
.Y(n_705)
);

CKINVDCx11_ASAP7_75t_R g706 ( 
.A(n_625),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_650),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_630),
.B(n_429),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_658),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_640),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_654),
.B(n_423),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_649),
.B(n_490),
.Y(n_712)
);

BUFx4f_ASAP7_75t_L g713 ( 
.A(n_658),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_634),
.B(n_423),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_648),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_634),
.B(n_423),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_659),
.Y(n_718)
);

AO22x2_ASAP7_75t_L g719 ( 
.A1(n_655),
.A2(n_460),
.B1(n_464),
.B2(n_452),
.Y(n_719)
);

INVx4_ASAP7_75t_SL g720 ( 
.A(n_626),
.Y(n_720)
);

INVx5_ASAP7_75t_L g721 ( 
.A(n_626),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_660),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_650),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_652),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_662),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_649),
.B(n_520),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_634),
.B(n_423),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_652),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_635),
.B(n_436),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_599),
.B(n_485),
.Y(n_730)
);

AO22x2_ASAP7_75t_L g731 ( 
.A1(n_628),
.A2(n_609),
.B1(n_632),
.B2(n_661),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_669),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_612),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_619),
.Y(n_734)
);

INVx6_ASAP7_75t_L g735 ( 
.A(n_601),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_658),
.B(n_637),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_645),
.B(n_485),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

CKINVDCx8_ASAP7_75t_R g739 ( 
.A(n_636),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_667),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_615),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_658),
.B(n_454),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_601),
.Y(n_743)
);

INVx4_ASAP7_75t_SL g744 ( 
.A(n_626),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_609),
.A2(n_454),
.B1(n_440),
.B2(n_494),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_638),
.B(n_504),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_653),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_618),
.Y(n_748)
);

INVx5_ASAP7_75t_L g749 ( 
.A(n_626),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_658),
.B(n_453),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_621),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_621),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_639),
.A2(n_440),
.B1(n_443),
.B2(n_458),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_680),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_702),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_694),
.B(n_455),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_700),
.B(n_637),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_709),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_748),
.B(n_663),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_678),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_690),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_677),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_704),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_736),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_692),
.B(n_661),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_679),
.B(n_642),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_695),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_745),
.B(n_593),
.C(n_478),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_696),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_698),
.B(n_705),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_716),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_736),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_718),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_676),
.B(n_439),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_721),
.B(n_604),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_722),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_725),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_732),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_733),
.B(n_592),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_730),
.B(n_642),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_738),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_721),
.B(n_604),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_679),
.B(n_624),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_673),
.B(n_617),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_741),
.B(n_751),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_746),
.B(n_451),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_752),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_683),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_701),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_731),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_748),
.B(n_627),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_731),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_678),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_683),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_706),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_709),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_719),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_699),
.A2(n_753),
.B1(n_739),
.B2(n_719),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_681),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_746),
.A2(n_477),
.B1(n_647),
.B2(n_591),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_684),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_720),
.B(n_744),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_720),
.B(n_644),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_744),
.B(n_644),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_672),
.B(n_439),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_678),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_709),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_687),
.B(n_591),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_721),
.B(n_749),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_726),
.B(n_592),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_712),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_688),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_746),
.B(n_595),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_697),
.B(n_595),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_697),
.B(n_703),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_724),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_693),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_711),
.A2(n_188),
.B1(n_196),
.B2(n_192),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_749),
.B(n_604),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_750),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_697),
.B(n_603),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_681),
.B(n_671),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_681),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_749),
.B(n_604),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_708),
.B(n_653),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_757),
.A2(n_688),
.B1(n_691),
.B2(n_729),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_768),
.B(n_737),
.C(n_743),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_811),
.B(n_750),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_800),
.B(n_734),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_774),
.B(n_685),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_789),
.B(n_734),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_805),
.B(n_674),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_762),
.B(n_707),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_770),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_784),
.B(n_762),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_L g836 ( 
.A(n_757),
.B(n_463),
.C(n_742),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_756),
.B(n_675),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_803),
.B(n_686),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_803),
.B(n_686),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_773),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_780),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_798),
.A2(n_723),
.B1(n_735),
.B2(n_747),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_786),
.A2(n_432),
.B(n_671),
.C(n_182),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_808),
.A2(n_714),
.B1(n_727),
.B2(n_717),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_804),
.B(n_686),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_770),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_760),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_764),
.B(n_747),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_754),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_761),
.B(n_767),
.Y(n_850)
);

BUFx8_ASAP7_75t_L g851 ( 
.A(n_760),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_769),
.B(n_771),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_788),
.B(n_742),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_798),
.A2(n_182),
.B(n_670),
.C(n_713),
.Y(n_854)
);

NOR2x1_ASAP7_75t_R g855 ( 
.A(n_795),
.B(n_493),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_760),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_784),
.B(n_691),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_777),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_778),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_801),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_801),
.B(n_735),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_804),
.B(n_728),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_808),
.B(n_682),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_776),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_815),
.A2(n_717),
.B1(n_727),
.B2(n_714),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_825),
.B(n_689),
.Y(n_866)
);

O2A1O1Ixp5_ASAP7_75t_L g867 ( 
.A1(n_822),
.A2(n_601),
.B(n_196),
.C(n_233),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_810),
.B(n_670),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_755),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_793),
.B(n_715),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_810),
.B(n_623),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_766),
.B(n_623),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_815),
.A2(n_643),
.B1(n_636),
.B2(n_618),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_797),
.B(n_603),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_818),
.A2(n_643),
.B1(n_465),
.B2(n_451),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_790),
.A2(n_233),
.B(n_230),
.C(n_466),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_792),
.B(n_605),
.Y(n_877)
);

INVxp33_ASAP7_75t_L g878 ( 
.A(n_793),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_816),
.B(n_643),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_772),
.B(n_710),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_793),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_781),
.B(n_605),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_787),
.B(n_651),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_806),
.B(n_710),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_785),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_763),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_806),
.B(n_740),
.Y(n_887)
);

INVx8_ASAP7_75t_L g888 ( 
.A(n_802),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_765),
.B(n_651),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_806),
.B(n_740),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_817),
.A2(n_440),
.B1(n_187),
.B2(n_223),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_766),
.B(n_618),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_794),
.Y(n_893)
);

OAI22xp33_ASAP7_75t_L g894 ( 
.A1(n_759),
.A2(n_466),
.B1(n_452),
.B2(n_459),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_775),
.A2(n_611),
.B(n_604),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_765),
.B(n_618),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_812),
.B(n_444),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_758),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_818),
.B(n_457),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_783),
.B(n_618),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_758),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_759),
.A2(n_618),
.B1(n_440),
.B2(n_520),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_785),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_854),
.A2(n_802),
.B(n_230),
.C(n_809),
.Y(n_904)
);

BUFx4f_ASAP7_75t_L g905 ( 
.A(n_888),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_834),
.B(n_783),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_849),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_851),
.Y(n_908)
);

NOR2x1p5_ASAP7_75t_L g909 ( 
.A(n_836),
.B(n_799),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_846),
.B(n_820),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_831),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_864),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_885),
.B(n_791),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_903),
.Y(n_914)
);

OR2x6_ASAP7_75t_SL g915 ( 
.A(n_835),
.B(n_813),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_860),
.B(n_813),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_850),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_863),
.B(n_444),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_840),
.B(n_779),
.Y(n_919)
);

AO22x1_ASAP7_75t_L g920 ( 
.A1(n_830),
.A2(n_809),
.B1(n_823),
.B2(n_799),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_880),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_850),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_852),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_893),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_868),
.B(n_831),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_SL g926 ( 
.A(n_827),
.B(n_821),
.C(n_814),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_852),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_858),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_859),
.B(n_779),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_899),
.A2(n_759),
.B(n_823),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_829),
.A2(n_876),
.B(n_842),
.Y(n_931)
);

INVx8_ASAP7_75t_L g932 ( 
.A(n_888),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_826),
.A2(n_183),
.B1(n_232),
.B2(n_218),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_894),
.B(n_819),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_873),
.A2(n_824),
.B1(n_819),
.B2(n_821),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_877),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_841),
.B(n_814),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_869),
.B(n_796),
.Y(n_938)
);

AO22x1_ASAP7_75t_L g939 ( 
.A1(n_851),
.A2(n_824),
.B1(n_807),
.B2(n_444),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_888),
.B(n_775),
.Y(n_940)
);

OAI21xp33_ASAP7_75t_SL g941 ( 
.A1(n_884),
.A2(n_453),
.B(n_782),
.Y(n_941)
);

BUFx12f_ASAP7_75t_SL g942 ( 
.A(n_848),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_L g943 ( 
.A(n_861),
.B(n_457),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_828),
.B(n_782),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_828),
.B(n_594),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_SL g946 ( 
.A(n_867),
.B(n_459),
.C(n_445),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_897),
.B(n_443),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_879),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_833),
.B(n_594),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_L g950 ( 
.A(n_843),
.B(n_463),
.C(n_443),
.Y(n_950)
);

OAI221xp5_ASAP7_75t_L g951 ( 
.A1(n_865),
.A2(n_844),
.B1(n_902),
.B2(n_832),
.C(n_837),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_862),
.B(n_184),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_875),
.A2(n_533),
.B1(n_626),
.B2(n_594),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_853),
.B(n_611),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_886),
.B(n_616),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_866),
.B(n_611),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_887),
.B(n_189),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_926),
.B(n_895),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_931),
.B(n_870),
.C(n_890),
.Y(n_959)
);

OAI321xp33_ASAP7_75t_L g960 ( 
.A1(n_934),
.A2(n_896),
.A3(n_877),
.B1(n_874),
.B2(n_889),
.C(n_871),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_920),
.A2(n_930),
.B(n_916),
.C(n_944),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_907),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_932),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_941),
.A2(n_839),
.B(n_838),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_935),
.A2(n_845),
.B(n_857),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_950),
.A2(n_891),
.B(n_197),
.C(n_204),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_912),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_946),
.A2(n_900),
.B(n_892),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_953),
.A2(n_878),
.B1(n_898),
.B2(n_856),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_939),
.A2(n_616),
.B(n_847),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_940),
.B(n_881),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_914),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_911),
.B(n_872),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_925),
.B(n_882),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_L g975 ( 
.A(n_909),
.B(n_901),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_948),
.B(n_855),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_917),
.B(n_882),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_922),
.B(n_883),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_L g979 ( 
.A(n_908),
.B(n_932),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_904),
.A2(n_952),
.B(n_947),
.C(n_951),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_905),
.A2(n_883),
.B(n_901),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_936),
.B(n_901),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_957),
.A2(n_933),
.B(n_918),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_905),
.A2(n_611),
.B(n_548),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_923),
.B(n_533),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_940),
.A2(n_611),
.B(n_534),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_943),
.A2(n_199),
.B(n_216),
.C(n_213),
.Y(n_987)
);

NOR2xp67_ASAP7_75t_L g988 ( 
.A(n_927),
.B(n_1),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_924),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_932),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_942),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_937),
.A2(n_219),
.B(n_221),
.C(n_183),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_910),
.A2(n_913),
.B(n_906),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_906),
.A2(n_929),
.B(n_919),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_915),
.B(n_666),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_938),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_928),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_949),
.B(n_626),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_919),
.A2(n_500),
.B(n_498),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_945),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_929),
.A2(n_183),
.B(n_426),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_956),
.A2(n_235),
.B(n_226),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_955),
.A2(n_540),
.B(n_420),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_921),
.B(n_188),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_954),
.A2(n_428),
.B(n_427),
.Y(n_1005)
);

OAI321xp33_ASAP7_75t_L g1006 ( 
.A1(n_926),
.A2(n_418),
.A3(n_431),
.B1(n_430),
.B2(n_427),
.C(n_428),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_905),
.B(n_218),
.Y(n_1007)
);

INVx11_ASAP7_75t_L g1008 ( 
.A(n_908),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_908),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_931),
.A2(n_540),
.B(n_431),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_905),
.B(n_218),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_931),
.A2(n_430),
.B(n_503),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_931),
.A2(n_540),
.B(n_508),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_905),
.B(n_232),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_911),
.B(n_1),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_993),
.B(n_2),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_994),
.B(n_2),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_974),
.B(n_4),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_983),
.A2(n_518),
.B(n_507),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_1009),
.B(n_4),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_995),
.B(n_5),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_L g1022 ( 
.A(n_1010),
.B(n_417),
.C(n_492),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_SL g1023 ( 
.A1(n_1004),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_991),
.A2(n_519),
.B1(n_546),
.B2(n_529),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_980),
.A2(n_525),
.B(n_523),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_958),
.B(n_232),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_963),
.B(n_6),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_961),
.A2(n_530),
.B(n_528),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_1009),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_989),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1012),
.A2(n_532),
.B(n_524),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_1013),
.A2(n_524),
.B(n_514),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_SL g1033 ( 
.A1(n_1007),
.A2(n_547),
.B(n_537),
.C(n_536),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_964),
.A2(n_524),
.B(n_514),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_959),
.A2(n_514),
.B1(n_516),
.B2(n_515),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_962),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1026),
.A2(n_975),
.B1(n_979),
.B2(n_969),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1016),
.A2(n_988),
.B1(n_992),
.B2(n_1015),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1029),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1017),
.A2(n_1011),
.B1(n_1014),
.B2(n_985),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1034),
.A2(n_1001),
.B(n_960),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_1035),
.B(n_990),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1023),
.A2(n_987),
.B(n_966),
.C(n_1006),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_1021),
.A2(n_982),
.B(n_970),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1029),
.B(n_990),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1036),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1018),
.A2(n_984),
.B(n_968),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_1030),
.A2(n_976),
.B(n_986),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1022),
.A2(n_1000),
.B1(n_965),
.B2(n_990),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1020),
.A2(n_1019),
.B(n_1025),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_SL g1051 ( 
.A1(n_1028),
.A2(n_1002),
.B(n_963),
.C(n_1003),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_1029),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_1027),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_R g1054 ( 
.A(n_1027),
.B(n_1009),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1024),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1031),
.B(n_971),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1032),
.A2(n_981),
.B(n_1005),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1033),
.B(n_1008),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1029),
.B(n_973),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1026),
.A2(n_978),
.B(n_977),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1017),
.B(n_996),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1051),
.A2(n_999),
.B(n_967),
.C(n_972),
.Y(n_1062)
);

BUFx8_ASAP7_75t_SL g1063 ( 
.A(n_1039),
.Y(n_1063)
);

AND2x2_ASAP7_75t_SL g1064 ( 
.A(n_1048),
.B(n_971),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1052),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1046),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_1054),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1053),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1064),
.A2(n_1050),
.B(n_1047),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1068),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1070),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1069),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1070),
.Y(n_1073)
);

BUFx2_ASAP7_75t_R g1074 ( 
.A(n_1072),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1071),
.A2(n_1050),
.B(n_1064),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1073),
.A2(n_1065),
.B(n_1068),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_1075),
.A2(n_1067),
.B1(n_1048),
.B2(n_1038),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_1076),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_1065),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1078),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1080),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1079),
.A2(n_1074),
.B(n_1066),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_1059),
.Y(n_1083)
);

AO21x2_ASAP7_75t_L g1084 ( 
.A1(n_1082),
.A2(n_1045),
.B(n_1042),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_1081),
.B1(n_1058),
.B2(n_1038),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1083),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1084),
.B(n_1062),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_L g1088 ( 
.A1(n_1086),
.A2(n_1084),
.B1(n_1041),
.B2(n_1061),
.C(n_1063),
.Y(n_1088)
);

INVxp67_ASAP7_75t_SL g1089 ( 
.A(n_1087),
.Y(n_1089)
);

INVx5_ASAP7_75t_L g1090 ( 
.A(n_1088),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1088),
.B(n_1055),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1091),
.B(n_1056),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1089),
.B(n_1056),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1090),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1093),
.B(n_1090),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1094),
.B(n_1037),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1095),
.A2(n_1092),
.B1(n_1063),
.B2(n_1057),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_1049),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1098),
.B(n_1040),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_1060),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1100),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1102),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1101),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1103),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1106),
.B(n_7),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_8),
.Y(n_1108)
);

NOR2x1p5_ASAP7_75t_SL g1109 ( 
.A(n_1106),
.B(n_1044),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1109),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1108),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1107),
.Y(n_1112)
);

AO22x2_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_1113)
);

XNOR2x1_ASAP7_75t_L g1114 ( 
.A(n_1112),
.B(n_10),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1114),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1113),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1116),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1115),
.B(n_1111),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1118),
.B(n_996),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1117),
.B(n_996),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1120),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1119),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1122),
.B(n_11),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1121),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1124),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1123),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1124),
.B(n_11),
.Y(n_1127)
);

O2A1O1Ixp5_ASAP7_75t_SL g1128 ( 
.A1(n_1125),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1128)
);

AOI221x1_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.C(n_16),
.Y(n_1129)
);

OAI221xp5_ASAP7_75t_SL g1130 ( 
.A1(n_1127),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1130),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1128),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1132),
.B(n_1129),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1131),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1133),
.B(n_17),
.Y(n_1135)
);

AO21x2_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_18),
.B(n_19),
.Y(n_1136)
);

OAI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1135),
.A2(n_1136),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_19),
.C(n_20),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1137),
.B(n_21),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_SL g1140 ( 
.A(n_1138),
.B(n_24),
.C(n_25),
.Y(n_1140)
);

AOI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1139),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1140),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1142),
.B(n_29),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_L g1144 ( 
.A(n_1141),
.B(n_30),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1142),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1145),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_31),
.Y(n_1147)
);

AO22x2_ASAP7_75t_L g1148 ( 
.A1(n_1143),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1146),
.Y(n_1149)
);

INVxp67_ASAP7_75t_SL g1150 ( 
.A(n_1147),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1149),
.Y(n_1151)
);

NOR4xp25_ASAP7_75t_L g1152 ( 
.A(n_1150),
.B(n_1148),
.C(n_33),
.D(n_34),
.Y(n_1152)
);

NAND2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_32),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_34),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1154),
.A2(n_35),
.B(n_36),
.C(n_39),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1153),
.A2(n_36),
.B(n_39),
.Y(n_1156)
);

NOR4xp25_ASAP7_75t_L g1157 ( 
.A(n_1155),
.B(n_40),
.C(n_41),
.D(n_42),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1156),
.B(n_40),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1158),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1157),
.B(n_42),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1159),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1160),
.B(n_43),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1159),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1161),
.B(n_43),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1163),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_1162),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1166),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1164),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1167),
.A2(n_1165),
.B1(n_45),
.B2(n_46),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1168),
.B(n_44),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1169),
.A2(n_1043),
.B1(n_49),
.B2(n_51),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1170),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1172),
.A2(n_1171),
.B1(n_52),
.B2(n_53),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1172),
.A2(n_48),
.B1(n_55),
.B2(n_58),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1173),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1174),
.Y(n_1176)
);

AOI22x1_ASAP7_75t_L g1177 ( 
.A1(n_1176),
.A2(n_60),
.B1(n_63),
.B2(n_65),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_SL g1178 ( 
.A1(n_1175),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1176),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1178),
.A2(n_76),
.B(n_77),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1177),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1179),
.Y(n_1182)
);

OAI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1177),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1183)
);

AOI221xp5_ASAP7_75t_L g1184 ( 
.A1(n_1182),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.C(n_86),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1181),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1180),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1183),
.Y(n_1187)
);

AOI222xp33_ASAP7_75t_L g1188 ( 
.A1(n_1185),
.A2(n_87),
.B1(n_88),
.B2(n_92),
.C1(n_94),
.C2(n_95),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1186),
.A2(n_96),
.B(n_98),
.Y(n_1189)
);

XNOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1187),
.B(n_99),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_1184),
.A2(n_101),
.B(n_102),
.Y(n_1191)
);

NAND2x1_ASAP7_75t_SL g1192 ( 
.A(n_1185),
.B(n_103),
.Y(n_1192)
);

AOI22x1_ASAP7_75t_L g1193 ( 
.A1(n_1185),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1185),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_1194)
);

OAI222xp33_ASAP7_75t_L g1195 ( 
.A1(n_1185),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.C1(n_118),
.C2(n_119),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1185),
.A2(n_997),
.B1(n_121),
.B2(n_122),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1185),
.A2(n_120),
.B(n_123),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1185),
.B(n_125),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1185),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_1199)
);

AOI221xp5_ASAP7_75t_L g1200 ( 
.A1(n_1191),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.C(n_132),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1190),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1192),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1198),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1197),
.A2(n_142),
.B(n_143),
.Y(n_1204)
);

XNOR2xp5_ASAP7_75t_L g1205 ( 
.A(n_1193),
.B(n_145),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1196),
.A2(n_146),
.B(n_147),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1189),
.Y(n_1207)
);

XNOR2xp5_ASAP7_75t_L g1208 ( 
.A(n_1194),
.B(n_148),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1207),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1203),
.A2(n_1199),
.B1(n_1188),
.B2(n_1195),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1205),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1208),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1206),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1204),
.Y(n_1214)
);

XNOR2x2_ASAP7_75t_L g1215 ( 
.A(n_1200),
.B(n_149),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1201),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1209),
.A2(n_1210),
.B(n_1213),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_SL g1218 ( 
.A1(n_1216),
.A2(n_1202),
.B1(n_151),
.B2(n_153),
.Y(n_1218)
);

AOI222xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1212),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.C1(n_157),
.C2(n_158),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1217),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1220),
.A2(n_1214),
.B1(n_1211),
.B2(n_1215),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1221),
.Y(n_1222)
);

AO21x2_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1218),
.B(n_1219),
.Y(n_1223)
);

OAI221xp5_ASAP7_75t_R g1224 ( 
.A1(n_1223),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.C(n_162),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1224),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1225),
.A2(n_171),
.B(n_173),
.Y(n_1226)
);

AOI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1226),
.A2(n_174),
.B(n_176),
.C(n_177),
.Y(n_1227)
);

AOI211xp5_ASAP7_75t_L g1228 ( 
.A1(n_1227),
.A2(n_178),
.B(n_998),
.C(n_997),
.Y(n_1228)
);


endmodule