module fake_ariane_891_n_163 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_163);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_163;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_124;
wire n_119;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_19;
wire n_40;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_21;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_121;
wire n_93;
wire n_118;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_22;
wire n_43;
wire n_87;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVxp33_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_7),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_20),
.A2(n_15),
.B1(n_23),
.B2(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_31),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_44),
.B(n_45),
.C(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_36),
.B(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_50),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_45),
.B(n_37),
.Y(n_62)
);

AOI21x1_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_48),
.B(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_43),
.B(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_43),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_43),
.B(n_46),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_35),
.B(n_41),
.C(n_47),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_43),
.B(n_40),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_48),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_43),
.B(n_41),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_46),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_38),
.B(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_65),
.B(n_68),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_49),
.Y(n_90)
);

AOI21x1_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_66),
.B(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

AO31x2_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_60),
.A3(n_56),
.B(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_92),
.Y(n_99)
);

OAI221xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_49),
.B1(n_73),
.B2(n_76),
.C(n_79),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_82),
.B(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_71),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_60),
.B1(n_75),
.B2(n_88),
.C(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_89),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_86),
.C(n_91),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_91),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_86),
.Y(n_112)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_106),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_95),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_104),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_103),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_74),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_128),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_126),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_122),
.B1(n_120),
.B2(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

CKINVDCx6p67_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_115),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_123),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_125),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_131),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_139),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_135),
.Y(n_149)
);

OAI211xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_134),
.B(n_136),
.C(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_141),
.B1(n_144),
.B2(n_143),
.C(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_148),
.B(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_132),
.B1(n_144),
.B2(n_139),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_132),
.B1(n_143),
.B2(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_158),
.B(n_154),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_158),
.B1(n_147),
.B2(n_135),
.C(n_149),
.Y(n_163)
);


endmodule