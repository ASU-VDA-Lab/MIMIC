module fake_jpeg_25522_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_44),
.Y(n_59)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_32),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_32),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_17),
.B1(n_16),
.B2(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_71),
.B1(n_75),
.B2(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_35),
.Y(n_101)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_37),
.A2(n_17),
.B1(n_16),
.B2(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_24),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_41),
.Y(n_115)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_43),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_39),
.A2(n_17),
.B1(n_16),
.B2(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_21),
.B1(n_18),
.B2(n_31),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_78),
.A2(n_92),
.B1(n_113),
.B2(n_33),
.Y(n_145)
);

OA22x2_ASAP7_75t_SL g79 ( 
.A1(n_73),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_81),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_19),
.B1(n_18),
.B2(n_24),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_80),
.A2(n_98),
.B1(n_33),
.B2(n_30),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_90),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_105),
.B1(n_54),
.B2(n_74),
.Y(n_131)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_86),
.Y(n_128)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_46),
.B1(n_26),
.B2(n_27),
.Y(n_92)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_96),
.Y(n_142)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_25),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_59),
.B1(n_72),
.B2(n_64),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_63),
.B(n_15),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_35),
.B1(n_46),
.B2(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_107),
.Y(n_141)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_115),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_42),
.C(n_36),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_40),
.C(n_23),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_47),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_60),
.B1(n_29),
.B2(n_30),
.Y(n_134)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_55),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_42),
.B1(n_40),
.B2(n_47),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_60),
.B1(n_33),
.B2(n_30),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_70),
.B(n_1),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_144),
.B(n_111),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_25),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_23),
.C(n_104),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_134),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_133),
.B1(n_145),
.B2(n_107),
.Y(n_150)
);

OAI22x1_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_25),
.B1(n_29),
.B2(n_20),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_93),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_137),
.B1(n_108),
.B2(n_76),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_79),
.A2(n_20),
.B1(n_30),
.B2(n_23),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_29),
.B(n_33),
.C(n_23),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_84),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_146),
.A2(n_86),
.B1(n_82),
.B2(n_96),
.Y(n_159)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_94),
.A3(n_115),
.B1(n_110),
.B2(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_148),
.B(n_149),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_89),
.B(n_111),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_151),
.B(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_83),
.B1(n_112),
.B2(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_83),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_153),
.B(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_14),
.C(n_13),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_100),
.C(n_91),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_123),
.B(n_138),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_87),
.B1(n_90),
.B2(n_95),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_172),
.B1(n_0),
.B2(n_4),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_124),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_100),
.B1(n_106),
.B2(n_99),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_167),
.B1(n_174),
.B2(n_134),
.Y(n_181)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_165),
.B(n_170),
.Y(n_208)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_136),
.B1(n_144),
.B2(n_130),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_132),
.C(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_114),
.B1(n_99),
.B2(n_102),
.Y(n_172)
);

AOI22x1_ASAP7_75t_SL g173 ( 
.A1(n_125),
.A2(n_14),
.B1(n_12),
.B2(n_2),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_0),
.C(n_1),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_179),
.C(n_127),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_120),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_10),
.C(n_3),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_181),
.B(n_200),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_138),
.B(n_118),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_205),
.B(n_206),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_149),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_193),
.C(n_207),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_195),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_191),
.B(n_196),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_124),
.B(n_127),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_178),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_168),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

AO22x1_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_132),
.B1(n_135),
.B2(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_141),
.B1(n_143),
.B2(n_126),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_202),
.B1(n_156),
.B2(n_164),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_154),
.A2(n_141),
.B1(n_126),
.B2(n_116),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_0),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_4),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_9),
.B(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_218),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_223),
.B1(n_224),
.B2(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_225),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_178),
.B(n_165),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_227),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_175),
.B1(n_161),
.B2(n_147),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_151),
.B1(n_174),
.B2(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_188),
.A2(n_171),
.B1(n_166),
.B2(n_179),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_236),
.B1(n_211),
.B2(n_203),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_186),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_229),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_194),
.A3(n_191),
.B1(n_190),
.B2(n_209),
.C1(n_181),
.C2(n_185),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_238),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_4),
.C(n_5),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_183),
.C(n_8),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_234)
);

OAI22x1_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_207),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_184),
.A2(n_9),
.B(n_7),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_202),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_211),
.A2(n_8),
.B1(n_9),
.B2(n_196),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_180),
.B1(n_198),
.B2(n_183),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_213),
.B1(n_225),
.B2(n_221),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_180),
.B1(n_204),
.B2(n_201),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_213),
.B1(n_216),
.B2(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_254),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_248),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_252),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_187),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_260),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_8),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_214),
.B(n_8),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_222),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_269),
.B1(n_277),
.B2(n_232),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_220),
.C(n_235),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_260),
.C(n_261),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_235),
.B1(n_219),
.B2(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_230),
.B1(n_223),
.B2(n_236),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_262),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_287),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_250),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_298),
.C(n_259),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_255),
.B1(n_215),
.B2(n_236),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_292),
.B1(n_224),
.B2(n_248),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_255),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_215),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_252),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_279),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_238),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_263),
.C(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_306),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_273),
.B1(n_263),
.B2(n_267),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_300),
.A2(n_302),
.B1(n_310),
.B2(n_240),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_307),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_257),
.B(n_246),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_282),
.B1(n_278),
.B2(n_265),
.Y(n_304)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_276),
.B(n_274),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_277),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_288),
.C(n_297),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_291),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_315),
.C(n_319),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_292),
.B1(n_284),
.B2(n_271),
.Y(n_314)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_276),
.C(n_267),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_303),
.C(n_301),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_270),
.B1(n_275),
.B2(n_290),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_316),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_325),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_300),
.B1(n_295),
.B2(n_234),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_254),
.B(n_237),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_314),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_321),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_312),
.C(n_323),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_331),
.B(n_333),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_329),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_327),
.B(n_319),
.Y(n_339)
);


endmodule