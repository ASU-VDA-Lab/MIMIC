module fake_jpeg_9493_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_69),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_29),
.B1(n_22),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_66),
.B1(n_16),
.B2(n_17),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_29),
.B1(n_31),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_16),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_17),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_31),
.B1(n_18),
.B2(n_24),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_16),
.Y(n_94)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_78),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_31),
.B1(n_17),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_76),
.A2(n_86),
.B1(n_98),
.B2(n_105),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_42),
.C(n_45),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_83),
.C(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_106),
.B1(n_19),
.B2(n_23),
.Y(n_116)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_82),
.B(n_84),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_34),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_34),
.C(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_88),
.B(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_91),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_27),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_35),
.B1(n_32),
.B2(n_19),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_68),
.B1(n_26),
.B2(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_28),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_61),
.Y(n_138)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_104),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_35),
.B1(n_32),
.B2(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_19),
.B(n_23),
.C(n_69),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_112),
.A2(n_120),
.B1(n_126),
.B2(n_135),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_114),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_120),
.C(n_141),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_49),
.C(n_52),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_132),
.C(n_100),
.Y(n_171)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_77),
.A2(n_63),
.B1(n_61),
.B2(n_58),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_25),
.B1(n_33),
.B2(n_58),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_80),
.C(n_74),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_75),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_63),
.B1(n_61),
.B2(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_74),
.A2(n_25),
.B1(n_33),
.B2(n_57),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_97),
.B1(n_78),
.B2(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_94),
.B(n_81),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_142),
.A2(n_148),
.B(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_75),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_153),
.C(n_171),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_151),
.Y(n_175)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_154),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_99),
.B(n_87),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_125),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_162),
.B1(n_169),
.B2(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_84),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_109),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx10_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_88),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_165),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_89),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_25),
.B(n_34),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_108),
.B1(n_97),
.B2(n_73),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_127),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_85),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_9),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_10),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_132),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_184),
.C(n_194),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_190),
.Y(n_213)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_137),
.A3(n_114),
.B1(n_116),
.B2(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_126),
.B1(n_119),
.B2(n_124),
.Y(n_182)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_119),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_144),
.B(n_174),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_124),
.C(n_111),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_186),
.B(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_195),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_139),
.B1(n_121),
.B2(n_25),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_198),
.B1(n_207),
.B2(n_172),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_197),
.B1(n_199),
.B2(n_204),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_117),
.C(n_8),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_208),
.B(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_202),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_202),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_215),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_212),
.A2(n_225),
.B(n_226),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_173),
.B1(n_163),
.B2(n_148),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_214),
.A2(n_235),
.B(n_189),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_187),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_231),
.C(n_234),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_160),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_218),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_180),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_230),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_183),
.A2(n_154),
.B1(n_149),
.B2(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_149),
.B1(n_164),
.B2(n_147),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_R g250 ( 
.A1(n_233),
.A2(n_198),
.B(n_207),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_166),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_147),
.B(n_117),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_200),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_249),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_248),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_198),
.B(n_184),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_201),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_177),
.B1(n_199),
.B2(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_179),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_236),
.B1(n_252),
.B2(n_242),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_194),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_257),
.B1(n_258),
.B2(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_195),
.C(n_203),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_216),
.C(n_235),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_209),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_256),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_227),
.A2(n_188),
.B1(n_205),
.B2(n_201),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_221),
.B1(n_218),
.B2(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_272),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_223),
.B1(n_226),
.B2(n_233),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_262),
.B1(n_267),
.B2(n_270),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_265),
.B(n_269),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_222),
.B1(n_212),
.B2(n_217),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_205),
.B1(n_213),
.B2(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_238),
.B(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_276),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_249),
.C(n_237),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_7),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_277),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_243),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_254),
.B(n_9),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_0),
.C(n_3),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_0),
.C(n_3),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_15),
.C(n_4),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_284),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_239),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_286),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_243),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_251),
.Y(n_290)
);

AOI32xp33_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_266),
.A3(n_263),
.B1(n_259),
.B2(n_261),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_244),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_251),
.Y(n_293)
);

NAND4xp25_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.C(n_11),
.D(n_14),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_255),
.C(n_256),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_297),
.A2(n_282),
.B1(n_280),
.B2(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_274),
.B(n_255),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_300),
.Y(n_314)
);

AO221x1_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_260),
.B1(n_9),
.B2(n_13),
.C(n_6),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_272),
.B(n_268),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_11),
.B(n_14),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_304),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_5),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_285),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_15),
.B(n_4),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_3),
.B(n_5),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_306),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_281),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_301),
.C(n_300),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_5),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_317),
.A2(n_298),
.B(n_5),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_324),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_295),
.B(n_314),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_295),
.C(n_315),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_327),
.A2(n_328),
.B(n_315),
.Y(n_330)
);

INVx11_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_319),
.B(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_328),
.B1(n_326),
.B2(n_325),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_318),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_310),
.Y(n_334)
);


endmodule