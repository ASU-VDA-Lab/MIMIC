module fake_netlist_5_1342_n_1887 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1887);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1887;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_81),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_117),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_84),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_171),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_133),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_26),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_49),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_91),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_43),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_46),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_51),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_54),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_63),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_47),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_40),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_15),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_116),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_42),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_172),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_8),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_37),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_45),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_13),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_44),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_50),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_62),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_103),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_60),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_104),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_132),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_85),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_69),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_118),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_18),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_152),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_72),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_174),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_114),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_71),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_181),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_12),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_65),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_28),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_48),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_45),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_124),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_162),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_56),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_173),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_60),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_110),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_49),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_44),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_107),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_139),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_178),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_182),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_66),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_54),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_86),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_137),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_95),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_144),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_68),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_159),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_156),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_122),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_18),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_64),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_50),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_74),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_128),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_90),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_29),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_43),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_92),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_20),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_96),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_180),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_150),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_113),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_19),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_64),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_8),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_21),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_123),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_76),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_17),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_20),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_99),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_108),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_102),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_88),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_129),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_28),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_30),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_130),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_52),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_134),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_77),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_46),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_35),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_177),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_57),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_16),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_89),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_109),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_37),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_19),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_125),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_98),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_40),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_93),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_5),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_168),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_73),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_155),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_4),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_34),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_14),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_1),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_14),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_32),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_120),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_26),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_184),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_1),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_67),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_100),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_94),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_146),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_5),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_131),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_0),
.Y(n_364)
);

CKINVDCx11_ASAP7_75t_R g365 ( 
.A(n_52),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_32),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_31),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_365),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_224),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_235),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_265),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_229),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_185),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_244),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_216),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_220),
.B(n_269),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_211),
.B(n_0),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_245),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_186),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_191),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_246),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_248),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_265),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_284),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_265),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_254),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_211),
.B(n_3),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_265),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_265),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_189),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_276),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_260),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_276),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_276),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_247),
.B(n_3),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_262),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_276),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_267),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_194),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_276),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_268),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_296),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_191),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_247),
.B(n_6),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_189),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_274),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_279),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_281),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_270),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_282),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_285),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_296),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_288),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_186),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_359),
.B(n_6),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_291),
.Y(n_417)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_286),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_249),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_247),
.B(n_9),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_219),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_296),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_293),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_296),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_296),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_319),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_347),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_298),
.B(n_9),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_303),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_297),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_303),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_249),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_298),
.B(n_10),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_200),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_299),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_303),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_238),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_303),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_303),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_257),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_255),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_326),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_222),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_358),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_306),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_222),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_L g448 ( 
.A(n_298),
.B(n_10),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_227),
.B(n_11),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_307),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_240),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_240),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_233),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_201),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_309),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_250),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_250),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_263),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_201),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_189),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_369),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_370),
.B(n_320),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_189),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_460),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_397),
.B(n_187),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_437),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_374),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_378),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_390),
.A2(n_256),
.B(n_227),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_187),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_421),
.B(n_188),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_380),
.B(n_255),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_371),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_381),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_371),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_383),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_403),
.B(n_256),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_382),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_386),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_385),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_392),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_429),
.B(n_188),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_420),
.B(n_316),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_438),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_373),
.Y(n_496)
);

OA21x2_ASAP7_75t_L g497 ( 
.A1(n_405),
.A2(n_292),
.B(n_263),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_460),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_433),
.B(n_442),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_460),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_399),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_460),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_391),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_396),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_393),
.Y(n_509)
);

NAND2x1p5_ASAP7_75t_L g510 ( 
.A(n_395),
.B(n_189),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_409),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_434),
.B(n_190),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_398),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_376),
.B(n_243),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_R g515 ( 
.A(n_446),
.B(n_356),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_377),
.B(n_190),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_394),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_394),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_401),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_406),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_400),
.Y(n_522)
);

CKINVDCx8_ASAP7_75t_R g523 ( 
.A(n_368),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_400),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_402),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_407),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_SL g531 ( 
.A(n_372),
.B(n_202),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g532 ( 
.A(n_408),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_423),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_410),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_425),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_519),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_316),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_517),
.B(n_411),
.Y(n_541)
);

AOI22x1_ASAP7_75t_L g542 ( 
.A1(n_510),
.A2(n_375),
.B1(n_494),
.B2(n_483),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_412),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_472),
.A2(n_387),
.B1(n_454),
.B2(n_379),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_503),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_500),
.B(n_395),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_465),
.B(n_414),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_500),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_467),
.B(n_417),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_517),
.B(n_431),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_519),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_466),
.B(n_384),
.Y(n_554)
);

BUFx6f_ASAP7_75t_SL g555 ( 
.A(n_503),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_514),
.B(n_436),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_L g557 ( 
.A1(n_472),
.A2(n_350),
.B1(n_308),
.B2(n_353),
.Y(n_557)
);

NAND2x1p5_ASAP7_75t_L g558 ( 
.A(n_500),
.B(n_192),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_473),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_490),
.B(n_450),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_473),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_466),
.B(n_418),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_490),
.A2(n_455),
.B1(n_416),
.B2(n_404),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_512),
.B(n_471),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_532),
.B(n_404),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_534),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_512),
.B(n_471),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_515),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_534),
.Y(n_569)
);

AND2x2_ASAP7_75t_SL g570 ( 
.A(n_483),
.B(n_449),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_462),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_530),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_507),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_494),
.B(n_448),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_534),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_469),
.Y(n_578)
);

BUFx4f_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_494),
.B(n_474),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_474),
.B(n_448),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_510),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_473),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_474),
.B(n_444),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_475),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_496),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_530),
.B(n_426),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_510),
.B(n_333),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_510),
.B(n_290),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_462),
.B(n_333),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_530),
.B(n_475),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_476),
.B(n_290),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_478),
.B(n_458),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_480),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_464),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_486),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_484),
.B(n_290),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_485),
.A2(n_441),
.B1(n_445),
.B2(n_443),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_497),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_480),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_482),
.B(n_426),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_482),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_489),
.B(n_422),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_507),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_488),
.B(n_444),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_488),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_491),
.B(n_458),
.Y(n_610)
);

BUFx8_ASAP7_75t_SL g611 ( 
.A(n_486),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_481),
.B(n_261),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_508),
.B(n_290),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_493),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_493),
.B(n_498),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_498),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_531),
.A2(n_353),
.B1(n_419),
.B2(n_424),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_502),
.B(n_430),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_505),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_513),
.B(n_453),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_464),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_497),
.A2(n_292),
.B1(n_237),
.B2(n_332),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_509),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_481),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_520),
.B(n_290),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_526),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_497),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_509),
.B(n_457),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_516),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_521),
.B(n_427),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_518),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_522),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_507),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_507),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_527),
.B(n_428),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_464),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_522),
.B(n_430),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_507),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_524),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_525),
.B(n_447),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_528),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_528),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_529),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_529),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_507),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_533),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_526),
.B(n_193),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_536),
.Y(n_654)
);

BUFx4f_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_536),
.B(n_432),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_464),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_537),
.B(n_321),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_532),
.A2(n_205),
.B1(n_212),
.B2(n_209),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_463),
.Y(n_661)
);

INVxp33_ASAP7_75t_L g662 ( 
.A(n_537),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_463),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_470),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_470),
.B(n_432),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_499),
.B(n_439),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_499),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_499),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_463),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_470),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_463),
.A2(n_311),
.B1(n_313),
.B2(n_317),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_532),
.B(n_193),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_523),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_504),
.B(n_440),
.Y(n_676)
);

NOR2x1p5_ASAP7_75t_L g677 ( 
.A(n_523),
.B(n_202),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_504),
.B(n_321),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_506),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_506),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_506),
.B(n_440),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_479),
.B(n_195),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_463),
.Y(n_683)
);

AND2x2_ASAP7_75t_SL g684 ( 
.A(n_495),
.B(n_321),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_487),
.B(n_203),
.Y(n_686)
);

AND2x6_ASAP7_75t_SL g687 ( 
.A(n_674),
.B(n_339),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_562),
.B(n_495),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_564),
.B(n_567),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_606),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_541),
.A2(n_305),
.B(n_302),
.C(n_289),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_545),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_580),
.B(n_196),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_552),
.B(n_204),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_580),
.B(n_196),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_562),
.B(n_197),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_543),
.B(n_197),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_621),
.B(n_198),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_585),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_582),
.B(n_207),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_560),
.B(n_223),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_579),
.A2(n_492),
.B(n_487),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_684),
.B(n_198),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_599),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_547),
.B(n_199),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_684),
.B(n_199),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_685),
.B(n_351),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_549),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_570),
.B(n_225),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_550),
.B(n_554),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_570),
.B(n_232),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_626),
.B(n_242),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_577),
.B(n_321),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_626),
.B(n_242),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_554),
.B(n_205),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_596),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_584),
.B(n_242),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_548),
.B(n_209),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_572),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_661),
.B(n_253),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_586),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_596),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_597),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_579),
.A2(n_672),
.B(n_664),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_595),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_558),
.A2(n_624),
.B1(n_546),
.B2(n_542),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_595),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_546),
.B(n_212),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_608),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_597),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_577),
.B(n_321),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_575),
.B(n_258),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_577),
.B(n_602),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_584),
.B(n_312),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_575),
.B(n_259),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_558),
.B(n_322),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_581),
.B(n_322),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_581),
.B(n_272),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_577),
.B(n_354),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_629),
.B(n_278),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_540),
.A2(n_336),
.B1(n_346),
.B2(n_360),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_540),
.A2(n_331),
.B1(n_361),
.B2(n_328),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_629),
.B(n_540),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_540),
.A2(n_329),
.B1(n_343),
.B2(n_283),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_625),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_608),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_571),
.B(n_312),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_625),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_629),
.B(n_540),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_652),
.B(n_312),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_557),
.B(n_239),
.C(n_241),
.Y(n_751)
);

NAND2x1_ASAP7_75t_L g752 ( 
.A(n_561),
.B(n_661),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_540),
.B(n_492),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_594),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_568),
.B(n_535),
.Y(n_755)
);

BUFx8_ASAP7_75t_L g756 ( 
.A(n_555),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_577),
.B(n_492),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_602),
.B(n_354),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_662),
.B(n_323),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_602),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_563),
.A2(n_352),
.B(n_366),
.C(n_362),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_602),
.B(n_501),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_602),
.B(n_501),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_610),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_665),
.A2(n_354),
.B1(n_364),
.B2(n_243),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_592),
.B(n_501),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_632),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_568),
.B(n_323),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_593),
.B(n_463),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_578),
.B(n_337),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_681),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_603),
.B(n_463),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_556),
.A2(n_337),
.B1(n_363),
.B2(n_340),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_605),
.B(n_463),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_665),
.A2(n_354),
.B1(n_243),
.B2(n_315),
.Y(n_775)
);

BUFx6f_ASAP7_75t_SL g776 ( 
.A(n_539),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_665),
.A2(n_354),
.B1(n_315),
.B2(n_463),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_609),
.B(n_340),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_614),
.B(n_341),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_544),
.B(n_341),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_662),
.B(n_345),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_632),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_610),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_594),
.B(n_345),
.Y(n_784)
);

AOI22x1_ASAP7_75t_L g785 ( 
.A1(n_664),
.A2(n_363),
.B1(n_217),
.B2(n_208),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_600),
.B(n_315),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_579),
.B(n_661),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_660),
.Y(n_788)
);

INVx8_ASAP7_75t_L g789 ( 
.A(n_565),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_615),
.B(n_221),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_590),
.A2(n_264),
.B1(n_266),
.B2(n_310),
.Y(n_791)
);

AND2x2_ASAP7_75t_SL g792 ( 
.A(n_589),
.B(n_447),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_617),
.B(n_226),
.Y(n_793)
);

BUFx5_ASAP7_75t_L g794 ( 
.A(n_683),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_630),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_228),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_590),
.A2(n_300),
.B1(n_230),
.B2(n_231),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_631),
.B(n_234),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_633),
.B(n_236),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_644),
.B(n_251),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_L g801 ( 
.A(n_613),
.B(n_314),
.C(n_252),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_628),
.B(n_367),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_630),
.Y(n_803)
);

INVx8_ASAP7_75t_L g804 ( 
.A(n_565),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_645),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_645),
.B(n_451),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_681),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_539),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_646),
.B(n_271),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_647),
.B(n_273),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_663),
.B(n_275),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_649),
.B(n_277),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_663),
.B(n_280),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_620),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_539),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_622),
.A2(n_591),
.B1(n_654),
.B2(n_651),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_653),
.B(n_294),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_663),
.B(n_295),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_669),
.B(n_301),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_587),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_559),
.B(n_304),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_635),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_635),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_559),
.B(n_574),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_636),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_559),
.B(n_318),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_636),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_613),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_627),
.B(n_344),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_627),
.B(n_348),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_643),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_612),
.B(n_206),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_643),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_648),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_648),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_669),
.B(n_683),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_574),
.B(n_349),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_355),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_616),
.B(n_357),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_555),
.B(n_206),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_669),
.B(n_208),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_672),
.A2(n_588),
.B(n_668),
.C(n_667),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_681),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_574),
.B(n_457),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_565),
.A2(n_330),
.B1(n_214),
.B2(n_215),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_583),
.B(n_456),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_680),
.B(n_456),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_538),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_683),
.B(n_327),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_555),
.B(n_210),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_588),
.A2(n_680),
.B1(n_551),
.B2(n_538),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_677),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_565),
.A2(n_325),
.B1(n_210),
.B2(n_327),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_689),
.B(n_583),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_689),
.B(n_583),
.Y(n_855)
);

O2A1O1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_709),
.A2(n_658),
.B(n_589),
.C(n_656),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_710),
.B(n_690),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_843),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_843),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_710),
.B(n_598),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_711),
.A2(n_618),
.B1(n_639),
.B2(n_634),
.Y(n_861)
);

AOI22x1_ASAP7_75t_L g862 ( 
.A1(n_820),
.A2(n_667),
.B1(n_640),
.B2(n_657),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_743),
.A2(n_561),
.B1(n_673),
.B2(n_667),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_726),
.A2(n_612),
.B1(n_658),
.B2(n_678),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_718),
.B(n_598),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_728),
.A2(n_640),
.B(n_657),
.C(n_598),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_694),
.B(n_660),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_725),
.A2(n_678),
.B1(n_367),
.B2(n_566),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_761),
.A2(n_604),
.B(n_619),
.C(n_641),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_713),
.A2(n_739),
.B(n_731),
.Y(n_870)
);

AOI21xp33_ASAP7_75t_L g871 ( 
.A1(n_838),
.A2(n_601),
.B(n_215),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_847),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_718),
.B(n_640),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_693),
.A2(n_686),
.B(n_682),
.C(n_666),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_749),
.A2(n_561),
.B1(n_657),
.B2(n_671),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_847),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_704),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_696),
.B(n_214),
.C(n_217),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_697),
.B(n_679),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_754),
.A2(n_828),
.B1(n_733),
.B2(n_760),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_713),
.A2(n_676),
.B(n_573),
.Y(n_882)
);

AO21x1_ASAP7_75t_L g883 ( 
.A1(n_731),
.A2(n_573),
.B(n_607),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_760),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_752),
.A2(n_655),
.B(n_573),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_739),
.A2(n_576),
.B(n_551),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_771),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_760),
.Y(n_888)
);

AO32x1_ASAP7_75t_L g889 ( 
.A1(n_816),
.A2(n_569),
.A3(n_553),
.B1(n_566),
.B2(n_576),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_824),
.A2(n_655),
.B(n_642),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_697),
.A2(n_561),
.B1(n_675),
.B2(n_660),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_814),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_808),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_688),
.B(n_218),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_760),
.B(n_675),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_728),
.A2(n_553),
.B(n_569),
.C(n_670),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_705),
.A2(n_675),
.B1(n_607),
.B2(n_642),
.Y(n_897)
);

AND2x6_ASAP7_75t_L g898 ( 
.A(n_757),
.B(n_638),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_771),
.B(n_607),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_733),
.A2(n_642),
.B(n_650),
.Y(n_900)
);

OAI21xp33_ASAP7_75t_L g901 ( 
.A1(n_715),
.A2(n_342),
.B(n_324),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_762),
.A2(n_650),
.B(n_638),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_788),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_758),
.A2(n_670),
.B(n_451),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_696),
.B(n_338),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_721),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_695),
.A2(n_841),
.B(n_738),
.C(n_735),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_770),
.B(n_650),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_776),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_763),
.A2(n_650),
.B(n_638),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_727),
.A2(n_338),
.B1(n_330),
.B2(n_334),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_729),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_839),
.B(n_638),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_701),
.B(n_637),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_807),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_746),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_715),
.B(n_452),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_841),
.A2(n_324),
.B(n_334),
.C(n_335),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_755),
.B(n_335),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_737),
.A2(n_637),
.B1(n_342),
.B2(n_611),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_717),
.B(n_11),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_740),
.A2(n_176),
.B1(n_167),
.B2(n_165),
.Y(n_922)
);

NAND3xp33_ASAP7_75t_L g923 ( 
.A(n_773),
.B(n_838),
.C(n_781),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_787),
.A2(n_161),
.B(n_160),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_807),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_737),
.B(n_611),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_787),
.A2(n_158),
.B(n_154),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_836),
.A2(n_149),
.B(n_147),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_734),
.B(n_21),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_700),
.A2(n_145),
.B1(n_143),
.B2(n_140),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_699),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_699),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_759),
.B(n_22),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_736),
.B(n_136),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_836),
.A2(n_126),
.B(n_119),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_724),
.A2(n_101),
.B(n_87),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_712),
.B(n_22),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_753),
.A2(n_83),
.B(n_80),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_764),
.B(n_24),
.Y(n_939)
);

BUFx4f_ASAP7_75t_L g940 ( 
.A(n_789),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_842),
.A2(n_78),
.B(n_25),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_714),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_702),
.A2(n_24),
.B(n_25),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_776),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_783),
.B(n_27),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_795),
.B(n_803),
.Y(n_946)
);

O2A1O1Ixp5_ASAP7_75t_L g947 ( 
.A1(n_732),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_947)
);

NAND2xp33_ASAP7_75t_L g948 ( 
.A(n_794),
.B(n_31),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_716),
.A2(n_33),
.B(n_36),
.C(n_38),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_806),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_844),
.A2(n_36),
.B(n_38),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_805),
.B(n_39),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_750),
.B(n_692),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_811),
.A2(n_39),
.B(n_41),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_765),
.A2(n_62),
.B1(n_53),
.B2(n_55),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_708),
.B(n_719),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_806),
.B(n_48),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_722),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_789),
.Y(n_959)
);

AO32x2_ASAP7_75t_L g960 ( 
.A1(n_797),
.A2(n_53),
.A3(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_791),
.A2(n_58),
.B(n_59),
.Y(n_961)
);

OAI22xp33_ASAP7_75t_L g962 ( 
.A1(n_832),
.A2(n_59),
.B1(n_61),
.B2(n_853),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_722),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_806),
.B(n_61),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_821),
.B(n_826),
.Y(n_965)
);

OAI321xp33_ASAP7_75t_L g966 ( 
.A1(n_829),
.A2(n_775),
.A3(n_845),
.B1(n_736),
.B2(n_703),
.C(n_706),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_837),
.B(n_829),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_723),
.Y(n_968)
);

OAI21xp33_ASAP7_75t_L g969 ( 
.A1(n_747),
.A2(n_802),
.B(n_751),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_723),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_815),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_801),
.A2(n_822),
.B(n_834),
.C(n_850),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_840),
.A2(n_850),
.B(n_825),
.C(n_827),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_846),
.A2(n_720),
.B(n_811),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_851),
.A2(n_848),
.B(n_833),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_698),
.B(n_799),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_819),
.B(n_818),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_720),
.A2(n_819),
.B(n_818),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_813),
.A2(n_774),
.B(n_772),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_768),
.B(n_840),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_780),
.A2(n_784),
.B(n_786),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_756),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_769),
.A2(n_766),
.B(n_827),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_792),
.B(n_782),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_707),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_730),
.B(n_835),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_SL g987 ( 
.A1(n_691),
.A2(n_849),
.B(n_830),
.C(n_778),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_794),
.B(n_790),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_794),
.B(n_796),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_849),
.A2(n_798),
.B(n_800),
.C(n_809),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_730),
.A2(n_748),
.B(n_833),
.C(n_831),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_810),
.A2(n_812),
.B(n_817),
.C(n_793),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_745),
.A2(n_782),
.B(n_823),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_779),
.B(n_785),
.C(n_852),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_794),
.B(n_777),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_741),
.A2(n_744),
.B1(n_742),
.B2(n_835),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_848),
.A2(n_767),
.B(n_823),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_707),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_707),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_745),
.A2(n_825),
.B1(n_748),
.B2(n_767),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_794),
.A2(n_789),
.B(n_804),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_804),
.A2(n_687),
.B(n_756),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_804),
.A2(n_689),
.B1(n_711),
.B2(n_709),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_713),
.A2(n_739),
.B(n_731),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_843),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_752),
.A2(n_582),
.B(n_579),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_710),
.B(n_580),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_713),
.A2(n_739),
.B(n_731),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_689),
.A2(n_710),
.B(n_728),
.C(n_694),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_689),
.A2(n_709),
.B(n_711),
.C(n_546),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_760),
.B(n_771),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_689),
.A2(n_709),
.B(n_711),
.C(n_546),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_752),
.A2(n_582),
.B(n_579),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_752),
.A2(n_582),
.B(n_579),
.Y(n_1014)
);

BUFx8_ASAP7_75t_L g1015 ( 
.A(n_776),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_689),
.B(n_564),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_760),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_752),
.A2(n_582),
.B(n_579),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_689),
.B(n_564),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_689),
.B(n_710),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_689),
.B(n_564),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_752),
.A2(n_582),
.B(n_579),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_688),
.B(n_562),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_689),
.B(n_564),
.Y(n_1024)
);

AO22x1_ASAP7_75t_L g1025 ( 
.A1(n_838),
.A2(n_689),
.B1(n_751),
.B2(n_736),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_704),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_704),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_689),
.B(n_710),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_689),
.B(n_564),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_689),
.B(n_710),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_847),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_760),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_694),
.A2(n_689),
.B(n_731),
.C(n_713),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_1006),
.A2(n_1014),
.B(n_1013),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_977),
.A2(n_978),
.B(n_974),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_906),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_854),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_997),
.A2(n_886),
.B(n_975),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_983),
.A2(n_910),
.B(n_902),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_857),
.B(n_1020),
.Y(n_1040)
);

AO21x1_ASAP7_75t_L g1041 ( 
.A1(n_1020),
.A2(n_1030),
.B(n_941),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_900),
.A2(n_890),
.B(n_979),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_1017),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_959),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1030),
.B(n_1016),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1033),
.A2(n_1009),
.B(n_1008),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1023),
.B(n_877),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_882),
.A2(n_883),
.A3(n_866),
.B(n_896),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_988),
.A2(n_989),
.B(n_995),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_L g1051 ( 
.A(n_959),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_858),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_SL g1053 ( 
.A1(n_871),
.A2(n_861),
.B(n_923),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_970),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_970),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_993),
.A2(n_885),
.B(n_862),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1033),
.A2(n_1004),
.B(n_1010),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_855),
.A2(n_967),
.B(n_965),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_1024),
.A2(n_1029),
.B(n_905),
.C(n_1012),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_991),
.A2(n_904),
.B(n_873),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_986),
.A2(n_875),
.B(n_899),
.Y(n_1061)
);

AO31x2_ASAP7_75t_L g1062 ( 
.A1(n_973),
.A2(n_1003),
.A3(n_972),
.B(n_981),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_914),
.A2(n_865),
.B(n_863),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_976),
.A2(n_990),
.B(n_966),
.C(n_907),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_857),
.B(n_867),
.C(n_878),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_1027),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1028),
.A2(n_1007),
.B1(n_864),
.B2(n_933),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_917),
.B(n_860),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1017),
.A2(n_1032),
.B(n_881),
.Y(n_1069)
);

AOI21xp33_ASAP7_75t_L g1070 ( 
.A1(n_918),
.A2(n_961),
.B(n_954),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1017),
.A2(n_1032),
.B(n_992),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1032),
.A2(n_1017),
.B(n_984),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_976),
.B(n_867),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_942),
.B(n_892),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_880),
.B(n_950),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1032),
.A2(n_996),
.B(n_908),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_958),
.A2(n_1000),
.B(n_1011),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_859),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_1011),
.A2(n_931),
.B(n_968),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_950),
.B(n_946),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_912),
.B(n_916),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_874),
.A2(n_987),
.B(n_856),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_912),
.B(n_916),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_932),
.A2(n_963),
.B(n_935),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_942),
.B(n_994),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_969),
.B(n_953),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_884),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_948),
.A2(n_936),
.B(n_1031),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_928),
.A2(n_927),
.B(n_924),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1026),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_938),
.A2(n_887),
.B(n_915),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_894),
.B(n_1026),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_925),
.A2(n_869),
.B(n_864),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_884),
.Y(n_1094)
);

AND2x6_ASAP7_75t_L g1095 ( 
.A(n_872),
.B(n_876),
.Y(n_1095)
);

AO22x1_ASAP7_75t_L g1096 ( 
.A1(n_926),
.A2(n_998),
.B1(n_955),
.B2(n_999),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1005),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_971),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_956),
.A2(n_934),
.B(n_888),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_879),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_888),
.A2(n_895),
.B(n_897),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_985),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_957),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_921),
.B(n_929),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_937),
.B(n_901),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_943),
.A2(n_889),
.A3(n_939),
.B(n_952),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_926),
.B(n_920),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_911),
.A2(n_962),
.B1(n_945),
.B2(n_964),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_898),
.B(n_891),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_SL g1110 ( 
.A1(n_962),
.A2(n_980),
.B(n_930),
.C(n_922),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_959),
.B(n_893),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_940),
.A2(n_889),
.B(n_898),
.Y(n_1112)
);

OAI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_911),
.A2(n_919),
.B(n_868),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_985),
.B(n_999),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_959),
.B(n_1002),
.Y(n_1115)
);

AOI21x1_ASAP7_75t_L g1116 ( 
.A1(n_951),
.A2(n_898),
.B(n_947),
.Y(n_1116)
);

AO22x1_ASAP7_75t_L g1117 ( 
.A1(n_909),
.A2(n_944),
.B1(n_1015),
.B2(n_898),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_949),
.A2(n_868),
.B(n_947),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_949),
.A2(n_898),
.B(n_960),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_903),
.B(n_982),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_960),
.A2(n_1030),
.B1(n_1020),
.B2(n_1016),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_960),
.A2(n_752),
.B(n_760),
.Y(n_1122)
);

OR2x6_ASAP7_75t_L g1123 ( 
.A(n_1027),
.B(n_789),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_906),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1020),
.A2(n_1030),
.B(n_689),
.C(n_1009),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_906),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1033),
.A2(n_1009),
.B(n_1020),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_882),
.A2(n_883),
.A3(n_1009),
.B(n_726),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1020),
.A2(n_1030),
.B1(n_1016),
.B2(n_1019),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_870),
.A2(n_913),
.B(n_974),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1020),
.A2(n_1030),
.B1(n_1016),
.B2(n_1019),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1011),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_882),
.A2(n_883),
.A3(n_1009),
.B(n_726),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_906),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_906),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_906),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_858),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_997),
.A2(n_886),
.B(n_975),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_SL g1150 ( 
.A1(n_981),
.A2(n_941),
.B(n_1001),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1007),
.B(n_857),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_882),
.A2(n_883),
.A3(n_1009),
.B(n_726),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_1017),
.B(n_760),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_997),
.A2(n_886),
.B(n_975),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1033),
.A2(n_1009),
.B(n_1020),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1007),
.B(n_857),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1033),
.A2(n_1009),
.B(n_1020),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_905),
.B(n_923),
.C(n_871),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_882),
.A2(n_883),
.A3(n_1009),
.B(n_726),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_1017),
.B(n_760),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_905),
.B(n_923),
.C(n_871),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_997),
.A2(n_886),
.B(n_975),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1020),
.A2(n_1030),
.B1(n_923),
.B2(n_689),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1020),
.A2(n_1030),
.B1(n_1016),
.B2(n_1019),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_SL g1171 ( 
.A1(n_933),
.A2(n_711),
.B(n_709),
.Y(n_1171)
);

O2A1O1Ixp5_ASAP7_75t_L g1172 ( 
.A1(n_1025),
.A2(n_694),
.B(n_1009),
.C(n_1020),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_870),
.A2(n_913),
.B(n_974),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1033),
.A2(n_1009),
.B(n_1020),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1007),
.B(n_857),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_906),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1011),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1006),
.A2(n_752),
.B(n_760),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1020),
.B(n_1030),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_857),
.B(n_1020),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_997),
.A2(n_886),
.B(n_975),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1020),
.A2(n_1030),
.B1(n_923),
.B2(n_689),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_1156),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1053),
.A2(n_1127),
.B(n_1134),
.C(n_1170),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1036),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1144),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1040),
.B(n_1182),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_1123),
.B(n_1117),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1142),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1045),
.B(n_1124),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1052),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1134),
.A2(n_1137),
.B(n_1170),
.C(n_1130),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1097),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1147),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1045),
.B(n_1124),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1128),
.B(n_1129),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1177),
.B(n_1107),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1178),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1114),
.B(n_1074),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1125),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1035),
.A2(n_1088),
.B(n_1059),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_L g1205 ( 
.A(n_1163),
.B(n_1166),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1081),
.Y(n_1206)
);

AOI222xp33_ASAP7_75t_L g1207 ( 
.A1(n_1113),
.A2(n_1175),
.B1(n_1153),
.B2(n_1128),
.C1(n_1155),
.C2(n_1168),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_1043),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1081),
.Y(n_1209)
);

OAI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1169),
.A2(n_1184),
.B(n_1073),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1145),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1131),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1111),
.B(n_1123),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1137),
.B(n_1041),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1066),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1051),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1043),
.B(n_1051),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1043),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1105),
.B(n_1104),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1090),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1111),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1047),
.Y(n_1222)
);

INVx5_ASAP7_75t_L g1223 ( 
.A(n_1043),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1129),
.A2(n_1139),
.B1(n_1181),
.B2(n_1135),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1035),
.A2(n_1063),
.B(n_1057),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1123),
.B(n_1115),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1054),
.Y(n_1227)
);

INVx3_ASAP7_75t_SL g1228 ( 
.A(n_1120),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1135),
.B(n_1139),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1083),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1104),
.B(n_1073),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1092),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1140),
.A2(n_1153),
.B(n_1181),
.C(n_1143),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1140),
.B(n_1143),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1098),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1103),
.B(n_1155),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1158),
.B(n_1168),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1158),
.B(n_1175),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1055),
.Y(n_1239)
);

INVx3_ASAP7_75t_SL g1240 ( 
.A(n_1120),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1057),
.A2(n_1046),
.B(n_1159),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1083),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1044),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_1086),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1044),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1096),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1102),
.B(n_1100),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1050),
.B(n_1068),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1068),
.B(n_1080),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1085),
.B(n_1065),
.Y(n_1250)
);

CKINVDCx6p67_ASAP7_75t_R g1251 ( 
.A(n_1095),
.Y(n_1251)
);

AND2x4_ASAP7_75t_SL g1252 ( 
.A(n_1138),
.B(n_1179),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1087),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1087),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1108),
.A2(n_1067),
.B1(n_1095),
.B2(n_1110),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1067),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1108),
.B(n_1075),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1156),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1094),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1075),
.B(n_1064),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1046),
.A2(n_1132),
.B(n_1159),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1179),
.B(n_1095),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1094),
.B(n_1072),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_L g1264 ( 
.A(n_1109),
.B(n_1161),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1132),
.B(n_1176),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1161),
.A2(n_1176),
.B(n_1122),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1070),
.B(n_1121),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1165),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1077),
.B(n_1076),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1062),
.B(n_1121),
.Y(n_1270)
);

CKINVDCx14_ASAP7_75t_R g1271 ( 
.A(n_1109),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1034),
.A2(n_1126),
.B(n_1148),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1172),
.B(n_1062),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1165),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1171),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1146),
.A2(n_1180),
.B(n_1174),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1062),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1079),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1118),
.A2(n_1093),
.B(n_1119),
.C(n_1099),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1071),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1069),
.B(n_1101),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1091),
.B(n_1084),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1112),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_1116),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1151),
.A2(n_1162),
.B(n_1042),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1061),
.B(n_1049),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1150),
.Y(n_1287)
);

O2A1O1Ixp5_ASAP7_75t_SL g1288 ( 
.A1(n_1106),
.A2(n_1173),
.B(n_1136),
.C(n_1039),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1133),
.B(n_1141),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1133),
.B(n_1141),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1089),
.A2(n_1056),
.B(n_1149),
.C(n_1183),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1060),
.A2(n_1038),
.B(n_1167),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1154),
.B(n_1164),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1106),
.B(n_1154),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1154),
.B(n_1164),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1164),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1048),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1060),
.B(n_1157),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1156),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1052),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1169),
.B(n_1184),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1036),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1040),
.B(n_1020),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1127),
.A2(n_1020),
.B(n_1030),
.C(n_689),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1144),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1052),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1040),
.B(n_1182),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1169),
.A2(n_1030),
.B1(n_1020),
.B2(n_1016),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_1043),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1040),
.A2(n_1030),
.B1(n_1020),
.B2(n_1182),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1053),
.A2(n_1009),
.B(n_1030),
.C(n_1020),
.Y(n_1313)
);

AND2x2_ASAP7_75t_SL g1314 ( 
.A(n_1169),
.B(n_948),
.Y(n_1314)
);

OAI321xp33_ASAP7_75t_L g1315 ( 
.A1(n_1163),
.A2(n_1166),
.A3(n_962),
.B1(n_1113),
.B2(n_1030),
.C(n_1020),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1051),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1058),
.A2(n_1082),
.B(n_1037),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1090),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1036),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1040),
.B(n_1020),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1127),
.A2(n_1020),
.B(n_1030),
.C(n_689),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1078),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1043),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1040),
.B(n_1020),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1040),
.A2(n_1030),
.B1(n_1020),
.B2(n_1182),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1169),
.A2(n_1030),
.B1(n_1020),
.B2(n_1016),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1111),
.B(n_959),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1111),
.B(n_959),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1090),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1144),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1040),
.B(n_1182),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1308),
.B(n_1333),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1235),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1312),
.A2(n_1327),
.B1(n_1308),
.B2(n_1333),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1193),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1195),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1196),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1189),
.A2(n_1321),
.B1(n_1326),
.B2(n_1303),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1220),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1300),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1246),
.A2(n_1256),
.B1(n_1255),
.B2(n_1315),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1307),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1312),
.A2(n_1327),
.B1(n_1205),
.B2(n_1301),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1212),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1231),
.B(n_1199),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1208),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1323),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1208),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1257),
.B(n_1207),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1208),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1199),
.B(n_1229),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1188),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1281),
.B(n_1269),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1277),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1306),
.Y(n_1357)
);

BUFx2_ASAP7_75t_R g1358 ( 
.A(n_1332),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1301),
.A2(n_1314),
.B1(n_1210),
.B2(n_1328),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1203),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1219),
.B(n_1236),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1187),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1206),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1314),
.A2(n_1271),
.B1(n_1229),
.B2(n_1237),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1220),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1319),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1320),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1289),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1319),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1331),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1237),
.B(n_1200),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1290),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1297),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1234),
.A2(n_1238),
.B1(n_1197),
.B2(n_1192),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1244),
.B(n_1198),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1331),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1209),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1250),
.A2(n_1309),
.B1(n_1296),
.B2(n_1244),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1223),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1309),
.A2(n_1325),
.B1(n_1310),
.B2(n_1304),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1230),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1318),
.B(n_1248),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1242),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1233),
.B(n_1249),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1260),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1227),
.Y(n_1386)
);

BUFx2_ASAP7_75t_R g1387 ( 
.A(n_1228),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1201),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1239),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1233),
.B(n_1224),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1292),
.A2(n_1285),
.B(n_1276),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1287),
.A2(n_1214),
.B1(n_1264),
.B2(n_1280),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1305),
.A2(n_1322),
.B1(n_1232),
.B2(n_1222),
.Y(n_1393)
);

INVx5_ASAP7_75t_L g1394 ( 
.A(n_1223),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1247),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1253),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1204),
.A2(n_1225),
.B(n_1214),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1267),
.A2(n_1265),
.B1(n_1226),
.B2(n_1261),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1254),
.Y(n_1399)
);

AO21x1_ASAP7_75t_L g1400 ( 
.A1(n_1313),
.A2(n_1186),
.B(n_1194),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1232),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1305),
.A2(n_1322),
.B1(n_1224),
.B2(n_1191),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1288),
.A2(n_1272),
.B(n_1317),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1223),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1259),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1202),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1261),
.A2(n_1275),
.B1(n_1241),
.B2(n_1226),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1302),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1284),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1194),
.A2(n_1241),
.B(n_1266),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1225),
.A2(n_1291),
.B(n_1279),
.Y(n_1411)
);

BUFx5_ASAP7_75t_L g1412 ( 
.A(n_1278),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1311),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1211),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1215),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1190),
.A2(n_1228),
.B1(n_1240),
.B2(n_1216),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1190),
.A2(n_1213),
.B1(n_1316),
.B2(n_1216),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1284),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1185),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1221),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1283),
.A2(n_1263),
.B(n_1298),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1273),
.A2(n_1294),
.B(n_1270),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1282),
.A2(n_1286),
.B(n_1293),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1240),
.Y(n_1425)
);

AO21x1_ASAP7_75t_SL g1426 ( 
.A1(n_1251),
.A2(n_1295),
.B(n_1284),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1217),
.A2(n_1185),
.B(n_1299),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1284),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1263),
.A2(n_1213),
.B1(n_1295),
.B2(n_1316),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1286),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1282),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1243),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1299),
.B(n_1274),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1258),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1262),
.B(n_1330),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1258),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1217),
.A2(n_1311),
.B(n_1268),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1268),
.A2(n_1245),
.B(n_1258),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1329),
.A2(n_1330),
.B1(n_1262),
.B2(n_1252),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1329),
.A2(n_1245),
.B1(n_1258),
.B2(n_1324),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1218),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1218),
.Y(n_1442)
);

AO21x1_ASAP7_75t_L g1443 ( 
.A1(n_1311),
.A2(n_1218),
.B(n_1324),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1311),
.A2(n_1166),
.B1(n_1163),
.B2(n_1308),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1324),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1324),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1193),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1193),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1193),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1231),
.B(n_1257),
.Y(n_1450)
);

CKINVDCx11_ASAP7_75t_R g1451 ( 
.A(n_1228),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1193),
.Y(n_1452)
);

INVx6_ASAP7_75t_L g1453 ( 
.A(n_1208),
.Y(n_1453)
);

BUFx8_ASAP7_75t_L g1454 ( 
.A(n_1201),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1193),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1301),
.A2(n_1166),
.B1(n_1163),
.B2(n_923),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1193),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1285),
.A2(n_1204),
.B(n_1272),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1308),
.A2(n_1053),
.B1(n_923),
.B2(n_1163),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1356),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1410),
.A2(n_1403),
.B(n_1397),
.Y(n_1461)
);

AOI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1390),
.A2(n_1402),
.B(n_1384),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1450),
.B(n_1361),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1370),
.Y(n_1464)
);

AOI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1393),
.A2(n_1400),
.B(n_1391),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1370),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1359),
.A2(n_1336),
.B1(n_1351),
.B2(n_1456),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1424),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1394),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1450),
.B(n_1361),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1334),
.B(n_1340),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1414),
.Y(n_1472)
);

INVxp33_ASAP7_75t_L g1473 ( 
.A(n_1408),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1368),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1423),
.B(n_1371),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1423),
.B(n_1372),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1424),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1459),
.A2(n_1345),
.B(n_1444),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1353),
.B(n_1347),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1430),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1412),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1458),
.A2(n_1411),
.B(n_1400),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1412),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1412),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1371),
.B(n_1351),
.Y(n_1485)
);

INVxp67_ASAP7_75t_SL g1486 ( 
.A(n_1341),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1385),
.B(n_1431),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1346),
.B(n_1382),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1354),
.Y(n_1489)
);

AO21x1_ASAP7_75t_SL g1490 ( 
.A1(n_1392),
.A2(n_1373),
.B(n_1417),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_SL g1491 ( 
.A(n_1387),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_SL g1492 ( 
.A(n_1354),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1373),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1420),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1417),
.Y(n_1495)
);

INVx5_ASAP7_75t_L g1496 ( 
.A(n_1394),
.Y(n_1496)
);

AO21x1_ASAP7_75t_SL g1497 ( 
.A1(n_1378),
.A2(n_1407),
.B(n_1422),
.Y(n_1497)
);

OA21x2_ASAP7_75t_L g1498 ( 
.A1(n_1409),
.A2(n_1419),
.B(n_1428),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1409),
.A2(n_1419),
.B(n_1428),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1457),
.B(n_1385),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1382),
.B(n_1398),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1337),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1375),
.B(n_1363),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1357),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1415),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1375),
.B(n_1377),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1355),
.B(n_1416),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1365),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1338),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1357),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1339),
.Y(n_1511)
);

CKINVDCx16_ASAP7_75t_R g1512 ( 
.A(n_1388),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1342),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1406),
.B(n_1366),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1369),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1344),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1376),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1411),
.B(n_1401),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1374),
.A2(n_1427),
.B(n_1447),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1448),
.Y(n_1520)
);

AOI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1443),
.A2(n_1427),
.B(n_1405),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1449),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1452),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1455),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1443),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1381),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1383),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1436),
.B(n_1434),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1433),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1395),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1379),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1388),
.Y(n_1532)
);

CKINVDCx8_ASAP7_75t_R g1533 ( 
.A(n_1394),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1396),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1399),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1426),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1437),
.A2(n_1404),
.B(n_1429),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1389),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1488),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1479),
.B(n_1343),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1460),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1494),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1467),
.A2(n_1364),
.B1(n_1471),
.B2(n_1478),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1536),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1518),
.B(n_1380),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1494),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1525),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1475),
.B(n_1426),
.Y(n_1548)
);

INVx4_ASAP7_75t_R g1549 ( 
.A(n_1491),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1518),
.B(n_1425),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1536),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1463),
.B(n_1349),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1470),
.B(n_1386),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1498),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1499),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1464),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1515),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1501),
.B(n_1442),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1508),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1529),
.B(n_1486),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1466),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1493),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1485),
.B(n_1495),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1493),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1485),
.B(n_1445),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1503),
.B(n_1446),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1481),
.B(n_1446),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1503),
.B(n_1435),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1476),
.B(n_1335),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1481),
.B(n_1394),
.Y(n_1572)
);

INVx5_ASAP7_75t_L g1573 ( 
.A(n_1536),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1506),
.B(n_1335),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1517),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1483),
.B(n_1394),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1497),
.A2(n_1418),
.B1(n_1451),
.B2(n_1454),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1480),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1497),
.A2(n_1451),
.B1(n_1454),
.B2(n_1421),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1476),
.B(n_1362),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1508),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1472),
.A2(n_1360),
.B1(n_1362),
.B2(n_1367),
.C(n_1435),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1506),
.B(n_1367),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1517),
.B(n_1454),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1482),
.B(n_1360),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1512),
.B(n_1358),
.Y(n_1586)
);

NAND2x1_ASAP7_75t_L g1587 ( 
.A(n_1507),
.B(n_1453),
.Y(n_1587)
);

AOI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1473),
.A2(n_1440),
.B1(n_1439),
.B2(n_1438),
.C(n_1432),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1558),
.B(n_1500),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1578),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1562),
.B(n_1500),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1543),
.A2(n_1512),
.B1(n_1507),
.B2(n_1532),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1563),
.B(n_1500),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1579),
.A2(n_1462),
.B(n_1465),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1577),
.A2(n_1588),
.B1(n_1540),
.B2(n_1582),
.C(n_1539),
.Y(n_1595)
);

NAND4xp25_ASAP7_75t_L g1596 ( 
.A(n_1551),
.B(n_1514),
.C(n_1505),
.D(n_1511),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1542),
.B(n_1482),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1557),
.A2(n_1530),
.B1(n_1509),
.B2(n_1511),
.C(n_1513),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1565),
.B(n_1551),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1584),
.B(n_1462),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1502),
.Y(n_1601)
);

NAND3xp33_ASAP7_75t_L g1602 ( 
.A(n_1585),
.B(n_1514),
.C(n_1523),
.Y(n_1602)
);

OAI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1545),
.A2(n_1465),
.B(n_1524),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1559),
.B(n_1522),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1571),
.B(n_1522),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1571),
.B(n_1509),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1586),
.B(n_1504),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1585),
.B(n_1545),
.C(n_1520),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1547),
.A2(n_1507),
.B1(n_1496),
.B2(n_1492),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1567),
.A2(n_1507),
.B1(n_1490),
.B2(n_1519),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1548),
.A2(n_1521),
.B(n_1526),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1548),
.A2(n_1521),
.B(n_1526),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1567),
.A2(n_1507),
.B1(n_1490),
.B2(n_1519),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1516),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1547),
.A2(n_1527),
.B(n_1531),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1550),
.A2(n_1527),
.B(n_1531),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1561),
.B(n_1510),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1561),
.B(n_1520),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1581),
.B(n_1523),
.Y(n_1620)
);

OAI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1587),
.A2(n_1524),
.B1(n_1534),
.B2(n_1535),
.C(n_1468),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1574),
.B(n_1489),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1581),
.B(n_1534),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1583),
.B(n_1432),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1550),
.A2(n_1519),
.B1(n_1537),
.B2(n_1528),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1560),
.B(n_1535),
.C(n_1538),
.Y(n_1626)
);

OAI221xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1560),
.A2(n_1487),
.B1(n_1553),
.B2(n_1554),
.C(n_1546),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1568),
.B(n_1477),
.Y(n_1628)
);

OA211x2_ASAP7_75t_L g1629 ( 
.A1(n_1587),
.A2(n_1533),
.B(n_1496),
.C(n_1469),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1569),
.B(n_1477),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1569),
.B(n_1477),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1552),
.A2(n_1531),
.B(n_1474),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1569),
.B(n_1484),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1573),
.B(n_1496),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1544),
.A2(n_1469),
.B(n_1350),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1564),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1590),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1630),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1590),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1626),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1597),
.B(n_1602),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1617),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1617),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1628),
.B(n_1631),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1633),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1633),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1606),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1626),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1605),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1566),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1619),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1592),
.A2(n_1482),
.B1(n_1461),
.B2(n_1570),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1620),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1608),
.B(n_1601),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1623),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1600),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1608),
.B(n_1555),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1603),
.B(n_1541),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1593),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1603),
.B(n_1541),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1556),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1645),
.B(n_1599),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1653),
.A2(n_1595),
.B(n_1594),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1637),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1655),
.B(n_1604),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1655),
.B(n_1641),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1655),
.B(n_1627),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1641),
.B(n_1636),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1642),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1598),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1642),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1642),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1645),
.B(n_1609),
.Y(n_1675)
);

OAI21xp33_ASAP7_75t_L g1676 ( 
.A1(n_1640),
.A2(n_1596),
.B(n_1611),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1637),
.B(n_1634),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1657),
.B(n_1607),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1636),
.B(n_1591),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1589),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1645),
.B(n_1613),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1637),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1640),
.B(n_1612),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1649),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1639),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1647),
.B(n_1615),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1646),
.B(n_1632),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1643),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1649),
.B(n_1616),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1646),
.B(n_1572),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1639),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1647),
.B(n_1570),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1646),
.B(n_1572),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1618),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1646),
.B(n_1572),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1660),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1638),
.B(n_1572),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1576),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1624),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1690),
.B(n_1638),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1678),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1697),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1670),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1678),
.B(n_1639),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1670),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1672),
.Y(n_1709)
);

XNOR2xp5_ASAP7_75t_L g1710 ( 
.A(n_1668),
.B(n_1549),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1673),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1699),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1690),
.B(n_1638),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1673),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1669),
.B(n_1651),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1669),
.B(n_1651),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1674),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1678),
.B(n_1639),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1665),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1672),
.B(n_1648),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1674),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1648),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1687),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1677),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1677),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1684),
.Y(n_1726)
);

NAND2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1687),
.B(n_1653),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1680),
.B(n_1622),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1675),
.B(n_1638),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1667),
.B(n_1658),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1667),
.B(n_1658),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1684),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1691),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1691),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1675),
.B(n_1638),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1665),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1671),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1679),
.B(n_1644),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1671),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1679),
.B(n_1644),
.Y(n_1740)
);

AO21x1_ASAP7_75t_L g1741 ( 
.A1(n_1664),
.A2(n_1658),
.B(n_1659),
.Y(n_1741)
);

AOI21xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1664),
.A2(n_1549),
.B(n_1659),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1683),
.B(n_1700),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1671),
.Y(n_1744)
);

OAI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1676),
.A2(n_1661),
.B(n_1662),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1710),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1710),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1706),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1723),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1706),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1743),
.B(n_1683),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1704),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1715),
.B(n_1668),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1721),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1709),
.B(n_1702),
.Y(n_1756)
);

NAND3x1_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_1692),
.C(n_1689),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1692),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1704),
.B(n_1686),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1729),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1743),
.B(n_1686),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1720),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1721),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1745),
.A2(n_1681),
.B1(n_1666),
.B2(n_1695),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1707),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1724),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1715),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1741),
.B(n_1666),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1727),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1728),
.B(n_1742),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1707),
.Y(n_1771)
);

INVx3_ASAP7_75t_SL g1772 ( 
.A(n_1730),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1716),
.B(n_1681),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1707),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1716),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1722),
.B(n_1663),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1727),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1738),
.B(n_1700),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1729),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1724),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1730),
.B(n_1682),
.Y(n_1781)
);

OAI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1769),
.A2(n_1735),
.B(n_1731),
.Y(n_1782)
);

AND2x2_ASAP7_75t_SL g1783 ( 
.A(n_1770),
.B(n_1735),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1756),
.B(n_1769),
.Y(n_1784)
);

NAND5xp2_ASAP7_75t_SL g1785 ( 
.A(n_1761),
.B(n_1703),
.C(n_1713),
.D(n_1738),
.E(n_1740),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1748),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1750),
.B(n_1746),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1747),
.B(n_1731),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1752),
.B(n_1740),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1752),
.B(n_1703),
.Y(n_1790)
);

AOI21xp33_ASAP7_75t_L g1791 ( 
.A1(n_1757),
.A2(n_1719),
.B(n_1732),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1772),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1777),
.A2(n_1736),
.B1(n_1718),
.B2(n_1719),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1777),
.A2(n_1713),
.B(n_1661),
.C(n_1739),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1754),
.B(n_1708),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1772),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1748),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1749),
.B(n_1678),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1772),
.B(n_1768),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1751),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1767),
.B(n_1718),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1757),
.A2(n_1629),
.B1(n_1662),
.B2(n_1701),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1762),
.B(n_1693),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1751),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1758),
.A2(n_1718),
.B(n_1714),
.Y(n_1805)
);

AO22x1_ASAP7_75t_L g1806 ( 
.A1(n_1759),
.A2(n_1725),
.B1(n_1726),
.B2(n_1711),
.Y(n_1806)
);

INVxp67_ASAP7_75t_SL g1807 ( 
.A(n_1753),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1792),
.B(n_1761),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1796),
.Y(n_1809)
);

NAND2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1796),
.B(n_1759),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1796),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1792),
.B(n_1775),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1807),
.B(n_1759),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1786),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1787),
.B(n_1754),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1797),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1799),
.A2(n_1779),
.B1(n_1760),
.B2(n_1759),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1795),
.B(n_1773),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1788),
.B(n_1760),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1789),
.B(n_1779),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1783),
.Y(n_1821)
);

OAI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1799),
.A2(n_1773),
.B1(n_1764),
.B2(n_1776),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1790),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1784),
.B(n_1781),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1782),
.B(n_1765),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1801),
.B(n_1765),
.Y(n_1827)
);

OAI31xp33_ASAP7_75t_L g1828 ( 
.A1(n_1822),
.A2(n_1793),
.A3(n_1794),
.B(n_1791),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_L g1829 ( 
.A(n_1822),
.B(n_1817),
.C(n_1813),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1825),
.A2(n_1785),
.B1(n_1791),
.B2(n_1806),
.C(n_1805),
.Y(n_1830)
);

NOR3xp33_ASAP7_75t_L g1831 ( 
.A(n_1812),
.B(n_1798),
.C(n_1804),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1808),
.B(n_1778),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1808),
.B(n_1771),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1821),
.A2(n_1802),
.B1(n_1803),
.B2(n_1771),
.C(n_1774),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1819),
.A2(n_1778),
.B(n_1774),
.Y(n_1835)
);

AOI21xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1810),
.A2(n_1763),
.B(n_1755),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1815),
.A2(n_1763),
.B(n_1755),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1810),
.A2(n_1780),
.B(n_1766),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1809),
.B(n_1766),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1818),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1829),
.B(n_1811),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1830),
.A2(n_1820),
.B1(n_1823),
.B2(n_1826),
.Y(n_1842)
);

AOI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1828),
.A2(n_1826),
.B(n_1827),
.C(n_1818),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1840),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1832),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1836),
.B(n_1820),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1831),
.B(n_1838),
.C(n_1834),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1833),
.B(n_1827),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1835),
.B(n_1814),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1839),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1837),
.Y(n_1851)
);

OAI211xp5_ASAP7_75t_L g1852 ( 
.A1(n_1828),
.A2(n_1824),
.B(n_1816),
.C(n_1780),
.Y(n_1852)
);

AOI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1828),
.A2(n_1732),
.B(n_1733),
.C(n_1737),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1847),
.A2(n_1733),
.B1(n_1744),
.B2(n_1737),
.C(n_1717),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1848),
.B(n_1734),
.Y(n_1855)
);

NAND2x1p5_ASAP7_75t_L g1856 ( 
.A(n_1841),
.B(n_1379),
.Y(n_1856)
);

NOR3xp33_ASAP7_75t_L g1857 ( 
.A(n_1852),
.B(n_1744),
.C(n_1621),
.Y(n_1857)
);

NAND4xp25_ASAP7_75t_L g1858 ( 
.A(n_1843),
.B(n_1629),
.C(n_1635),
.D(n_1701),
.Y(n_1858)
);

NAND3x1_ASAP7_75t_L g1859 ( 
.A(n_1842),
.B(n_1694),
.C(n_1693),
.Y(n_1859)
);

INVxp67_ASAP7_75t_SL g1860 ( 
.A(n_1856),
.Y(n_1860)
);

NOR2x1_ASAP7_75t_L g1861 ( 
.A(n_1855),
.B(n_1851),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1857),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1859),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1854),
.B(n_1848),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1858),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1858),
.A2(n_1845),
.B1(n_1853),
.B2(n_1846),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_SL g1867 ( 
.A(n_1866),
.B(n_1844),
.C(n_1850),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1862),
.B(n_1849),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1861),
.A2(n_1688),
.B(n_1685),
.C(n_1694),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1864),
.B(n_1685),
.Y(n_1870)
);

OAI211xp5_ASAP7_75t_L g1871 ( 
.A1(n_1860),
.A2(n_1533),
.B(n_1635),
.C(n_1441),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1863),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1868),
.B(n_1865),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1872),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1870),
.B(n_1696),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1874),
.B(n_1867),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1876),
.A2(n_1873),
.B1(n_1871),
.B2(n_1875),
.C(n_1869),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1688),
.B(n_1685),
.Y(n_1878)
);

OA21x2_ASAP7_75t_L g1879 ( 
.A1(n_1877),
.A2(n_1688),
.B(n_1696),
.Y(n_1879)
);

OA21x2_ASAP7_75t_L g1880 ( 
.A1(n_1878),
.A2(n_1698),
.B(n_1663),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1879),
.A2(n_1656),
.B1(n_1654),
.B2(n_1652),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1880),
.B(n_1878),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1881),
.B(n_1698),
.Y(n_1883)
);

XOR2x1_ASAP7_75t_L g1884 ( 
.A(n_1882),
.B(n_1348),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1884),
.A2(n_1883),
.B1(n_1441),
.B2(n_1652),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1885),
.A2(n_1652),
.B1(n_1654),
.B2(n_1656),
.C(n_1648),
.Y(n_1886)
);

AOI211xp5_ASAP7_75t_L g1887 ( 
.A1(n_1886),
.A2(n_1413),
.B(n_1350),
.C(n_1352),
.Y(n_1887)
);


endmodule