module fake_jpeg_3774_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_32),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_37),
.Y(n_62)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_44),
.B(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_24),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_2),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_30),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_47),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_55),
.B(n_32),
.C(n_8),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_3),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_54),
.B(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_14),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_5),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_51),
.B1(n_55),
.B2(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_65),
.B1(n_72),
.B2(n_48),
.Y(n_107)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_6),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_91),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_108),
.B1(n_111),
.B2(n_84),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_48),
.B1(n_45),
.B2(n_68),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_111),
.B(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_86),
.B1(n_103),
.B2(n_100),
.Y(n_124)
);

AOI22x1_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_64),
.B1(n_53),
.B2(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_88),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_64),
.B1(n_57),
.B2(n_59),
.Y(n_111)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_102),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_77),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_119),
.C(n_121),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_94),
.B1(n_75),
.B2(n_85),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_123),
.B(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_124),
.C(n_125),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_84),
.C(n_74),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_84),
.B(n_74),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_90),
.C(n_95),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_109),
.C(n_105),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_130),
.B(n_137),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_109),
.A3(n_90),
.B1(n_10),
.B2(n_99),
.C1(n_82),
.C2(n_76),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_99),
.B(n_91),
.C(n_106),
.D(n_97),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_118),
.B(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_143),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_113),
.C(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_145),
.Y(n_148)
);

NOR2x1_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_116),
.C(n_97),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_138),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_151),
.C(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

OAI221xp5_ASAP7_75t_L g154 ( 
.A1(n_148),
.A2(n_146),
.B1(n_141),
.B2(n_133),
.C(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_149),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_153),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_157),
.B(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_160),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule