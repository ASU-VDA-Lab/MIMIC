module fake_jpeg_5860_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_33),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_16),
.C(n_28),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_18),
.C(n_21),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_48),
.B1(n_55),
.B2(n_72),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_20),
.B(n_26),
.C(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_32),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_23),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_62),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_24),
.B1(n_32),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_59),
.B1(n_25),
.B2(n_16),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_24),
.B1(n_29),
.B2(n_25),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_25),
.B(n_29),
.C(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_38),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_81)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_38),
.A2(n_12),
.B(n_10),
.Y(n_72)
);

OA22x2_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_51),
.B1(n_71),
.B2(n_69),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_84),
.B1(n_64),
.B2(n_50),
.Y(n_115)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_80),
.B(n_93),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_60),
.B1(n_70),
.B2(n_49),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_43),
.B1(n_40),
.B2(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_19),
.B1(n_27),
.B2(n_21),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_50),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_95),
.B1(n_49),
.B2(n_65),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_21),
.B1(n_18),
.B2(n_11),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_52),
.C(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_101),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_47),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_45),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_108),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_76),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_34),
.C(n_39),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_112),
.B(n_30),
.Y(n_138)
);

AOI22x1_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_39),
.B1(n_43),
.B2(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_73),
.Y(n_136)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_75),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_134),
.B(n_138),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_82),
.B1(n_97),
.B2(n_63),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_114),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_75),
.B1(n_63),
.B2(n_57),
.Y(n_132)
);

OR2x2_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_0),
.Y(n_134)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_56),
.B1(n_49),
.B2(n_54),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_56),
.B1(n_70),
.B2(n_85),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_65),
.B1(n_92),
.B2(n_116),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_30),
.B(n_85),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_150),
.B(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_104),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_158),
.B1(n_166),
.B2(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_156),
.B(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_100),
.B1(n_111),
.B2(n_108),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_105),
.B1(n_111),
.B2(n_101),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_169),
.B(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_174),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_101),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_120),
.B1(n_109),
.B2(n_102),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_70),
.B1(n_78),
.B2(n_94),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_39),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_131),
.C(n_133),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_79),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_144),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_128),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_189),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_160),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_138),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_131),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_192),
.B(n_156),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_148),
.C(n_125),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_197),
.C(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_151),
.B1(n_141),
.B2(n_132),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_199),
.B(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_154),
.A2(n_146),
.B1(n_150),
.B2(n_141),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_140),
.C(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_134),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_159),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_217),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_157),
.B1(n_155),
.B2(n_161),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_211),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_153),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_214),
.C(n_223),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_216),
.A2(n_86),
.B1(n_78),
.B2(n_66),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_162),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_161),
.B(n_134),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_177),
.C(n_170),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_172),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_194),
.C(n_179),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_79),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_227),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_149),
.B(n_107),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_168),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_231),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_79),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_201),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_116),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_179),
.B1(n_190),
.B2(n_195),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_229),
.B1(n_221),
.B2(n_226),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_252),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_213),
.C(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_207),
.C(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_249),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_1),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_169),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_152),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_253),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_152),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_246),
.C(n_243),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_216),
.B1(n_224),
.B2(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_229),
.B(n_221),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_239),
.C(n_233),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_149),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_235),
.A2(n_206),
.B1(n_149),
.B2(n_66),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_270),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_2),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_267),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_147),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_65),
.B1(n_74),
.B2(n_147),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_242),
.B(n_12),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_147),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_232),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_233),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_286),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_255),
.B(n_249),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_288),
.C(n_268),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_243),
.C(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_264),
.C(n_262),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_239),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_241),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_277),
.B1(n_280),
.B2(n_256),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_302),
.A3(n_282),
.B1(n_288),
.B2(n_285),
.C1(n_74),
.C2(n_11),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_265),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_294),
.B(n_297),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_279),
.A2(n_287),
.B1(n_269),
.B2(n_258),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_298),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_263),
.C(n_255),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_89),
.C(n_66),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_301),
.C(n_22),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_43),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_306),
.C(n_311),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_15),
.C(n_14),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_2),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_74),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_308),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_22),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_10),
.C2(n_7),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_14),
.C(n_3),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_313),
.B(n_309),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_22),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_7),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_22),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_8),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_6),
.C(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_318),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_22),
.B(n_6),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_319),
.B(n_9),
.Y(n_324)
);

NAND4xp25_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_3),
.C(n_6),
.D(n_8),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_6),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_9),
.B1(n_315),
.B2(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_9),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_326),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_328),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_323),
.B(n_329),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_327),
.Y(n_332)
);


endmodule