module fake_jpeg_21388_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_127;
wire n_76;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_13),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_72),
.Y(n_95)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_52),
.B1(n_80),
.B2(n_86),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_63),
.B1(n_62),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_52),
.B1(n_82),
.B2(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_1),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_70),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_65),
.B1(n_75),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_56),
.B1(n_57),
.B2(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_108),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_87),
.B1(n_85),
.B2(n_78),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_96),
.B1(n_79),
.B2(n_78),
.Y(n_113)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_64),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_1),
.Y(n_125)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_126),
.B1(n_8),
.B2(n_9),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_50),
.B(n_61),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_121),
.B(n_127),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_123),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_61),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_111),
.C(n_121),
.Y(n_133)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_66),
.B1(n_68),
.B2(n_74),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_66),
.B1(n_77),
.B2(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_77),
.B1(n_69),
.B2(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_76),
.B(n_54),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_54),
.B(n_5),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_102),
.B1(n_60),
.B2(n_58),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_122),
.B1(n_118),
.B2(n_11),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_3),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_30),
.C(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_28),
.C(n_41),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_141),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_33),
.B(n_40),
.C(n_39),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_140),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_146),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_155),
.B1(n_152),
.B2(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_133),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_147),
.B(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_147),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_36),
.B(n_22),
.C(n_25),
.D(n_27),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_138),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_49),
.B1(n_32),
.B2(n_34),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_136),
.C(n_129),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_38),
.B(n_151),
.C(n_14),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g168 ( 
.A(n_167),
.Y(n_168)
);


endmodule