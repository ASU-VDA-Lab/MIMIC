module fake_jpeg_5850_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_8),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_22),
.Y(n_47)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_16),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_21),
.B(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_60),
.B1(n_25),
.B2(n_26),
.Y(n_78)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_23),
.B1(n_19),
.B2(n_39),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_42),
.B1(n_38),
.B2(n_16),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_21),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_73),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_52),
.B1(n_56),
.B2(n_48),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_37),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_79),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_61),
.B1(n_57),
.B2(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_52),
.B1(n_61),
.B2(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_67),
.B1(n_40),
.B2(n_15),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_92),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_89),
.B(n_94),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_53),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_45),
.B1(n_38),
.B2(n_54),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_49),
.B1(n_51),
.B2(n_76),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_46),
.C(n_44),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_96),
.C(n_69),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_44),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_70),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_40),
.B1(n_75),
.B2(n_41),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_70),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_47),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_114),
.C(n_36),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_110),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_47),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_41),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_119),
.B1(n_120),
.B2(n_92),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_74),
.C(n_46),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_117),
.Y(n_130)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_80),
.B1(n_78),
.B2(n_62),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_121),
.B(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_59),
.B(n_22),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_59),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_22),
.B(n_37),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_26),
.B(n_25),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_86),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_138),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_119),
.B(n_108),
.C(n_112),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_90),
.B1(n_101),
.B2(n_85),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

XNOR2x2_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_128),
.C(n_132),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_90),
.A3(n_102),
.B1(n_86),
.B2(n_83),
.C1(n_84),
.C2(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_81),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_98),
.B1(n_99),
.B2(n_34),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_141),
.B(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_107),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_82),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_41),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_21),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_75),
.B1(n_41),
.B2(n_25),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_63),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_118),
.B1(n_127),
.B2(n_140),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_161),
.B1(n_105),
.B2(n_26),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_153),
.B(n_142),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_103),
.B(n_115),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_163),
.B1(n_135),
.B2(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_119),
.B1(n_108),
.B2(n_117),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_160),
.B1(n_158),
.B2(n_149),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_135),
.B1(n_141),
.B2(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_110),
.B1(n_123),
.B2(n_104),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_34),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_104),
.C(n_105),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_139),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_167),
.B(n_168),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_138),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_130),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_162),
.C(n_148),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_160),
.B(n_159),
.C(n_154),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_179),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_34),
.B1(n_29),
.B2(n_18),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_159),
.B1(n_161),
.B2(n_72),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_184),
.B(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_190),
.C(n_192),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_189),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_153),
.C(n_155),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_72),
.C(n_29),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_177),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_197),
.C(n_4),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_173),
.B1(n_170),
.B2(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_198),
.B1(n_202),
.B2(n_1),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_199),
.B(n_203),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_166),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_172),
.B1(n_29),
.B2(n_0),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_9),
.B(n_1),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_0),
.B1(n_18),
.B2(n_3),
.Y(n_202)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_182),
.B(n_191),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_209),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_208),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_207),
.C(n_211),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_4),
.C(n_5),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_5),
.Y(n_208)
);

OAI221xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.C(n_11),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_10),
.C(n_11),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_200),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_220),
.C(n_221),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_12),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_12),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_213),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_212),
.Y(n_226)
);

AOI321xp33_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_218),
.C(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_13),
.Y(n_228)
);


endmodule