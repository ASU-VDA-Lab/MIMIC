module fake_jpeg_389_n_677 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_677);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_677;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_70),
.Y(n_211)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_74),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_76),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_77),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_7),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_91),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_18),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_83),
.Y(n_209)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_87),
.B(n_130),
.Y(n_166)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_90),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_35),
.B(n_7),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_17),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_101),
.B(n_112),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_17),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_45),
.Y(n_119)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_54),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_128),
.Y(n_157)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_21),
.Y(n_127)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_23),
.B(n_6),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_24),
.Y(n_129)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_24),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_25),
.Y(n_197)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_21),
.Y(n_132)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_76),
.A2(n_50),
.B1(n_46),
.B2(n_44),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_133),
.A2(n_167),
.B1(n_210),
.B2(n_227),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_50),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_138),
.B(n_173),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_83),
.A2(n_33),
.B1(n_58),
.B2(n_57),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_139),
.A2(n_178),
.B1(n_188),
.B2(n_204),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_152),
.B(n_225),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_44),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_155),
.B(n_0),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_119),
.A2(n_50),
.B1(n_46),
.B2(n_44),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_77),
.B(n_55),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_37),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_174),
.B(n_16),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_61),
.A2(n_29),
.B1(n_46),
.B2(n_21),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_62),
.A2(n_29),
.B1(n_59),
.B2(n_33),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_197),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_58),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_67),
.Y(n_199)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_70),
.B(n_57),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_65),
.A2(n_55),
.B1(n_53),
.B2(n_48),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_96),
.A2(n_29),
.B1(n_48),
.B2(n_43),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_213),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_60),
.B(n_34),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_75),
.Y(n_247)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_118),
.Y(n_221)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_92),
.Y(n_222)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_73),
.Y(n_223)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_79),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_82),
.Y(n_226)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_81),
.A2(n_75),
.B1(n_60),
.B2(n_105),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_229),
.B(n_237),
.Y(n_312)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_230),
.Y(n_353)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_231),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_38),
.B1(n_37),
.B2(n_43),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_234),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_236),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_172),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_238),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_211),
.A2(n_38),
.B1(n_53),
.B2(n_34),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_239),
.A2(n_267),
.B1(n_294),
.B2(n_295),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_188),
.A2(n_90),
.B1(n_116),
.B2(n_113),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_244),
.A2(n_177),
.B1(n_165),
.B2(n_193),
.Y(n_324)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_144),
.Y(n_246)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_246),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_265),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_137),
.B(n_0),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_248),
.B(n_261),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_172),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_249),
.B(n_260),
.Y(n_319)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_251),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_252),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_138),
.B(n_107),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_253),
.Y(n_361)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_157),
.B(n_151),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_259),
.B(n_263),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_151),
.A2(n_103),
.B(n_99),
.C(n_86),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_0),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_215),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_157),
.B(n_95),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_201),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_282),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_220),
.A2(n_106),
.B1(n_9),
.B2(n_11),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_181),
.Y(n_268)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_268),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_134),
.A2(n_5),
.B1(n_14),
.B2(n_12),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_269),
.A2(n_271),
.B1(n_274),
.B2(n_292),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_143),
.B(n_0),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_272),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_210),
.A2(n_9),
.B1(n_14),
.B2(n_3),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_149),
.B(n_1),
.Y(n_272)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_168),
.Y(n_273)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_273),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_205),
.A2(n_9),
.B1(n_14),
.B2(n_3),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_275),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_142),
.B(n_5),
.C(n_14),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_303),
.C(n_163),
.Y(n_322)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_150),
.Y(n_277)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_212),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_279),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_216),
.B(n_1),
.Y(n_279)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_283),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_197),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_287),
.Y(n_315)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_187),
.Y(n_285)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_203),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_198),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_145),
.B(n_1),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_289),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_147),
.B(n_1),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_296),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_178),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_182),
.B(n_4),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_297),
.Y(n_318)
);

BUFx2_ASAP7_75t_SL g294 ( 
.A(n_180),
.Y(n_294)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_183),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_203),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_305),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_156),
.A2(n_4),
.B1(n_11),
.B2(n_12),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_301),
.A2(n_304),
.B1(n_309),
.B2(n_2),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_216),
.B(n_2),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_209),
.A2(n_2),
.B1(n_16),
.B2(n_164),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_169),
.B(n_16),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_158),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_307),
.Y(n_338)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_195),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_159),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_310),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_189),
.A2(n_2),
.B1(n_16),
.B2(n_170),
.Y(n_309)
);

INVx3_ASAP7_75t_SL g310 ( 
.A(n_228),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_165),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_311),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_252),
.A2(n_133),
.B(n_167),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_316),
.A2(n_333),
.B(n_307),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_369),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_324),
.A2(n_371),
.B1(n_291),
.B2(n_281),
.Y(n_401)
);

AOI32xp33_ASAP7_75t_L g330 ( 
.A1(n_235),
.A2(n_175),
.A3(n_194),
.B1(n_179),
.B2(n_184),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_251),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_248),
.B(n_261),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_331),
.B(n_349),
.C(n_351),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_252),
.A2(n_227),
.B(n_135),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_270),
.B(n_209),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_339),
.B(n_341),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_272),
.B(n_288),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_254),
.A2(n_202),
.B1(n_193),
.B2(n_177),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_342),
.A2(n_344),
.B1(n_345),
.B2(n_358),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_235),
.A2(n_260),
.B1(n_247),
.B2(n_255),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_289),
.A2(n_161),
.B1(n_154),
.B2(n_186),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_279),
.B(n_303),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_350),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_253),
.B(n_148),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_279),
.B(n_153),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_253),
.B(n_136),
.C(n_140),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_186),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_355),
.B(n_357),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_241),
.B(n_202),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_240),
.A2(n_228),
.B1(n_183),
.B2(n_141),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_359),
.A2(n_231),
.B1(n_245),
.B2(n_296),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_146),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_363),
.B(n_322),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_304),
.A2(n_146),
.B1(n_244),
.B2(n_280),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_310),
.B1(n_286),
.B2(n_300),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_242),
.B(n_146),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_280),
.A2(n_238),
.B1(n_243),
.B2(n_250),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_312),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_374),
.B(n_380),
.Y(n_423)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_314),
.B(n_262),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_377),
.B(n_382),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_319),
.A2(n_280),
.B1(n_277),
.B2(n_297),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_378),
.A2(n_383),
.B1(n_384),
.B2(n_391),
.Y(n_425)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_338),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_381),
.A2(n_411),
.B1(n_420),
.B2(n_353),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_367),
.B(n_298),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_371),
.A2(n_280),
.B1(n_257),
.B2(n_250),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_SL g457 ( 
.A(n_386),
.B(n_328),
.C(n_320),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_316),
.A2(n_299),
.B(n_302),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_387),
.A2(n_393),
.B(n_347),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_362),
.B(n_278),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_388),
.A2(n_390),
.B(n_405),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_372),
.Y(n_389)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_389),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_326),
.A2(n_233),
.B1(n_285),
.B2(n_283),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_404),
.B1(n_356),
.B2(n_369),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_346),
.A2(n_361),
.B(n_362),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_315),
.B(n_256),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_395),
.B(n_329),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_326),
.A2(n_233),
.B1(n_311),
.B2(n_236),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_396),
.B(n_410),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_400),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_401),
.A2(n_415),
.B1(n_416),
.B2(n_360),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_333),
.A2(n_264),
.B(n_258),
.Y(n_402)
);

OA22x2_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_325),
.B1(n_358),
.B2(n_360),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_339),
.A2(n_232),
.B1(n_246),
.B2(n_275),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_346),
.A2(n_232),
.B(n_273),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_331),
.B(n_230),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_363),
.C(n_347),
.Y(n_431)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_409),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_324),
.A2(n_290),
.B1(n_268),
.B2(n_295),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_418),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_320),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_334),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_313),
.A2(n_343),
.B1(n_341),
.B2(n_321),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_321),
.A2(n_335),
.B1(n_327),
.B2(n_318),
.Y(n_416)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_317),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_327),
.B(n_348),
.Y(n_418)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_364),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_332),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_349),
.B(n_351),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_422),
.A2(n_334),
.B(n_337),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_426),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_381),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_433),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_429),
.A2(n_419),
.B1(n_385),
.B2(n_431),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_430),
.A2(n_435),
.B(n_460),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_456),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_381),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_347),
.B(n_357),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_391),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_437),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_387),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_350),
.C(n_355),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_407),
.C(n_406),
.Y(n_468)
);

AO22x1_ASAP7_75t_L g440 ( 
.A1(n_378),
.A2(n_345),
.B1(n_364),
.B2(n_368),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_445),
.Y(n_481)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_410),
.A2(n_317),
.B1(n_323),
.B2(n_356),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_442),
.A2(n_413),
.B1(n_405),
.B2(n_420),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_449),
.B(n_376),
.Y(n_466)
);

OA22x2_ASAP7_75t_L g451 ( 
.A1(n_376),
.A2(n_368),
.B1(n_337),
.B2(n_332),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_396),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_381),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_452),
.B(n_453),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_394),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_462),
.C(n_389),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_402),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_366),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_459),
.B(n_463),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_393),
.A2(n_366),
.B(n_353),
.Y(n_460)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_419),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_461),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_464),
.B(n_472),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_465),
.A2(n_466),
.B1(n_469),
.B2(n_484),
.Y(n_511)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_424),
.Y(n_467)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_467),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_468),
.B(n_495),
.C(n_434),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_437),
.A2(n_383),
.B1(n_436),
.B2(n_425),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_423),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_425),
.A2(n_450),
.B1(n_435),
.B2(n_446),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_474),
.A2(n_482),
.B1(n_490),
.B2(n_494),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_462),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_475),
.B(n_476),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_432),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_427),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_477),
.B(n_480),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_479),
.A2(n_440),
.B(n_454),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_427),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_450),
.A2(n_446),
.B1(n_384),
.B2(n_398),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_487),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_451),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_398),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_497),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_458),
.A2(n_406),
.B1(n_403),
.B2(n_374),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_491),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_429),
.A2(n_402),
.B1(n_380),
.B2(n_403),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_422),
.C(n_400),
.Y(n_495)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_455),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_443),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_451),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_440),
.A2(n_397),
.B1(n_399),
.B2(n_412),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_498),
.A2(n_482),
.B1(n_474),
.B2(n_471),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_451),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_499),
.B(n_404),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_430),
.B(n_460),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_501),
.A2(n_443),
.B(n_447),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_456),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_509),
.Y(n_539)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_503),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_485),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_504),
.B(n_538),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_506),
.A2(n_514),
.B(n_528),
.Y(n_547)
);

AND3x1_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_426),
.C(n_457),
.Y(n_507)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_473),
.B(n_478),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g562 ( 
.A(n_508),
.B(n_527),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_438),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_447),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_510),
.A2(n_518),
.B1(n_524),
.B2(n_526),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_494),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_472),
.B(n_377),
.Y(n_513)
);

CKINVDCx14_ASAP7_75t_R g551 ( 
.A(n_513),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_426),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_516),
.B(n_533),
.C(n_534),
.Y(n_556)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_470),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_520),
.B(n_522),
.Y(n_546)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_491),
.Y(n_521)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_521),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_434),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_493),
.Y(n_523)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_523),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_489),
.A2(n_499),
.B1(n_497),
.B2(n_487),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_488),
.B(n_426),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_490),
.B(n_379),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_421),
.Y(n_554)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_493),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_531),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_453),
.C(n_454),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_486),
.B(n_375),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_535),
.B(n_492),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_466),
.A2(n_448),
.B1(n_444),
.B2(n_417),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_536),
.A2(n_469),
.B1(n_500),
.B2(n_483),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_481),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_470),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_510),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_541),
.B(n_548),
.Y(n_587)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_544),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_545),
.A2(n_555),
.B1(n_563),
.B2(n_433),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_547),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_529),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_519),
.A2(n_524),
.B1(n_517),
.B2(n_505),
.Y(n_549)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_549),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g550 ( 
.A1(n_511),
.A2(n_485),
.B(n_486),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_550),
.B(n_570),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_525),
.B(n_464),
.Y(n_552)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_552),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_517),
.A2(n_501),
.B(n_479),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_553),
.A2(n_506),
.B(n_536),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_559),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_505),
.A2(n_476),
.B1(n_475),
.B2(n_492),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_502),
.B(n_444),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_480),
.C(n_477),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_508),
.C(n_533),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_525),
.A2(n_537),
.B1(n_535),
.B2(n_519),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_448),
.Y(n_565)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_565),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_509),
.B(n_439),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_566),
.B(n_567),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_526),
.B(n_409),
.Y(n_568)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_568),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_522),
.B(n_439),
.Y(n_570)
);

AO22x1_ASAP7_75t_SL g572 ( 
.A1(n_540),
.A2(n_527),
.B1(n_507),
.B2(n_516),
.Y(n_572)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_572),
.Y(n_598)
);

FAx1_ASAP7_75t_SL g574 ( 
.A(n_560),
.B(n_562),
.CI(n_556),
.CON(n_574),
.SN(n_574)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_574),
.B(n_575),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_552),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_579),
.B(n_556),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_580),
.A2(n_569),
.B(n_561),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_555),
.A2(n_545),
.B1(n_563),
.B2(n_544),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_583),
.A2(n_588),
.B1(n_591),
.B2(n_592),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_547),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_584),
.A2(n_581),
.B(n_587),
.Y(n_614)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_543),
.Y(n_586)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_586),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_557),
.A2(n_534),
.B1(n_532),
.B2(n_515),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_558),
.B(n_532),
.Y(n_589)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_589),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_546),
.B(n_515),
.C(n_452),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_594),
.C(n_559),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_540),
.A2(n_428),
.B1(n_411),
.B2(n_408),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_546),
.B(n_411),
.C(n_329),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_596),
.B(n_600),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_584),
.A2(n_553),
.B(n_542),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_597),
.A2(n_606),
.B(n_608),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_615),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_539),
.C(n_566),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_590),
.B(n_539),
.C(n_567),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_602),
.B(n_612),
.C(n_600),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_583),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_611),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_577),
.A2(n_549),
.B(n_568),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_577),
.A2(n_551),
.B(n_565),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_609),
.A2(n_613),
.B(n_614),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_595),
.A2(n_564),
.B1(n_562),
.B2(n_554),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_610),
.A2(n_582),
.B1(n_593),
.B2(n_578),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_370),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_573),
.B(n_370),
.C(n_328),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_575),
.A2(n_580),
.B(n_581),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_SL g615 ( 
.A(n_576),
.B(n_573),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_616),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_599),
.B(n_576),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_619),
.B(n_620),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_595),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_622),
.B(n_612),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_613),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_623),
.B(n_627),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_601),
.A2(n_571),
.B1(n_592),
.B2(n_585),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_624),
.A2(n_607),
.B1(n_605),
.B2(n_606),
.Y(n_642)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_609),
.Y(n_625)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_625),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_589),
.Y(n_627)
);

MAJx2_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_604),
.C(n_608),
.Y(n_640)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_616),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_630),
.B(n_631),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_593),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_603),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_632),
.B(n_604),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_603),
.B(n_585),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_634),
.Y(n_644)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_637),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_645),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_642),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_629),
.A2(n_597),
.B(n_598),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_643),
.A2(n_633),
.B(n_639),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_629),
.A2(n_607),
.B1(n_571),
.B2(n_611),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_620),
.B(n_610),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_646),
.B(n_618),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_621),
.A2(n_598),
.B(n_574),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g659 ( 
.A1(n_647),
.A2(n_633),
.B(n_617),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_631),
.B(n_611),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_648),
.B(n_649),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_622),
.B(n_615),
.C(n_594),
.Y(n_649)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_650),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_651),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_638),
.B(n_636),
.C(n_649),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_655),
.A2(n_659),
.B(n_660),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_635),
.B(n_628),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g667 ( 
.A(n_656),
.B(n_658),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_641),
.B(n_626),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_636),
.B(n_626),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_654),
.B(n_644),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_661),
.A2(n_666),
.B(n_657),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_652),
.B(n_640),
.C(n_643),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_662),
.B(n_655),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_650),
.A2(n_646),
.B(n_645),
.Y(n_666)
);

AOI211xp5_ASAP7_75t_L g668 ( 
.A1(n_664),
.A2(n_663),
.B(n_667),
.C(n_665),
.Y(n_668)
);

AO21x2_ASAP7_75t_L g673 ( 
.A1(n_668),
.A2(n_670),
.B(n_671),
.Y(n_673)
);

AOI21xp33_ASAP7_75t_L g672 ( 
.A1(n_669),
.A2(n_627),
.B(n_634),
.Y(n_672)
);

NAND4xp25_ASAP7_75t_L g670 ( 
.A(n_661),
.B(n_657),
.C(n_653),
.D(n_617),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_672),
.A2(n_578),
.B(n_619),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_674),
.A2(n_673),
.B(n_582),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_675),
.A2(n_574),
.B(n_572),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_572),
.Y(n_677)
);


endmodule