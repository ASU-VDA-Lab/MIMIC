module real_jpeg_5754_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_1),
.Y(n_154)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_1),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_2),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_2),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_2),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_2),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_2),
.B(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_3),
.B(n_30),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_3),
.B(n_294),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_3),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_4),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_4),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_4),
.B(n_131),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_4),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_4),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_5),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_153),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_5),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_5),
.B(n_331),
.Y(n_330)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_8),
.B(n_156),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_8),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_8),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_9),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_9),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_9),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_9),
.B(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_10),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_10),
.Y(n_319)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_12),
.B(n_52),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_12),
.B(n_85),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_12),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_12),
.B(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_13),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_14),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_14),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_15),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_15),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_15),
.B(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_15),
.B(n_328),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_16),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_17),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_17),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_17),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_17),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_17),
.B(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_302),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_254),
.B(n_301),
.Y(n_19)
);

AOI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_214),
.B(n_253),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_162),
.B(n_213),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_123),
.B(n_161),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_89),
.B(n_122),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_66),
.B(n_88),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_44),
.B(n_65),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_37),
.B(n_43),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_35),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_42),
.Y(n_157)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_42),
.Y(n_192)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_56),
.C(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_64),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_87),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_87),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_73),
.C(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_72),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_106),
.C(n_107),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_82),
.Y(n_329)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_86),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_92),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_105),
.C(n_108),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_96),
.C(n_99),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_97),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_118),
.C(n_120),
.Y(n_159)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_116),
.Y(n_294)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_117),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_160),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_138),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_126),
.B(n_137),
.C(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_187),
.C(n_188),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_151),
.C(n_158),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_143),
.C(n_146),
.Y(n_184)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_145),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_148),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_158),
.B2(n_159),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_155),
.Y(n_183)
);

BUFx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_211),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_211),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_185),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_165),
.B(n_166),
.C(n_185),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_181),
.B2(n_182),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_231),
.C(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_174),
.C(n_180),
.Y(n_226)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_190),
.C(n_210),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_198),
.B1(n_209),
.B2(n_210),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_193),
.B(n_197),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.Y(n_197)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_197),
.B(n_218),
.C(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_199),
.B(n_206),
.C(n_207),
.Y(n_251)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_252),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_252),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_229),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_217),
.B(n_228),
.C(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_225),
.B2(n_227),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_220),
.B(n_223),
.C(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_224),
.Y(n_296)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_229),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_234),
.C(n_246),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_246),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_240),
.C(n_242),
.Y(n_268)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_250),
.C(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_251),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_299),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_282),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_259),
.B(n_267),
.C(n_270),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_260),
.B(n_262),
.C(n_264),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_274),
.C(n_279),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_274),
.Y(n_281)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_279),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_347),
.C(n_348),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_287),
.B1(n_297),
.B2(n_298),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_298),
.C(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_293),
.C(n_295),
.Y(n_336)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_349),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_346),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_346),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_333),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_320),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_316),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_345),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_338)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_339),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_341),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);


endmodule