module fake_jpeg_15804_n_56 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_56);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_56;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_7),
.B(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_15),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_9),
.A3(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_21),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_0),
.CON(n_28),
.SN(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_20),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_31),
.B1(n_5),
.B2(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_43),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_24),
.C(n_12),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_24),
.B1(n_11),
.B2(n_19),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_38),
.B1(n_48),
.B2(n_45),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

OAI21x1_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_50),
.B(n_51),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_55),
.Y(n_56)
);


endmodule