module real_aes_7197_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_140;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g445 ( .A1(n_0), .A2(n_145), .B(n_446), .C(n_449), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_1), .B(n_440), .Y(n_450) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g143 ( .A(n_3), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_4), .B(n_146), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_5), .A2(n_435), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_6), .A2(n_168), .B(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_7), .A2(n_39), .B1(n_133), .B2(n_191), .Y(n_231) );
AOI222xp33_ASAP7_75t_L g101 ( .A1(n_8), .A2(n_19), .B1(n_102), .B2(n_696), .C1(n_697), .C2(n_701), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_8), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_9), .B(n_168), .Y(n_176) );
AND2x6_ASAP7_75t_L g148 ( .A(n_10), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_11), .A2(n_148), .B(n_426), .C(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_12), .B(n_40), .Y(n_108) );
INVx1_ASAP7_75t_L g127 ( .A(n_13), .Y(n_127) );
INVx1_ASAP7_75t_L g124 ( .A(n_14), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_15), .B(n_129), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_16), .B(n_146), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_17), .B(n_120), .Y(n_178) );
AO32x2_ASAP7_75t_L g229 ( .A1(n_18), .A2(n_119), .A3(n_162), .B1(n_168), .B2(n_230), .Y(n_229) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_20), .A2(n_100), .B1(n_704), .B2(n_713), .C1(n_721), .C2(n_727), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g715 ( .A1(n_20), .A2(n_30), .B1(n_110), .B2(n_716), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_20), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_21), .B(n_133), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_22), .B(n_120), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_23), .A2(n_54), .B1(n_133), .B2(n_191), .Y(n_232) );
AOI22xp33_ASAP7_75t_SL g193 ( .A1(n_24), .A2(n_79), .B1(n_129), .B2(n_133), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_25), .B(n_133), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_26), .A2(n_162), .B(n_426), .C(n_457), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_27), .A2(n_162), .B(n_426), .C(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_28), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_29), .B(n_164), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_30), .A2(n_110), .B1(n_111), .B2(n_112), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_30), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_31), .A2(n_435), .B(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_32), .B(n_164), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_33), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g131 ( .A(n_34), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_35), .A2(n_432), .B(n_475), .C(n_476), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_36), .B(n_133), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_37), .B(n_164), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_38), .B(n_213), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_41), .B(n_455), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_42), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_43), .B(n_146), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_44), .B(n_435), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_45), .A2(n_432), .B(n_475), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_46), .B(n_133), .Y(n_171) );
INVx1_ASAP7_75t_L g447 ( .A(n_47), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_48), .A2(n_88), .B1(n_191), .B2(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g500 ( .A(n_49), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_50), .B(n_133), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_51), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_52), .B(n_435), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_53), .B(n_141), .Y(n_175) );
AOI22xp33_ASAP7_75t_SL g182 ( .A1(n_55), .A2(n_59), .B1(n_129), .B2(n_133), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_56), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_57), .B(n_133), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_58), .B(n_133), .Y(n_210) );
INVx1_ASAP7_75t_L g149 ( .A(n_60), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_61), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_62), .B(n_440), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_63), .A2(n_135), .B(n_141), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_64), .B(n_133), .Y(n_144) );
INVx1_ASAP7_75t_L g123 ( .A(n_65), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_66), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_67), .B(n_146), .Y(n_478) );
AO32x2_ASAP7_75t_L g188 ( .A1(n_68), .A2(n_162), .A3(n_168), .B1(n_189), .B2(n_194), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_69), .B(n_147), .Y(n_491) );
INVx1_ASAP7_75t_L g158 ( .A(n_70), .Y(n_158) );
INVx1_ASAP7_75t_L g201 ( .A(n_71), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_72), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_73), .B(n_459), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_74), .A2(n_426), .B(n_428), .C(n_432), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_75), .B(n_129), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_76), .Y(n_509) );
INVx1_ASAP7_75t_L g708 ( .A(n_77), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_78), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_80), .B(n_191), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_81), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_82), .B(n_129), .Y(n_205) );
INVx2_ASAP7_75t_L g121 ( .A(n_83), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_84), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_85), .B(n_161), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_86), .B(n_129), .Y(n_172) );
OR2x2_ASAP7_75t_L g105 ( .A(n_87), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g417 ( .A(n_87), .Y(n_417) );
OR2x2_ASAP7_75t_L g712 ( .A(n_87), .B(n_700), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_89), .A2(n_98), .B1(n_129), .B2(n_130), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_90), .B(n_435), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_91), .Y(n_477) );
INVxp67_ASAP7_75t_L g512 ( .A(n_92), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_93), .B(n_129), .Y(n_156) );
INVx1_ASAP7_75t_L g429 ( .A(n_94), .Y(n_429) );
INVx1_ASAP7_75t_L g487 ( .A(n_95), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_96), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g502 ( .A(n_97), .B(n_164), .Y(n_502) );
INVxp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_109), .B1(n_415), .B2(n_418), .Y(n_103) );
INVx2_ASAP7_75t_L g702 ( .A(n_104), .Y(n_702) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g416 ( .A(n_106), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g700 ( .A(n_106), .Y(n_700) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g701 ( .A1(n_109), .A2(n_418), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_111), .A2(n_112), .B1(n_715), .B2(n_717), .Y(n_714) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR5x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_306), .C(n_364), .D(n_400), .E(n_407), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_252), .C(n_276), .Y(n_113) );
AOI221xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_184), .B1(n_218), .B2(n_223), .C(n_233), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_115), .A2(n_387), .B(n_389), .Y(n_386) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_165), .Y(n_115) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_116), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_151), .Y(n_116) );
INVx2_ASAP7_75t_L g222 ( .A(n_117), .Y(n_222) );
AND2x2_ASAP7_75t_L g235 ( .A(n_117), .B(n_167), .Y(n_235) );
AND2x2_ASAP7_75t_L g289 ( .A(n_117), .B(n_166), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_117), .B(n_152), .Y(n_304) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_125), .B(n_150), .Y(n_117) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_118), .A2(n_153), .B(n_163), .Y(n_152) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_119), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_120), .Y(n_168) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_121), .B(n_122), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_139), .B(n_148), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_132), .C(n_135), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_128), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_128), .A2(n_520), .B(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
INVx1_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
INVx3_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_133), .Y(n_431) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
AND2x6_ASAP7_75t_L g426 ( .A(n_134), .B(n_427), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_L g428 ( .A1(n_135), .A2(n_429), .B(n_430), .C(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_136), .A2(n_204), .B(n_205), .Y(n_203) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g459 ( .A(n_137), .Y(n_459) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_138), .Y(n_161) );
INVx1_ASAP7_75t_L g213 ( .A(n_138), .Y(n_213) );
INVx1_ASAP7_75t_L g427 ( .A(n_138), .Y(n_427) );
AND2x2_ASAP7_75t_L g436 ( .A(n_138), .B(n_142), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_144), .C(n_145), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_L g157 ( .A1(n_140), .A2(n_158), .B(n_159), .C(n_160), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_140), .A2(n_458), .B(n_460), .Y(n_457) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_145), .A2(n_174), .B(n_175), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_145), .A2(n_161), .B1(n_181), .B2(n_182), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_145), .A2(n_161), .B1(n_231), .B2(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_146), .A2(n_155), .B(n_156), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_146), .A2(n_171), .B(n_172), .Y(n_170) );
O2A1O1Ixp5_ASAP7_75t_SL g199 ( .A1(n_146), .A2(n_200), .B(n_201), .C(n_202), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_146), .B(n_512), .Y(n_511) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g189 ( .A1(n_147), .A2(n_161), .B1(n_190), .B2(n_193), .Y(n_189) );
BUFx3_ASAP7_75t_L g162 ( .A(n_148), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_148), .A2(n_170), .B(n_173), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_148), .A2(n_199), .B(n_203), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_148), .A2(n_209), .B(n_214), .Y(n_208) );
INVx4_ASAP7_75t_SL g433 ( .A(n_148), .Y(n_433) );
AND2x4_ASAP7_75t_L g435 ( .A(n_148), .B(n_436), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g488 ( .A(n_148), .B(n_436), .Y(n_488) );
AND2x2_ASAP7_75t_L g322 ( .A(n_151), .B(n_263), .Y(n_322) );
AND2x2_ASAP7_75t_L g355 ( .A(n_151), .B(n_167), .Y(n_355) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OR2x2_ASAP7_75t_L g262 ( .A(n_152), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g275 ( .A(n_152), .B(n_167), .Y(n_275) );
AND2x2_ASAP7_75t_L g282 ( .A(n_152), .B(n_263), .Y(n_282) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_152), .Y(n_291) );
AND2x2_ASAP7_75t_L g298 ( .A(n_152), .B(n_166), .Y(n_298) );
INVx1_ASAP7_75t_L g329 ( .A(n_152), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_157), .B(n_162), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_160), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g448 ( .A(n_161), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g179 ( .A(n_162), .B(n_180), .C(n_183), .Y(n_179) );
INVx2_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_164), .A2(n_198), .B(n_206), .Y(n_197) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_164), .A2(n_208), .B(n_217), .Y(n_207) );
INVx1_ASAP7_75t_L g465 ( .A(n_164), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_164), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_164), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g305 ( .A(n_165), .Y(n_305) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_177), .Y(n_165) );
INVx2_ASAP7_75t_L g261 ( .A(n_166), .Y(n_261) );
AND2x2_ASAP7_75t_L g283 ( .A(n_166), .B(n_222), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_166), .B(n_329), .Y(n_334) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_167), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g406 ( .A(n_167), .B(n_370), .Y(n_406) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_176), .Y(n_167) );
INVx4_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_168), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_168), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g220 ( .A(n_177), .Y(n_220) );
INVx3_ASAP7_75t_L g321 ( .A(n_177), .Y(n_321) );
OR2x2_ASAP7_75t_L g351 ( .A(n_177), .B(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_177), .B(n_261), .Y(n_377) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g264 ( .A(n_178), .Y(n_264) );
AO21x1_ASAP7_75t_L g263 ( .A1(n_180), .A2(n_183), .B(n_264), .Y(n_263) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_183), .A2(n_424), .B(n_437), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_183), .B(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g440 ( .A(n_183), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_183), .B(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_183), .A2(n_486), .B(n_493), .Y(n_485) );
AOI33xp33_ASAP7_75t_L g397 ( .A1(n_184), .A2(n_235), .A3(n_249), .B1(n_321), .B2(n_398), .B3(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_195), .Y(n_185) );
OR2x2_ASAP7_75t_L g250 ( .A(n_186), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_186), .B(n_247), .Y(n_309) );
OR2x2_ASAP7_75t_L g362 ( .A(n_186), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g288 ( .A(n_187), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g313 ( .A(n_187), .B(n_195), .Y(n_313) );
AND2x2_ASAP7_75t_L g380 ( .A(n_187), .B(n_225), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_187), .A2(n_280), .B(n_406), .Y(n_405) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g227 ( .A(n_188), .Y(n_227) );
INVx1_ASAP7_75t_L g240 ( .A(n_188), .Y(n_240) );
AND2x2_ASAP7_75t_L g259 ( .A(n_188), .B(n_229), .Y(n_259) );
AND2x2_ASAP7_75t_L g308 ( .A(n_188), .B(n_228), .Y(n_308) );
INVx2_ASAP7_75t_L g449 ( .A(n_192), .Y(n_449) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_192), .Y(n_479) );
INVx1_ASAP7_75t_L g462 ( .A(n_194), .Y(n_462) );
INVx2_ASAP7_75t_SL g350 ( .A(n_195), .Y(n_350) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
INVx2_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
INVx1_ASAP7_75t_L g401 ( .A(n_196), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_196), .B(n_295), .Y(n_414) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g241 ( .A(n_197), .Y(n_241) );
OR2x2_ASAP7_75t_L g247 ( .A(n_197), .B(n_248), .Y(n_247) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_197), .Y(n_258) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_207), .Y(n_225) );
AND2x2_ASAP7_75t_L g242 ( .A(n_207), .B(n_228), .Y(n_242) );
INVx1_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
INVx1_ASAP7_75t_L g255 ( .A(n_207), .Y(n_255) );
AND2x2_ASAP7_75t_L g280 ( .A(n_207), .B(n_229), .Y(n_280) );
INVx2_ASAP7_75t_L g296 ( .A(n_207), .Y(n_296) );
AND2x2_ASAP7_75t_L g389 ( .A(n_207), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_207), .B(n_270), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g244 ( .A(n_220), .Y(n_244) );
INVx1_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_220), .B(n_304), .Y(n_370) );
INVx1_ASAP7_75t_SL g330 ( .A(n_221), .Y(n_330) );
INVx2_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
AND2x2_ASAP7_75t_L g320 ( .A(n_222), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g336 ( .A(n_222), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
INVx1_ASAP7_75t_L g398 ( .A(n_224), .Y(n_398) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g253 ( .A(n_226), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g356 ( .A(n_226), .B(n_346), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_226), .A2(n_367), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_L g269 ( .A(n_227), .B(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
INVx1_ASAP7_75t_L g318 ( .A(n_227), .Y(n_318) );
OR2x2_ASAP7_75t_L g382 ( .A(n_228), .B(n_241), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_228), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g295 ( .A(n_229), .B(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g302 ( .A(n_229), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_236), .B1(n_243), .B2(n_245), .Y(n_233) );
OR2x2_ASAP7_75t_L g312 ( .A(n_234), .B(n_262), .Y(n_312) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_235), .A2(n_354), .B1(n_356), .B2(n_357), .C1(n_358), .C2(n_361), .Y(n_353) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_242), .Y(n_237) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g300 ( .A(n_239), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_241), .B(n_255), .Y(n_254) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
AND2x2_ASAP7_75t_L g373 ( .A(n_241), .B(n_242), .Y(n_373) );
INVx1_ASAP7_75t_L g391 ( .A(n_241), .Y(n_391) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g357 ( .A(n_244), .B(n_283), .Y(n_357) );
AND2x2_ASAP7_75t_L g399 ( .A(n_244), .B(n_275), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_246), .B(n_294), .Y(n_381) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_247), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g274 ( .A(n_251), .B(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g342 ( .A(n_251), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .B(n_260), .C(n_265), .Y(n_252) );
INVxp67_ASAP7_75t_L g266 ( .A(n_253), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_254), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_254), .B(n_301), .Y(n_396) );
BUFx3_ASAP7_75t_L g360 ( .A(n_255), .Y(n_360) );
INVx1_ASAP7_75t_L g267 ( .A(n_256), .Y(n_267) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g286 ( .A(n_258), .B(n_280), .Y(n_286) );
INVx1_ASAP7_75t_SL g326 ( .A(n_259), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
AND2x2_ASAP7_75t_L g339 ( .A(n_261), .B(n_322), .Y(n_339) );
INVx1_ASAP7_75t_SL g310 ( .A(n_262), .Y(n_310) );
INVx1_ASAP7_75t_L g337 ( .A(n_263), .Y(n_337) );
AOI31xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .A3(n_268), .B(n_271), .Y(n_265) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g358 ( .A(n_269), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g332 ( .A(n_270), .Y(n_332) );
BUFx2_ASAP7_75t_L g346 ( .A(n_270), .Y(n_346) );
AND2x2_ASAP7_75t_L g374 ( .A(n_270), .B(n_295), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g347 ( .A(n_274), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_275), .B(n_342), .Y(n_388) );
AND2x2_ASAP7_75t_L g395 ( .A(n_275), .B(n_321), .Y(n_395) );
AOI211xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B(n_284), .C(n_299), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_281), .A2(n_308), .B1(n_309), .B2(n_310), .C(n_311), .Y(n_307) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g315 ( .A(n_282), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
OAI32xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .A3(n_290), .B1(n_292), .B2(n_297), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_286), .A2(n_339), .B(n_340), .C(n_343), .Y(n_338) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
OAI21xp5_ASAP7_75t_SL g402 ( .A1(n_294), .A2(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g363 ( .A(n_295), .Y(n_363) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_301), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g349 ( .A(n_301), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NAND4xp25_ASAP7_75t_SL g306 ( .A(n_307), .B(n_319), .C(n_338), .D(n_353), .Y(n_306) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g367 ( .A(n_308), .B(n_360), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_310), .B(n_342), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_314), .B2(n_317), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_312), .A2(n_363), .B1(n_394), .B2(n_396), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_312), .A2(n_401), .B(n_402), .C(n_405), .Y(n_400) );
INVx2_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_349), .B1(n_366), .B2(n_367), .C1(n_368), .C2(n_371), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_322), .B(n_323), .C(n_327), .Y(n_319) );
INVx1_ASAP7_75t_L g385 ( .A(n_320), .Y(n_385) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_324), .A2(n_328), .B1(n_331), .B2(n_333), .Y(n_327) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g354 ( .A(n_336), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g412 ( .A(n_339), .Y(n_412) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B1(n_348), .B2(n_351), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_346), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g403 ( .A(n_351), .Y(n_403) );
INVx1_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_357), .Y(n_411) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND5xp2_ASAP7_75t_L g364 ( .A(n_365), .B(n_372), .C(n_386), .D(n_392), .E(n_397), .Y(n_364) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_375), .C(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI31xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .A3(n_382), .B(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g404 ( .A(n_380), .Y(n_404) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI222xp33_ASAP7_75t_L g407 ( .A1(n_394), .A2(n_396), .B1(n_408), .B2(n_411), .C1(n_412), .C2(n_413), .Y(n_407) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g703 ( .A(n_415), .Y(n_703) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR2x2_ASAP7_75t_L g699 ( .A(n_417), .B(n_700), .Y(n_699) );
OR3x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_604), .C(n_653), .Y(n_418) );
NAND5xp2_ASAP7_75t_L g419 ( .A(n_420), .B(n_538), .C(n_567), .D(n_575), .E(n_590), .Y(n_419) );
O2A1O1Ixp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_466), .B(n_482), .C(n_522), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_451), .Y(n_421) );
AND2x2_ASAP7_75t_L g533 ( .A(n_422), .B(n_530), .Y(n_533) );
AND2x2_ASAP7_75t_L g566 ( .A(n_422), .B(n_452), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_422), .B(n_470), .Y(n_659) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_439), .Y(n_422) );
INVx2_ASAP7_75t_L g469 ( .A(n_423), .Y(n_469) );
BUFx2_ASAP7_75t_L g633 ( .A(n_423), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_434), .Y(n_424) );
INVx5_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_SL g442 ( .A1(n_433), .A2(n_443), .B(n_444), .C(n_445), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_433), .A2(n_444), .B(n_509), .C(n_510), .Y(n_508) );
BUFx2_ASAP7_75t_L g455 ( .A(n_435), .Y(n_455) );
AND2x2_ASAP7_75t_L g451 ( .A(n_439), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g531 ( .A(n_439), .Y(n_531) );
AND2x2_ASAP7_75t_L g617 ( .A(n_439), .B(n_530), .Y(n_617) );
AND2x2_ASAP7_75t_L g672 ( .A(n_439), .B(n_469), .Y(n_672) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_450), .Y(n_439) );
INVx2_ASAP7_75t_L g475 ( .A(n_444), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g589 ( .A(n_451), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_451), .B(n_470), .Y(n_636) );
INVx5_ASAP7_75t_L g530 ( .A(n_452), .Y(n_530) );
AND2x4_ASAP7_75t_L g551 ( .A(n_452), .B(n_531), .Y(n_551) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_452), .Y(n_573) );
AND2x2_ASAP7_75t_L g648 ( .A(n_452), .B(n_633), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_452), .B(n_471), .Y(n_651) );
OR2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
AOI21xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_456), .B(n_462), .Y(n_453) );
INVx2_ASAP7_75t_L g461 ( .A(n_459), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_461), .A2(n_477), .B(n_478), .C(n_479), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_461), .A2(n_479), .B(n_500), .C(n_501), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_466), .B(n_531), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_466), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
AND2x2_ASAP7_75t_L g556 ( .A(n_468), .B(n_531), .Y(n_556) );
AND2x2_ASAP7_75t_L g574 ( .A(n_468), .B(n_471), .Y(n_574) );
INVx1_ASAP7_75t_L g594 ( .A(n_468), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_468), .B(n_530), .Y(n_639) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_468), .Y(n_681) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_469), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_470), .B(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_470), .Y(n_583) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_470), .A2(n_526), .B(n_587), .C(n_589), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_470), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g602 ( .A(n_470), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g606 ( .A(n_470), .B(n_530), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_470), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g621 ( .A(n_470), .B(n_531), .Y(n_621) );
AND2x2_ASAP7_75t_L g671 ( .A(n_470), .B(n_672), .Y(n_671) );
INVx5_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g535 ( .A(n_471), .Y(n_535) );
AND2x2_ASAP7_75t_L g576 ( .A(n_471), .B(n_529), .Y(n_576) );
AND2x2_ASAP7_75t_L g588 ( .A(n_471), .B(n_563), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_471), .B(n_617), .Y(n_635) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .Y(n_471) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_503), .Y(n_482) );
INVx1_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_495), .Y(n_483) );
OR2x2_ASAP7_75t_L g526 ( .A(n_484), .B(n_495), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_484), .B(n_533), .C(n_534), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_484), .B(n_505), .Y(n_543) );
OR2x2_ASAP7_75t_L g558 ( .A(n_484), .B(n_546), .Y(n_558) );
AND2x2_ASAP7_75t_L g564 ( .A(n_484), .B(n_514), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_484), .B(n_695), .Y(n_694) );
INVx5_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_485), .B(n_505), .Y(n_561) );
AND2x2_ASAP7_75t_L g600 ( .A(n_485), .B(n_515), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_485), .B(n_514), .Y(n_628) );
OR2x2_ASAP7_75t_L g631 ( .A(n_485), .B(n_514), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_489), .Y(n_486) );
INVx5_ASAP7_75t_SL g546 ( .A(n_495), .Y(n_546) );
OR2x2_ASAP7_75t_L g552 ( .A(n_495), .B(n_504), .Y(n_552) );
AND2x2_ASAP7_75t_L g568 ( .A(n_495), .B(n_569), .Y(n_568) );
AOI321xp33_ASAP7_75t_L g575 ( .A1(n_495), .A2(n_576), .A3(n_577), .B1(n_578), .B2(n_584), .C(n_586), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_495), .B(n_503), .Y(n_585) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_495), .Y(n_598) );
OR2x2_ASAP7_75t_L g645 ( .A(n_495), .B(n_543), .Y(n_645) );
AND2x2_ASAP7_75t_L g667 ( .A(n_495), .B(n_564), .Y(n_667) );
AND2x2_ASAP7_75t_L g686 ( .A(n_495), .B(n_505), .Y(n_686) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_514), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_505), .B(n_514), .Y(n_527) );
AND2x2_ASAP7_75t_L g536 ( .A(n_505), .B(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
AND2x2_ASAP7_75t_L g569 ( .A(n_505), .B(n_564), .Y(n_569) );
INVxp67_ASAP7_75t_L g599 ( .A(n_505), .Y(n_599) );
OR2x2_ASAP7_75t_L g641 ( .A(n_505), .B(n_546), .Y(n_641) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_513), .Y(n_505) );
OR2x2_ASAP7_75t_L g523 ( .A(n_514), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_SL g537 ( .A(n_514), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_514), .B(n_526), .Y(n_570) );
AND2x2_ASAP7_75t_L g619 ( .A(n_514), .B(n_563), .Y(n_619) );
AND2x2_ASAP7_75t_L g657 ( .A(n_514), .B(n_546), .Y(n_657) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_515), .B(n_546), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_525), .B(n_528), .C(n_532), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_523), .A2(n_525), .B1(n_650), .B2(n_652), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_525), .A2(n_548), .B1(n_603), .B2(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_SL g677 ( .A(n_526), .Y(n_677) );
INVx1_ASAP7_75t_SL g577 ( .A(n_527), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_529), .B(n_549), .Y(n_579) );
AOI222xp33_ASAP7_75t_L g590 ( .A1(n_529), .A2(n_570), .B1(n_577), .B2(n_591), .C1(n_595), .C2(n_601), .Y(n_590) );
AND2x2_ASAP7_75t_L g680 ( .A(n_529), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g555 ( .A(n_530), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_530), .B(n_550), .Y(n_625) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_530), .Y(n_662) );
AND2x2_ASAP7_75t_L g665 ( .A(n_530), .B(n_574), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_530), .B(n_681), .Y(n_691) );
INVx1_ASAP7_75t_L g582 ( .A(n_531), .Y(n_582) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_531), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_533), .A2(n_674), .B(n_675), .C(n_678), .Y(n_673) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_535), .B(n_597), .C(n_600), .Y(n_596) );
OR2x2_ASAP7_75t_L g624 ( .A(n_535), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_535), .B(n_551), .Y(n_652) );
OR2x2_ASAP7_75t_L g557 ( .A(n_537), .B(n_558), .Y(n_557) );
AOI211xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_541), .B(n_547), .C(n_559), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_540), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g646 ( .A(n_541), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_542), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g560 ( .A(n_545), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_546), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g614 ( .A(n_546), .B(n_564), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_546), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_546), .B(n_563), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_552), .B1(n_553), .B2(n_557), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_549), .B(n_621), .Y(n_620) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_551), .B(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_552), .A2(n_616), .B1(n_618), .B2(n_620), .C(n_622), .Y(n_615) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g670 ( .A(n_555), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g683 ( .A(n_555), .B(n_672), .Y(n_683) );
INVx1_ASAP7_75t_L g603 ( .A(n_556), .Y(n_603) );
INVx1_ASAP7_75t_L g674 ( .A(n_557), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_558), .A2(n_641), .B(n_664), .Y(n_663) );
AOI21xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_562), .B(n_565), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_570), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g607 ( .A(n_568), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_569), .A2(n_655), .B1(n_658), .B2(n_660), .C(n_663), .Y(n_654) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_577), .A2(n_667), .B1(n_668), .B2(n_670), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g643 ( .A(n_579), .Y(n_643) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp67_ASAP7_75t_SL g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_L g647 ( .A(n_583), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g612 ( .A(n_588), .Y(n_612) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_593), .B(n_617), .Y(n_669) );
INVxp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_599), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g685 ( .A(n_600), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g692 ( .A(n_600), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI211xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B(n_608), .C(n_642), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B(n_615), .C(n_634), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g695 ( .A(n_619), .Y(n_695) );
AND2x2_ASAP7_75t_L g632 ( .A(n_621), .B(n_633), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_630), .B2(n_632), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g640 ( .A(n_628), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g693 ( .A(n_629), .Y(n_693) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI31xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .A3(n_637), .B(n_640), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_646), .C(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
CKINVDCx16_ASAP7_75t_R g650 ( .A(n_651), .Y(n_650) );
NAND5xp2_ASAP7_75t_L g653 ( .A(n_654), .B(n_666), .C(n_673), .D(n_687), .E(n_690), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_665), .A2(n_691), .B1(n_692), .B2(n_694), .Y(n_690) );
INVx1_ASAP7_75t_SL g689 ( .A(n_667), .Y(n_689) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .B(n_684), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .Y(n_705) );
NOR2xp33_ASAP7_75t_SL g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g726 ( .A(n_707), .Y(n_726) );
INVx1_ASAP7_75t_L g725 ( .A(n_709), .Y(n_725) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_709), .A2(n_720), .B(n_726), .Y(n_728) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_711), .A2(n_714), .B(n_718), .Y(n_713) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g720 ( .A(n_712), .Y(n_720) );
INVx1_ASAP7_75t_L g717 ( .A(n_715), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
CKINVDCx6p67_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
endmodule