module fake_jpeg_1053_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_44),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_51),
.B1(n_46),
.B2(n_41),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_70),
.B1(n_47),
.B2(n_38),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_46),
.B1(n_41),
.B2(n_47),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_50),
.B1(n_40),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_50),
.B1(n_42),
.B2(n_56),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_77),
.B(n_4),
.Y(n_98)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_49),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_1),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_83),
.B1(n_19),
.B2(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_18),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_68),
.B1(n_64),
.B2(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_67),
.B1(n_53),
.B2(n_52),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_17),
.C(n_28),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_49),
.B1(n_62),
.B2(n_6),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_96),
.B1(n_13),
.B2(n_14),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_4),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_100),
.B(n_11),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_20),
.Y(n_104)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_21),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_7),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_112),
.C(n_92),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_8),
.B(n_10),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_93),
.B1(n_16),
.B2(n_26),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_8),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_88),
.C(n_13),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_11),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_24),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_108),
.B1(n_107),
.B2(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_137),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_129),
.B(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_120),
.B(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_132),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_142),
.B(n_143),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_135),
.C(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_145),
.A2(n_134),
.B1(n_137),
.B2(n_123),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_147),
.A2(n_122),
.B(n_103),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_150),
.C(n_148),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_122),
.B(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_15),
.B(n_27),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_37),
.Y(n_156)
);


endmodule