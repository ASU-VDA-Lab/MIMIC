module fake_jpeg_30746_n_537 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_537);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_1),
.B(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_21),
.B(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_81),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_21),
.B(n_14),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_92),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_36),
.B(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_14),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_93),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_50),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_50),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_109),
.B(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_115),
.B(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_49),
.B1(n_47),
.B2(n_51),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_118),
.A2(n_131),
.B1(n_160),
.B2(n_34),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_87),
.A2(n_26),
.B1(n_17),
.B2(n_48),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_32),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_77),
.B(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_141),
.B(n_153),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_90),
.A2(n_51),
.B1(n_44),
.B2(n_26),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_48),
.B1(n_43),
.B2(n_44),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_60),
.B(n_19),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_155),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_46),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_62),
.A2(n_33),
.B(n_32),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_62),
.A2(n_33),
.B(n_32),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_51),
.Y(n_184)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_68),
.A2(n_51),
.B1(n_44),
.B2(n_19),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_70),
.B(n_34),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_86),
.B1(n_69),
.B2(n_85),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_164),
.A2(n_166),
.B1(n_193),
.B2(n_196),
.Y(n_217)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_165),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_114),
.B1(n_64),
.B2(n_74),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_167),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_171),
.A2(n_192),
.B1(n_194),
.B2(n_30),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_176),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_104),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_177),
.Y(n_253)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_178),
.B(n_181),
.Y(n_243)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_180),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_108),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_186),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_89),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_105),
.B(n_97),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_102),
.B1(n_100),
.B2(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_135),
.A2(n_96),
.B1(n_95),
.B2(n_94),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_195),
.A2(n_151),
.B1(n_144),
.B2(n_121),
.Y(n_238)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_230)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_114),
.A2(n_56),
.B1(n_61),
.B2(n_63),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

AO22x2_ASAP7_75t_L g201 ( 
.A1(n_135),
.A2(n_88),
.B1(n_83),
.B2(n_82),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_211),
.B1(n_213),
.B2(n_137),
.Y(n_232)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_113),
.A2(n_17),
.B1(n_16),
.B2(n_30),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_127),
.B1(n_149),
.B2(n_162),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_120),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_128),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_212),
.Y(n_233)
);

NAND2x1_ASAP7_75t_SL g210 ( 
.A(n_131),
.B(n_43),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_137),
.B(n_151),
.Y(n_219)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_128),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_219),
.A2(n_182),
.B(n_156),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_184),
.B(n_117),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_227),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_107),
.B1(n_116),
.B2(n_148),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_240),
.B1(n_246),
.B2(n_205),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_226),
.A2(n_189),
.B1(n_211),
.B2(n_207),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_184),
.B(n_28),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_138),
.B(n_127),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_231),
.A2(n_236),
.B(n_0),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_232),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_208),
.B1(n_209),
.B2(n_190),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_250),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_186),
.A2(n_30),
.B(n_16),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_144),
.B1(n_148),
.B2(n_107),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_171),
.A2(n_116),
.B1(n_162),
.B2(n_121),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_154),
.B1(n_43),
.B2(n_134),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_163),
.B(n_46),
.C(n_45),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_201),
.A2(n_154),
.B1(n_134),
.B2(n_20),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_254),
.A2(n_268),
.B1(n_237),
.B2(n_273),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_217),
.B1(n_230),
.B2(n_226),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_186),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_259),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_189),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_244),
.A2(n_172),
.B1(n_185),
.B2(n_179),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_260),
.A2(n_285),
.B1(n_289),
.B2(n_245),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_223),
.B1(n_245),
.B2(n_221),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_180),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_227),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_170),
.B1(n_177),
.B2(n_202),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_264),
.A2(n_216),
.B1(n_232),
.B2(n_241),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_165),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_265),
.B(n_269),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_213),
.C(n_203),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_276),
.C(n_232),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_169),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_274),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_197),
.B1(n_187),
.B2(n_200),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_188),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_288),
.B(n_241),
.Y(n_292)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_198),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_220),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_275),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_196),
.C(n_173),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_28),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_38),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_279),
.Y(n_324)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

AO22x2_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_222),
.B1(n_253),
.B2(n_251),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_231),
.A2(n_42),
.B(n_38),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_287),
.B(n_245),
.Y(n_301)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_214),
.A2(n_146),
.B1(n_42),
.B2(n_43),
.Y(n_285)
);

AOI32xp33_ASAP7_75t_L g286 ( 
.A1(n_219),
.A2(n_45),
.A3(n_43),
.B1(n_10),
.B2(n_3),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_238),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_215),
.A2(n_10),
.B(n_1),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_214),
.A2(n_43),
.B1(n_10),
.B2(n_2),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_236),
.B(n_10),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_216),
.B1(n_237),
.B2(n_241),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_321),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_293),
.A2(n_307),
.B1(n_313),
.B2(n_314),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_232),
.B(n_235),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_294),
.A2(n_282),
.B(n_283),
.Y(n_344)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_279),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_300),
.A2(n_309),
.B1(n_275),
.B2(n_255),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_302),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_259),
.B(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_266),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_273),
.A2(n_223),
.B1(n_235),
.B2(n_221),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_308),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_247),
.B1(n_229),
.B2(n_248),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_311),
.A2(n_264),
.B1(n_260),
.B2(n_278),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_254),
.A2(n_223),
.B1(n_221),
.B2(n_248),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_247),
.B(n_229),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_251),
.C(n_253),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_276),
.C(n_262),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_304),
.B(n_281),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_327),
.B(n_345),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_328),
.B(n_340),
.C(n_332),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_301),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_337),
.B1(n_346),
.B2(n_302),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_263),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_325),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_339),
.B1(n_343),
.B2(n_348),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_257),
.B(n_290),
.Y(n_336)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_349),
.C(n_310),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_323),
.A2(n_256),
.B1(n_261),
.B2(n_266),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_294),
.A2(n_267),
.B1(n_256),
.B2(n_261),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_291),
.A2(n_267),
.B1(n_269),
.B2(n_288),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_315),
.B(n_303),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_304),
.B(n_277),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_323),
.A2(n_257),
.B1(n_276),
.B2(n_282),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_222),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_300),
.A2(n_270),
.B1(n_248),
.B2(n_285),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_350),
.A2(n_356),
.B1(n_311),
.B2(n_319),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_252),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_352),
.Y(n_386)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_309),
.A2(n_222),
.B1(n_252),
.B2(n_289),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_312),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_357),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_312),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_358),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_297),
.B(n_252),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_312),
.Y(n_377)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_360),
.A2(n_292),
.B(n_306),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_362),
.A2(n_368),
.B(n_371),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_363),
.B(n_364),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_360),
.A2(n_338),
.B(n_347),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_379),
.B(n_389),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_338),
.A2(n_320),
.B(n_302),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_338),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_376),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_342),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_384),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_303),
.Y(n_378)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_344),
.A2(n_295),
.B(n_310),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_351),
.A2(n_331),
.B1(n_337),
.B2(n_347),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_388),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_381),
.A2(n_395),
.B1(n_334),
.B2(n_339),
.Y(n_396)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

XOR2x2_ASAP7_75t_SL g387 ( 
.A(n_343),
.B(n_296),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_387),
.B(n_361),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_346),
.A2(n_296),
.B1(n_305),
.B2(n_293),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_344),
.A2(n_322),
.B(n_321),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_390),
.A2(n_335),
.B1(n_342),
.B2(n_353),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_357),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_358),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_318),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_393),
.C(n_394),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_317),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_330),
.A2(n_321),
.B1(n_319),
.B2(n_308),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_396),
.A2(n_398),
.B1(n_421),
.B2(n_369),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_381),
.A2(n_350),
.B1(n_356),
.B2(n_341),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_379),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_329),
.Y(n_403)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_329),
.Y(n_404)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_366),
.B(n_354),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_405),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_365),
.B(n_321),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_418),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_321),
.Y(n_413)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_414),
.A2(n_389),
.B1(n_388),
.B2(n_380),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_353),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_335),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_424),
.Y(n_426)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_372),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_420),
.A2(n_422),
.B1(n_423),
.B2(n_400),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_395),
.A2(n_326),
.B1(n_1),
.B2(n_2),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_370),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_326),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_373),
.A2(n_0),
.B(n_1),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_425),
.A2(n_371),
.B(n_391),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_398),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_363),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_429),
.B(n_430),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_392),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_431),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_409),
.A2(n_413),
.B1(n_412),
.B2(n_422),
.Y(n_432)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_417),
.B(n_394),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_434),
.B(n_435),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_393),
.Y(n_435)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_440),
.B(n_397),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_362),
.C(n_364),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_445),
.C(n_448),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_415),
.A2(n_387),
.B1(n_385),
.B2(n_383),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_415),
.A2(n_375),
.B1(n_376),
.B2(n_391),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_444),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_412),
.A2(n_375),
.B1(n_368),
.B2(n_2),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_0),
.C(n_1),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_0),
.C(n_3),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_396),
.B(n_3),
.C(n_4),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_449),
.B(n_399),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_451),
.B(n_458),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_406),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_454),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_406),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_406),
.C(n_419),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_456),
.B(n_460),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_436),
.B(n_400),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_457),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_406),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_414),
.C(n_402),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_427),
.B(n_397),
.C(n_405),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_464),
.B(n_438),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_404),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_426),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_470),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_426),
.C(n_439),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_488),
.C(n_455),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_466),
.A2(n_447),
.B1(n_450),
.B2(n_432),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_399),
.B1(n_445),
.B2(n_448),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_463),
.A2(n_437),
.B1(n_446),
.B2(n_436),
.Y(n_474)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_474),
.Y(n_503)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_475),
.B(n_479),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_453),
.A2(n_446),
.B1(n_447),
.B2(n_428),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_482),
.Y(n_498)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_468),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_483),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_444),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_487),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_462),
.A2(n_431),
.B(n_450),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_485),
.A2(n_486),
.B(n_473),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_428),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_401),
.C(n_403),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_500),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_490),
.B(n_495),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_451),
.B1(n_421),
.B2(n_454),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_491),
.A2(n_493),
.B1(n_481),
.B2(n_486),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_485),
.A2(n_458),
.B1(n_452),
.B2(n_407),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_459),
.C(n_455),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_497),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_418),
.B(n_407),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_459),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_423),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_420),
.C(n_449),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_410),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_424),
.B(n_7),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_481),
.C(n_484),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_472),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_507),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_472),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_508),
.B(n_513),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_497),
.C(n_496),
.Y(n_520)
);

FAx1_ASAP7_75t_SL g510 ( 
.A(n_490),
.B(n_410),
.CI(n_425),
.CON(n_510),
.SN(n_510)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_510),
.B(n_493),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_501),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_512),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_6),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_499),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_516),
.A2(n_492),
.B(n_503),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_517),
.A2(n_518),
.B(n_520),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_514),
.A2(n_515),
.B(n_511),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_522),
.A2(n_6),
.B(n_7),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_505),
.A2(n_491),
.B1(n_495),
.B2(n_8),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_SL g525 ( 
.A1(n_524),
.A2(n_512),
.B(n_514),
.C(n_8),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_527),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_521),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_7),
.C(n_8),
.Y(n_527)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_530),
.B(n_524),
.C(n_8),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_519),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_531),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_533),
.B(n_7),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_7),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_9),
.Y(n_536)
);

AO21x1_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_9),
.B(n_529),
.Y(n_537)
);


endmodule