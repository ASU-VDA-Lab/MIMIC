module fake_jpeg_20592_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_31),
.Y(n_38)
);

CKINVDCx9p33_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_15),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_18),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_21),
.B1(n_14),
.B2(n_11),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_27),
.B1(n_21),
.B2(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_55),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_30),
.B(n_31),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_58),
.C(n_2),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_19),
.B1(n_21),
.B2(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_38),
.B1(n_32),
.B2(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_19),
.B1(n_12),
.B2(n_17),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_17),
.B(n_19),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_43),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_20),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_66),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_3),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_57),
.B(n_58),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_7),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_10),
.B(n_9),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_53),
.C(n_51),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_3),
.C(n_4),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_51),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_49),
.B1(n_48),
.B2(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_79),
.B1(n_62),
.B2(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_50),
.B1(n_56),
.B2(n_5),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_87),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_82),
.B1(n_76),
.B2(n_73),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_63),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_80),
.B(n_81),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_81),
.C(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_61),
.C(n_8),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_73),
.B1(n_6),
.B2(n_4),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_87),
.B1(n_84),
.B2(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

AOI31xp33_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_96),
.A3(n_89),
.B(n_9),
.Y(n_102)
);

OAI21x1_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_4),
.B(n_99),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_101),
.Y(n_104)
);


endmodule