module fake_jpeg_18650_n_59 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_7),
.B(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_26),
.B1(n_3),
.B2(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_45),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_26),
.A3(n_24),
.B1(n_5),
.B2(n_6),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_13),
.Y(n_50)
);

AO21x2_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_2),
.B(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_17),
.B1(n_8),
.B2(n_11),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_23),
.B1(n_14),
.B2(n_15),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_19),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_49),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.C(n_41),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_44),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_46),
.B2(n_20),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_51),
.C(n_46),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_18),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_21),
.Y(n_57)
);

BUFx24_ASAP7_75t_SL g58 ( 
.A(n_57),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_22),
.Y(n_59)
);


endmodule