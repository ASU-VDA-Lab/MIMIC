module fake_jpeg_25823_n_264 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx13_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx8_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_30),
.Y(n_44)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_11),
.B1(n_12),
.B2(n_20),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g34 ( 
.A(n_14),
.B(n_18),
.CON(n_34),
.SN(n_34)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_11),
.B1(n_16),
.B2(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_31),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_27),
.B1(n_28),
.B2(n_11),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_59),
.B1(n_43),
.B2(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_49),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_32),
.C(n_29),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.C(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_35),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_26),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_14),
.B(n_18),
.C(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_15),
.Y(n_96)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_12),
.B1(n_40),
.B2(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_33),
.B1(n_30),
.B2(n_12),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_55),
.C(n_37),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_84),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_53),
.B1(n_59),
.B2(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_92),
.B1(n_90),
.B2(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_55),
.B(n_56),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_90),
.B(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_12),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_25),
.C(n_40),
.Y(n_118)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_37),
.B1(n_55),
.B2(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_2),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_15),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_37),
.B1(n_50),
.B2(n_57),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_101),
.B1(n_114),
.B2(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_37),
.B1(n_39),
.B2(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_104),
.B(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_115),
.B1(n_76),
.B2(n_20),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_29),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_24),
.B(n_48),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_39),
.B1(n_20),
.B2(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_116),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_141),
.B1(n_39),
.B2(n_66),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_89),
.C(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_127),
.C(n_129),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_124),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_24),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_92),
.C(n_79),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_136),
.B1(n_101),
.B2(n_109),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_77),
.C(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_135),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_70),
.B1(n_76),
.B2(n_78),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_39),
.B1(n_52),
.B2(n_40),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_78),
.B1(n_75),
.B2(n_62),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_100),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_145),
.B(n_147),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_20),
.B1(n_75),
.B2(n_65),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_48),
.Y(n_145)
);

XOR2x1_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_10),
.Y(n_147)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_167),
.B1(n_132),
.B2(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_166),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_21),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_162),
.C(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_61),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_61),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_77),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_77),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_39),
.B1(n_52),
.B2(n_40),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_132),
.B1(n_143),
.B2(n_137),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_58),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_140),
.C(n_122),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_147),
.B(n_126),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_151),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_178),
.B(n_149),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_145),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_131),
.B(n_146),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_187),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_190),
.B1(n_171),
.B2(n_166),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_200),
.B1(n_204),
.B2(n_188),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_155),
.B1(n_164),
.B2(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_202),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_164),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_205),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_170),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_158),
.C(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_178),
.C(n_190),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_154),
.B1(n_157),
.B2(n_161),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_178),
.B(n_182),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_149),
.B1(n_137),
.B2(n_23),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_58),
.B1(n_23),
.B2(n_25),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_210),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_215),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_186),
.B1(n_180),
.B2(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_218),
.C(n_214),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_219),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_21),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_203),
.B1(n_192),
.B2(n_201),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_184),
.B1(n_23),
.B2(n_13),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_16),
.B1(n_22),
.B2(n_19),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_19),
.C(n_21),
.Y(n_231)
);

OAI21x1_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_196),
.B(n_9),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_226),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_215),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_195),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_231),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_21),
.C(n_19),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_213),
.C(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_19),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_235),
.C(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_219),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_220),
.B(n_22),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_2),
.B(n_3),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_22),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_22),
.B1(n_16),
.B2(n_8),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_225),
.B1(n_16),
.B2(n_229),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_233),
.A3(n_234),
.B1(n_235),
.B2(n_232),
.C1(n_239),
.C2(n_25),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_3),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_9),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_36),
.C(n_8),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_3),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_4),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_241),
.B(n_248),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_4),
.B(n_5),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_253),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_249),
.B(n_6),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_5),
.B(n_6),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_258),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_261),
.A2(n_7),
.B(n_36),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_262),
.A2(n_7),
.B(n_36),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_263),
.B(n_36),
.Y(n_264)
);


endmodule