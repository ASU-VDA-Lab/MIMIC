module fake_netlist_6_4211_n_166 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_166);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_166;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_28;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_160;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_130;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_66;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_29;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_126;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_3),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_63),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_69),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_43),
.B1(n_37),
.B2(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_45),
.Y(n_89)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_72),
.B(n_54),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_80),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_70),
.B(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_71),
.B(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_78),
.B(n_83),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_71),
.C(n_72),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_82),
.B(n_64),
.C(n_41),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_73),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_84),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_81),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_100),
.B(n_97),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_73),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_41),
.B(n_46),
.C(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_98),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_107),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_108),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_113),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_116),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_113),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_117),
.A2(n_112),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_92),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_102),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_102),
.B(n_108),
.Y(n_132)
);

AOI222xp33_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_65),
.B1(n_46),
.B2(n_38),
.C1(n_34),
.C2(n_68),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_98),
.Y(n_134)
);

AOI211xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_92),
.B(n_77),
.C(n_85),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_97),
.B1(n_74),
.B2(n_76),
.Y(n_136)
);

OAI211xp5_ASAP7_75t_SL g137 ( 
.A1(n_133),
.A2(n_132),
.B(n_131),
.C(n_136),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_125),
.Y(n_138)
);

AOI221x1_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_121),
.B1(n_72),
.B2(n_66),
.C(n_62),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_85),
.B(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_121),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_135),
.A2(n_66),
.B(n_72),
.C(n_62),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_140),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_71),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

AND3x1_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_62),
.C(n_66),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_123),
.B1(n_62),
.B2(n_54),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_145),
.C(n_56),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_56),
.B1(n_54),
.B2(n_96),
.C(n_101),
.Y(n_155)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_101),
.B1(n_79),
.B2(n_86),
.C(n_110),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_153),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_151),
.B(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_R g160 ( 
.A(n_156),
.B(n_14),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI22x1_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_110),
.B1(n_79),
.B2(n_24),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_90),
.B1(n_99),
.B2(n_25),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_163),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_161),
.B1(n_158),
.B2(n_162),
.Y(n_166)
);


endmodule