module fake_netlist_6_1140_n_145 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_145);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_145;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_73;
wire n_138;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

OR2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_5),
.B(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_0),
.A2(n_24),
.B1(n_5),
.B2(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_10),
.B(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

NAND2x1p5_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx8_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVxp33_ASAP7_75t_SL g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_6),
.B(n_14),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_2),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_6),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_20),
.B(n_38),
.C(n_62),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_64),
.B(n_66),
.C(n_53),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_43),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_55),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_50),
.B1(n_60),
.B2(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_55),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_40),
.B1(n_52),
.B2(n_61),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_61),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_63),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_67),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_78),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_84),
.B(n_80),
.C(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

AO31x2_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_88),
.A3(n_92),
.B(n_93),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_75),
.B(n_85),
.C(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

OAI21x1_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_86),
.B(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_86),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_97),
.Y(n_122)
);

AO31x2_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_95),
.A3(n_103),
.B(n_108),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_102),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_108),
.Y(n_125)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_115),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_108),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_114),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_127),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_116),
.B(n_127),
.C(n_125),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_101),
.B(n_96),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_120),
.B(n_112),
.C(n_118),
.Y(n_137)
);

OAI211xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_132),
.B(n_96),
.C(n_113),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_117),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_108),
.B1(n_140),
.B2(n_141),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_144),
.Y(n_145)
);


endmodule