module fake_jpeg_30945_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_9),
.B(n_0),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_6),
.C(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_16),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_17),
.B1(n_1),
.B2(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_7),
.B1(n_8),
.B2(n_6),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_19),
.B1(n_21),
.B2(n_15),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_19),
.C(n_18),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_24),
.C(n_23),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.C(n_27),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_13),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_21),
.B1(n_17),
.B2(n_13),
.Y(n_35)
);

OAI221xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_13),
.B1(n_12),
.B2(n_16),
.C(n_14),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_35),
.C(n_14),
.Y(n_37)
);

AOI211xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_34),
.B(n_12),
.C(n_3),
.Y(n_38)
);


endmodule