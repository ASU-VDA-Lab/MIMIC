module fake_jpeg_22622_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_4),
.B(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_17),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2x1_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_19),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_22),
.CI(n_7),
.CON(n_27),
.SN(n_27)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_19),
.B1(n_11),
.B2(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_21),
.B1(n_20),
.B2(n_23),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_17),
.Y(n_28)
);

NOR2xp67_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_2),
.Y(n_32)
);

FAx1_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_0),
.CI(n_1),
.CON(n_29),
.SN(n_29)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_28),
.C(n_29),
.Y(n_34)
);

BUFx24_ASAP7_75t_SL g33 ( 
.A(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_30),
.B(n_27),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_37),
.C(n_20),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_5),
.C(n_0),
.Y(n_40)
);


endmodule