module fake_jpeg_9242_n_109 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_5),
.B(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_43),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_17),
.B1(n_21),
.B2(n_12),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_15),
.B1(n_25),
.B2(n_19),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_18),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_15),
.B(n_14),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_16),
.B1(n_18),
.B2(n_14),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_63),
.B1(n_42),
.B2(n_44),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_48),
.B(n_37),
.C(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_10),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_25),
.B(n_16),
.C(n_11),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_37),
.C(n_42),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_58),
.C(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_10),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_54),
.B1(n_62),
.B2(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_69),
.B1(n_64),
.B2(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_54),
.B(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_88),
.Y(n_95)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

AO221x1_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_60),
.B1(n_65),
.B2(n_50),
.C(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_79),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_89),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_82),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_78),
.C(n_81),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.C(n_90),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_72),
.C(n_75),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_101),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_71),
.B1(n_91),
.B2(n_87),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_88),
.B(n_83),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_68),
.B(n_85),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.B1(n_103),
.B2(n_52),
.C(n_89),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_70),
.C(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_52),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_50),
.Y(n_109)
);


endmodule