module real_jpeg_14228_n_17 (n_5, n_4, n_8, n_0, n_12, n_272, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_272;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_3),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_3),
.B(n_45),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_33),
.B(n_34),
.C(n_198),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_134),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_3),
.B(n_61),
.C(n_75),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_3),
.B(n_35),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_3),
.A2(n_64),
.B(n_223),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_3),
.A2(n_31),
.B1(n_34),
.B2(n_134),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_6),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_6),
.A2(n_31),
.B1(n_34),
.B2(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_98),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_6),
.A2(n_61),
.B1(n_63),
.B2(n_98),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_31),
.B1(n_34),
.B2(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_55),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_7),
.A2(n_55),
.B1(n_61),
.B2(n_63),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_61),
.B1(n_63),
.B2(n_79),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_31),
.B1(n_34),
.B2(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_42),
.B1(n_61),
.B2(n_63),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_12),
.A2(n_31),
.B1(n_34),
.B2(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_12),
.B(n_31),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_61),
.B1(n_63),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_68),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_31),
.B1(n_34),
.B2(n_47),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_14),
.A2(n_47),
.B1(n_61),
.B2(n_63),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_16),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_16),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_16),
.A2(n_39),
.B1(n_61),
.B2(n_63),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_21),
.B(n_102),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.C(n_90),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_22),
.A2(n_23),
.B1(n_82),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_56),
.B2(n_81),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_43),
.C(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_27),
.A2(n_40),
.B1(n_41),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_27),
.A2(n_40),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_27),
.A2(n_140),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_27),
.A2(n_171),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_30),
.A2(n_36),
.B(n_134),
.Y(n_198)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_34),
.A2(n_46),
.A3(n_50),
.B1(n_136),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_35),
.B(n_101),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_37),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_37),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_38),
.A2(n_40),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_40),
.A2(n_100),
.B(n_139),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_52),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_46),
.A2(n_48),
.B(n_134),
.C(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_49),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_49),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_49),
.A2(n_97),
.B(n_119),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_53),
.B(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_70),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_57),
.A2(n_70),
.B1(n_71),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_57),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_63),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_64),
.A2(n_69),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_64),
.A2(n_69),
.B1(n_152),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_64),
.A2(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_66),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_65),
.B(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_65),
.A2(n_66),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_66),
.B(n_201),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_69),
.A2(n_160),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_69),
.A2(n_200),
.B(n_228),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_69),
.B(n_134),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_73),
.B1(n_80),
.B2(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_78),
.B1(n_80),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_73),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_73),
.A2(n_80),
.B1(n_193),
.B2(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_88),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_77),
.A2(n_143),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_77),
.B(n_134),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_80),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_82),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_89),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_84),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_89),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_90),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.C(n_99),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_91),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_94),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_95),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_96),
.B(n_99),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_124),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_112),
.B2(n_113),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_111),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_109),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_107),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_107),
.A2(n_194),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_123),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_265),
.B(n_270),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_175),
.A3(n_184),
.B1(n_263),
.B2(n_264),
.C(n_272),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_161),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_129),
.B(n_161),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_146),
.C(n_154),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_145),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_138),
.C(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_154),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_165),
.C(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_173),
.C(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_177),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_204),
.B(n_262),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_202),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_186),
.B(n_202),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_195),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_187),
.A2(n_188),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_191),
.A2(n_195),
.B1(n_196),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_197),
.B(n_199),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_255),
.B(n_261),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_243),
.B(n_254),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_224),
.B(n_242),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_208),
.B(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_241),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_230),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_236),
.B(n_240),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_234),
.B(n_235),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_245),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_250),
.C(n_253),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_269),
.Y(n_270)
);


endmodule