module fake_jpeg_17253_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_70),
.Y(n_85)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_70),
.B1(n_45),
.B2(n_71),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_86),
.B1(n_89),
.B2(n_49),
.Y(n_99)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_60),
.B1(n_52),
.B2(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_63),
.B1(n_50),
.B2(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_46),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_48),
.C(n_44),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_98),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_0),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_96),
.B(n_103),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_114),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_115),
.B(n_55),
.C(n_4),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_65),
.B1(n_56),
.B2(n_53),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_1),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_113),
.Y(n_126)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_64),
.B1(n_61),
.B2(n_58),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_2),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_54),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_55),
.B1(n_57),
.B2(n_5),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_98),
.B1(n_106),
.B2(n_101),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_106),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_135),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_96),
.B1(n_121),
.B2(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_116),
.B1(n_118),
.B2(n_100),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_116),
.CI(n_104),
.CON(n_136),
.SN(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_118),
.B1(n_127),
.B2(n_131),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_136),
.C(n_134),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_138),
.B(n_137),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_147),
.B1(n_129),
.B2(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_145),
.C(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_128),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_154),
.C(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_21),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_156),
.C(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_111),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_18),
.B(n_41),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_17),
.B(n_40),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_16),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_19),
.B(n_38),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_14),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_13),
.C(n_37),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_22),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_11),
.B1(n_33),
.B2(n_32),
.Y(n_169)
);


endmodule