module fake_jpeg_945_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_55),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_60),
.B1(n_53),
.B2(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_51),
.B1(n_44),
.B2(n_43),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_50),
.B1(n_47),
.B2(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_57),
.B1(n_46),
.B2(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_42),
.B1(n_51),
.B2(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_65),
.B1(n_52),
.B2(n_43),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_98),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_92),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_58),
.B(n_46),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_49),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_41),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_1),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_50),
.B(n_3),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_18),
.C(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_19),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_116),
.C(n_88),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_77),
.B1(n_73),
.B2(n_4),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_12),
.B(n_13),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_6),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_9),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_9),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_14),
.A3(n_15),
.B1(n_22),
.B2(n_24),
.C1(n_27),
.C2(n_28),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_10),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_109),
.B(n_101),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_120),
.B(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_88),
.B(n_94),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_93),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_10),
.B(n_11),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_32),
.B(n_33),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_112),
.B1(n_35),
.B2(n_37),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_121),
.C(n_128),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_127),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_132),
.C(n_133),
.Y(n_141)
);

NAND4xp25_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_139),
.C(n_134),
.D(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_104),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_34),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_125),
.Y(n_147)
);


endmodule