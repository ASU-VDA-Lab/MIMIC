module fake_jpeg_31079_n_492 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_492);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_492;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_50),
.Y(n_148)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_17),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_7),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_71),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_7),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_67),
.Y(n_112)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_8),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_72),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_6),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_79),
.Y(n_114)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_84),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_4),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_95),
.Y(n_116)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_16),
.Y(n_96)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_42),
.B1(n_47),
.B2(n_25),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_100),
.A2(n_127),
.B1(n_39),
.B2(n_24),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_70),
.B1(n_85),
.B2(n_54),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_113),
.A2(n_119),
.B1(n_140),
.B2(n_64),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_47),
.B1(n_25),
.B2(n_42),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_61),
.A2(n_47),
.B1(n_25),
.B2(n_45),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_134),
.B1(n_136),
.B2(n_27),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_95),
.B1(n_89),
.B2(n_73),
.Y(n_127)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_37),
.B1(n_46),
.B2(n_30),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_92),
.A2(n_48),
.B1(n_36),
.B2(n_45),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g201 ( 
.A(n_137),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_82),
.A2(n_48),
.B1(n_44),
.B2(n_36),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_74),
.Y(n_159)
);

OR2x2_ASAP7_75t_SL g152 ( 
.A(n_56),
.B(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_152),
.B(n_24),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_77),
.A2(n_43),
.B1(n_27),
.B2(n_20),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_119),
.B1(n_134),
.B2(n_131),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_97),
.B1(n_86),
.B2(n_63),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_154),
.A2(n_157),
.B1(n_171),
.B2(n_181),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_98),
.B(n_79),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_156),
.B(n_160),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_91),
.B1(n_65),
.B2(n_60),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_159),
.B(n_164),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_44),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_51),
.A3(n_52),
.B1(n_81),
.B2(n_43),
.Y(n_164)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_177),
.B1(n_203),
.B2(n_123),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_46),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_167),
.B(n_170),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_51),
.C(n_66),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_169),
.B(n_191),
.C(n_199),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_66),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_100),
.A2(n_75),
.B1(n_50),
.B2(n_78),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_172),
.A2(n_149),
.B(n_122),
.C(n_2),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_74),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_176),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_112),
.B(n_39),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_102),
.A2(n_39),
.B1(n_24),
.B2(n_41),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_14),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_106),
.B(n_24),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_114),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_190),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_39),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_108),
.B(n_0),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_1),
.Y(n_247)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_109),
.B(n_16),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_12),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_198),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_139),
.B(n_2),
.C(n_3),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_132),
.B1(n_130),
.B2(n_122),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_0),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_0),
.B(n_1),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_126),
.A2(n_125),
.B1(n_144),
.B2(n_128),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_113),
.B1(n_127),
.B2(n_126),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_218),
.B1(n_220),
.B2(n_238),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_149),
.B(n_124),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_209),
.A2(n_226),
.B(n_228),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_210),
.A2(n_183),
.B1(n_185),
.B2(n_189),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_103),
.B(n_147),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_213),
.A2(n_201),
.B1(n_163),
.B2(n_195),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_216),
.B(n_229),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_166),
.A2(n_120),
.B1(n_103),
.B2(n_105),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_171),
.A2(n_105),
.B1(n_13),
.B2(n_2),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_3),
.B1(n_14),
.B2(n_15),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_178),
.A2(n_3),
.B1(n_15),
.B2(n_1),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_1),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_242),
.C(n_193),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_1),
.B1(n_15),
.B2(n_169),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_164),
.B(n_15),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_198),
.A2(n_155),
.B1(n_191),
.B2(n_157),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_238),
.B1(n_206),
.B2(n_220),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_253),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_158),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_258),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_256),
.B(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_202),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_259),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_261),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_202),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_161),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_262),
.B(n_267),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_162),
.B1(n_200),
.B2(n_173),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_265),
.B1(n_287),
.B2(n_239),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_188),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_223),
.C(n_229),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_245),
.A2(n_231),
.B1(n_213),
.B2(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_192),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_173),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_270),
.Y(n_325)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_179),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_225),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_271),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_175),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_272),
.B(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_201),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_225),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_274),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_181),
.Y(n_275)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_216),
.B(n_183),
.Y(n_277)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_214),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_278),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_219),
.B(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_223),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_248),
.B(n_204),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_236),
.B(n_204),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_285),
.A2(n_211),
.B(n_222),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_230),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_213),
.B1(n_236),
.B2(n_210),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_288),
.A2(n_213),
.B1(n_235),
.B2(n_226),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_296),
.B1(n_309),
.B2(n_252),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_213),
.B(n_209),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_304),
.B(n_312),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_261),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_298),
.C(n_317),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_243),
.C(n_211),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_299),
.A2(n_316),
.B1(n_320),
.B2(n_251),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_210),
.B(n_222),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_251),
.A2(n_210),
.B1(n_228),
.B2(n_239),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_224),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_319),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_275),
.A2(n_210),
.B(n_240),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_314),
.A2(n_285),
.B(n_277),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_186),
.B1(n_183),
.B2(n_168),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_265),
.A2(n_263),
.B1(n_260),
.B2(n_257),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_240),
.C(n_234),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_250),
.B(n_201),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_295),
.C(n_297),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_252),
.A2(n_174),
.B1(n_234),
.B2(n_244),
.Y(n_320)
);

NOR2x1p5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_310),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_328),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_327),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_349),
.C(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_332),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_335),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_334),
.A2(n_342),
.B1(n_294),
.B2(n_304),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_292),
.B(n_282),
.Y(n_336)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_339),
.A2(n_307),
.B(n_269),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_340),
.A2(n_352),
.B1(n_272),
.B2(n_280),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_341),
.B(n_345),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_309),
.A2(n_249),
.B1(n_266),
.B2(n_284),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_279),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_348),
.Y(n_363)
);

NAND2x1_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_266),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_344),
.A2(n_269),
.B(n_307),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_318),
.B(n_262),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_347),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_305),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_298),
.C(n_302),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_353),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_299),
.A2(n_286),
.B1(n_258),
.B2(n_276),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_281),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_255),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_355),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_325),
.B(n_267),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_321),
.B(n_253),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_356),
.B(n_357),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_270),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_301),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_359),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_301),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_369),
.C(n_383),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_370),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_342),
.B1(n_326),
.B2(n_340),
.Y(n_365)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_327),
.A2(n_293),
.B1(n_320),
.B2(n_324),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_366),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_310),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_368),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_289),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_289),
.C(n_312),
.Y(n_369)
);

OA22x2_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_290),
.B1(n_324),
.B2(n_322),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_326),
.A2(n_313),
.B1(n_300),
.B2(n_322),
.Y(n_372)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_280),
.B(n_273),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_373),
.A2(n_378),
.B(n_384),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_353),
.B1(n_355),
.B2(n_354),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_274),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_387),
.A2(n_365),
.B1(n_383),
.B2(n_372),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_336),
.Y(n_391)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_391),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_381),
.B(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_337),
.C(n_346),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_401),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_343),
.Y(n_399)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_399),
.Y(n_424)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_400),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_337),
.C(n_339),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_338),
.B(n_357),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_402),
.A2(n_360),
.B(n_363),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_345),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_403),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_385),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_406),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_356),
.Y(n_405)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_380),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_359),
.C(n_369),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_408),
.Y(n_425)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_332),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_397),
.A2(n_378),
.B(n_362),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_413),
.A2(n_416),
.B(n_402),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_409),
.B1(n_392),
.B2(n_388),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_397),
.A2(n_373),
.B(n_370),
.Y(n_416)
);

A2O1A1O1Ixp25_ASAP7_75t_L g417 ( 
.A1(n_387),
.A2(n_374),
.B(n_360),
.C(n_363),
.D(n_358),
.Y(n_417)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_417),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_418),
.Y(n_440)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_394),
.A2(n_370),
.B(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_426),
.Y(n_442)
);

NAND3xp33_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_347),
.C(n_329),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_421),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_370),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_388),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_444),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_422),
.B(n_403),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_434),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_389),
.C(n_407),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_435),
.C(n_436),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_425),
.B(n_410),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_389),
.C(n_398),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_390),
.C(n_396),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_390),
.C(n_396),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_441),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_428),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_401),
.C(n_368),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_445),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_413),
.A2(n_428),
.B(n_411),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_367),
.Y(n_445)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g447 ( 
.A(n_445),
.B(n_418),
.CI(n_405),
.CON(n_447),
.SN(n_447)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_448),
.Y(n_463)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_442),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_412),
.B(n_426),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_459),
.Y(n_466)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_444),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_458),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_439),
.A2(n_392),
.B1(n_429),
.B2(n_420),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_457),
.B1(n_427),
.B2(n_417),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_440),
.A2(n_424),
.B1(n_423),
.B2(n_393),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_443),
.A2(n_393),
.B1(n_395),
.B2(n_412),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_435),
.C(n_433),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_462),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_453),
.B(n_436),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_465),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_457),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_399),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_469),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_408),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_447),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_SL g473 ( 
.A1(n_470),
.A2(n_447),
.B(n_455),
.C(n_459),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_437),
.C(n_351),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_271),
.Y(n_479)
);

AOI21xp33_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_478),
.B(n_468),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_460),
.A2(n_450),
.B(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_475),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_350),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_479),
.Y(n_483)
);

OA21x2_ASAP7_75t_SL g478 ( 
.A1(n_463),
.A2(n_406),
.B(n_400),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_477),
.C(n_464),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_481),
.A2(n_254),
.B(n_208),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_482),
.A2(n_484),
.B(n_473),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_466),
.B(n_462),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_485),
.A2(n_486),
.B(n_487),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_480),
.A2(n_254),
.B(n_208),
.Y(n_487)
);

OAI21x1_ASAP7_75t_SL g488 ( 
.A1(n_485),
.A2(n_481),
.B(n_483),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_488),
.B(n_259),
.Y(n_490)
);

OAI221xp5_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_489),
.B1(n_259),
.B2(n_232),
.C(n_180),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_491),
.B(n_232),
.Y(n_492)
);


endmodule