module fake_jpeg_17419_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_47),
.Y(n_54)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_26),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_26),
.Y(n_53)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_26),
.B1(n_16),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_64),
.B1(n_68),
.B2(n_47),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_29),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_45),
.B1(n_16),
.B2(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_22),
.B1(n_16),
.B2(n_27),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_47),
.B1(n_43),
.B2(n_39),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_22),
.B1(n_18),
.B2(n_33),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_1),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_47),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_79),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_19),
.C(n_30),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_22),
.B1(n_43),
.B2(n_39),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_83),
.A2(n_110),
.B1(n_55),
.B2(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_97),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_85),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_88),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_18),
.B(n_33),
.C(n_35),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_63),
.B(n_23),
.C(n_25),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_33),
.B1(n_18),
.B2(n_35),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_25),
.B1(n_55),
.B2(n_39),
.Y(n_123)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_95),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_53),
.B(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_30),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_64),
.B1(n_59),
.B2(n_43),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_138),
.Y(n_148)
);

OR2x4_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_20),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_137),
.B1(n_140),
.B2(n_86),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_82),
.B(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_74),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_95),
.B(n_75),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_56),
.B1(n_52),
.B2(n_68),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_135),
.B1(n_84),
.B2(n_79),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_85),
.A2(n_52),
.B1(n_73),
.B2(n_31),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_30),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_94),
.B1(n_109),
.B2(n_96),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_142),
.A2(n_146),
.B1(n_161),
.B2(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_145),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_97),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_114),
.C(n_113),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_102),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_109),
.B(n_92),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_159),
.B(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_158),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_155),
.B1(n_165),
.B2(n_168),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx2_ASAP7_75t_R g153 ( 
.A(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_109),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_106),
.B(n_87),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_78),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_99),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_167),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_123),
.B(n_121),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_105),
.B1(n_104),
.B2(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_139),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_127),
.B1(n_139),
.B2(n_28),
.Y(n_207)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_103),
.B1(n_80),
.B2(n_91),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_31),
.B1(n_28),
.B2(n_21),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_178),
.Y(n_222)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_186),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_133),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_205),
.B(n_20),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_153),
.C(n_158),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_21),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_204),
.C(n_17),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_120),
.Y(n_195)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_115),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_124),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_200),
.B(n_10),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_127),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_144),
.B(n_89),
.C(n_132),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_127),
.B(n_111),
.C(n_30),
.D(n_21),
.Y(n_205)
);

CKINVDCx12_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_161),
.B1(n_155),
.B2(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_209),
.A2(n_211),
.B1(n_213),
.B2(n_217),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_161),
.B1(n_173),
.B2(n_139),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_204),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_196),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_20),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_201),
.A2(n_20),
.B1(n_17),
.B2(n_3),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_194),
.Y(n_251)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_1),
.B(n_2),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_203),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_15),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_3),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

OAI32xp33_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_178),
.A2(n_4),
.B(n_6),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_232),
.A2(n_12),
.B(n_13),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_199),
.B1(n_178),
.B2(n_14),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_177),
.B(n_176),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_11),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_246),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_199),
.B1(n_194),
.B2(n_184),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_237),
.B1(n_228),
.B2(n_210),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_193),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_175),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_187),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_186),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_249),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_215),
.C(n_209),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_218),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_174),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_216),
.B(n_192),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_232),
.B(n_213),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_SL g261 ( 
.A(n_229),
.B(n_196),
.C(n_184),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_269),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_241),
.B1(n_248),
.B2(n_250),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_214),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_275),
.C(n_251),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_273),
.B(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_227),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_231),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_281),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_219),
.B(n_237),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_219),
.B(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_291),
.C(n_292),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_296),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_286),
.B(n_295),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_239),
.B(n_211),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_256),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_231),
.C(n_253),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_282),
.C(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_257),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_267),
.B(n_254),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_252),
.B1(n_242),
.B2(n_261),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_300),
.C(n_303),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_270),
.B(n_278),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_R g301 ( 
.A(n_284),
.B(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_270),
.C(n_280),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_285),
.B(n_266),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_268),
.B(n_274),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_293),
.B1(n_221),
.B2(n_208),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_217),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_291),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_180),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_180),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_313),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_318),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_301),
.B1(n_307),
.B2(n_221),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_208),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_303),
.B(n_275),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_300),
.B(n_179),
.Y(n_321)
);

OAI221xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_179),
.B1(n_299),
.B2(n_181),
.C(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_318),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_328),
.B1(n_329),
.B2(n_15),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_298),
.B(n_288),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_12),
.B(n_13),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_324),
.A2(n_316),
.B(n_315),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_333),
.B(n_334),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_335),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_327),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_330),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_324),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_336),
.Y(n_341)
);


endmodule