module fake_jpeg_11453_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_82),
.Y(n_91)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_59),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_51),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_70),
.B1(n_71),
.B2(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_89),
.B1(n_95),
.B2(n_98),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_71),
.B1(n_76),
.B2(n_67),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_84),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_74),
.B(n_52),
.C(n_56),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_80),
.B(n_3),
.C(n_4),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_74),
.B1(n_52),
.B2(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_100),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_63),
.B1(n_57),
.B2(n_66),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_57),
.C(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_61),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_81),
.B(n_80),
.C(n_63),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_117),
.B1(n_34),
.B2(n_45),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_113),
.Y(n_136)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_1),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_2),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_24),
.B(n_48),
.C(n_47),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_3),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_4),
.C(n_5),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_43),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_26),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_130),
.CI(n_140),
.CON(n_141),
.SN(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_9),
.C(n_10),
.Y(n_130)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_138),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_9),
.B(n_11),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_119),
.B(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_139),
.B1(n_39),
.B2(n_41),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_16),
.A3(n_17),
.B1(n_19),
.B2(n_29),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_153),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_104),
.B(n_33),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_147),
.B(n_150),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_122),
.B1(n_121),
.B2(n_138),
.Y(n_157)
);

INVxp33_ASAP7_75t_SL g147 ( 
.A(n_132),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_126),
.A3(n_136),
.B1(n_135),
.B2(n_149),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_44),
.B(n_50),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_155),
.B(n_148),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.C(n_124),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_147),
.B1(n_148),
.B2(n_128),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_164),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_163),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_142),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_160),
.B(n_157),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_165),
.B(n_164),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_127),
.B(n_141),
.C(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_141),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_158),
.Y(n_171)
);


endmodule