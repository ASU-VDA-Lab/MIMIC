module fake_jpeg_29255_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_26),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_53),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_17),
.B1(n_33),
.B2(n_31),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_23),
.B(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_37),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_46),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_67),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_66),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_16),
.B1(n_34),
.B2(n_30),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_38),
.C(n_40),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_37),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_44),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_39),
.B(n_36),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_2),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_42),
.B1(n_37),
.B2(n_12),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_11),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_2),
.CI(n_3),
.CON(n_83),
.SN(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_5),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_9),
.B1(n_10),
.B2(n_15),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_18),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_93),
.C(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_6),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_21),
.C(n_7),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_70),
.C(n_73),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_86),
.B(n_92),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_89),
.C(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_97),
.C(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_97),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_94),
.Y(n_115)
);


endmodule