module fake_jpeg_20135_n_86 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_48),
.Y(n_52)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_2),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_66),
.B1(n_18),
.B2(n_21),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_22),
.C(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_2),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_16),
.B(n_17),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_61),
.B1(n_67),
.B2(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_23),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_24),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_73),
.C(n_26),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.C(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_81),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_73),
.B1(n_27),
.B2(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_25),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_30),
.Y(n_86)
);


endmodule