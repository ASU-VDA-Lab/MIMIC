module fake_jpeg_13419_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_0),
.CON(n_51),
.SN(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_35),
.C(n_43),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_56),
.B(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_46),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_64),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_45),
.B(n_49),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_4),
.B(n_6),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_2),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_45),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_47),
.B1(n_46),
.B2(n_37),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_71),
.B(n_70),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_17),
.C(n_29),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_82),
.C(n_83),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_67),
.B1(n_16),
.B2(n_19),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_12),
.C(n_13),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_85),
.B1(n_73),
.B2(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_86),
.C(n_81),
.Y(n_90)
);

OAI21x1_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_74),
.B(n_75),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_14),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_21),
.B(n_22),
.C(n_24),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_26),
.A3(n_28),
.B1(n_30),
.B2(n_80),
.C1(n_89),
.C2(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_76),
.Y(n_96)
);


endmodule