module fake_jpeg_28273_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_25),
.Y(n_59)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_43),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_23),
.C(n_8),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_34),
.B(n_20),
.C(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_55),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_24),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_23),
.B1(n_31),
.B2(n_37),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_54),
.B1(n_57),
.B2(n_38),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_55),
.B1(n_46),
.B2(n_53),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_68),
.B1(n_78),
.B2(n_86),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_85),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_37),
.B1(n_42),
.B2(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_37),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_25),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_39),
.B1(n_17),
.B2(n_24),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_81),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_38),
.B1(n_33),
.B2(n_22),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_60),
.B1(n_20),
.B2(n_21),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_16),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_16),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_96),
.B(n_72),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_109),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_60),
.B1(n_36),
.B2(n_40),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_102),
.B1(n_112),
.B2(n_117),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_71),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_60),
.B1(n_40),
.B2(n_21),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_40),
.B1(n_41),
.B2(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_87),
.Y(n_148)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_41),
.A3(n_40),
.B1(n_18),
.B2(n_44),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_89),
.B(n_81),
.C(n_66),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_67),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_138),
.Y(n_159)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_146),
.Y(n_156)
);

NOR2x1p5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_67),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_115),
.C(n_106),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_129),
.C(n_116),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_71),
.C(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_132),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_140),
.B(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_134),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_144),
.B(n_95),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_69),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_28),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_18),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_44),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_63),
.B(n_91),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_87),
.B1(n_84),
.B2(n_63),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_119),
.B1(n_93),
.B2(n_97),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_82),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_82),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_50),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_113),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_107),
.B(n_32),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_30),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_153),
.A2(n_154),
.B(n_167),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_96),
.B(n_107),
.Y(n_154)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_120),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_161),
.B(n_165),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_117),
.B1(n_101),
.B2(n_102),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_166),
.B1(n_171),
.B2(n_2),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_116),
.B(n_113),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_129),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_138),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_50),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_97),
.B1(n_118),
.B2(n_93),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_18),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_169),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_28),
.B(n_14),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_12),
.B1(n_15),
.B2(n_13),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_143),
.B1(n_140),
.B2(n_125),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_181),
.B1(n_144),
.B2(n_132),
.Y(n_185)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_174),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_6),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_1),
.B(n_2),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_126),
.A2(n_87),
.B1(n_108),
.B2(n_27),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_149),
.B1(n_135),
.B2(n_30),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_108),
.B1(n_40),
.B2(n_27),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_189),
.B1(n_210),
.B2(n_214),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_122),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_200),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_201),
.C(n_206),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_127),
.B1(n_146),
.B2(n_136),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_212),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_177),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_184),
.Y(n_217)
);

OAI22x1_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_30),
.B1(n_22),
.B2(n_19),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_199),
.B1(n_211),
.B2(n_181),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_22),
.B1(n_19),
.B2(n_9),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_22),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_6),
.C(n_12),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_209),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_6),
.B1(n_11),
.B2(n_9),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_5),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_154),
.C(n_153),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_158),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_217),
.B(n_225),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_232),
.B(n_167),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_213),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_193),
.B1(n_176),
.B2(n_201),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_159),
.C(n_158),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_231),
.C(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_207),
.C(n_200),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_152),
.B(n_157),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_184),
.B(n_152),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_233),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_159),
.C(n_151),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_174),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_194),
.B1(n_195),
.B2(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_189),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_218),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_191),
.B1(n_206),
.B2(n_187),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_231),
.C(n_219),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_253),
.C(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_151),
.C(n_180),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_192),
.B1(n_193),
.B2(n_5),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_263),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_215),
.B1(n_222),
.B2(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_236),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_271),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_220),
.C(n_228),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_220),
.C(n_227),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_232),
.C(n_224),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_225),
.B1(n_229),
.B2(n_11),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_272),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_254),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_244),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_239),
.B1(n_243),
.B2(n_241),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_242),
.B(n_239),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_245),
.B(n_271),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_251),
.B1(n_243),
.B2(n_241),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_265),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_299),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_262),
.B(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_297),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_246),
.B(n_13),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_283),
.B(n_277),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_284),
.C(n_3),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_13),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

NAND5xp2_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_277),
.C(n_284),
.D(n_282),
.E(n_288),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_305),
.B(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_312)
);

AOI31xp67_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_3),
.A3(n_4),
.B(n_296),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_4),
.B1(n_306),
.B2(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_3),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_299),
.C(n_290),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NAND4xp25_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.C(n_313),
.D(n_309),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_315),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule