module real_jpeg_18737_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_471),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_0),
.B(n_472),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_37),
.B1(n_40),
.B2(n_47),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_47),
.B1(n_101),
.B2(n_105),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_1),
.A2(n_47),
.B1(n_180),
.B2(n_185),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_1),
.A2(n_47),
.B1(n_263),
.B2(n_266),
.Y(n_262)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_3),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_3),
.Y(n_353)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_64),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_4),
.A2(n_64),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_5),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_53),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_53),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_53),
.B1(n_204),
.B2(n_209),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_7),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_60),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_7),
.A2(n_60),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_7),
.A2(n_60),
.B1(n_289),
.B2(n_291),
.Y(n_288)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_8),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_12),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_12),
.Y(n_221)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_146),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_54),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_18),
.B(n_54),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_28),
.B1(n_36),
.B2(n_48),
.Y(n_18)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_19),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_20),
.A2(n_28),
.B1(n_57),
.B2(n_62),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_20),
.A2(n_28),
.B1(n_57),
.B2(n_62),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_20),
.B(n_28),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_28),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_21),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_22),
.Y(n_304)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_28),
.A2(n_36),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_28),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_28)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_30),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_30),
.Y(n_348)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_32),
.Y(n_308)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_33),
.Y(n_194)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_34),
.Y(n_197)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_136),
.C(n_140),
.Y(n_54)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_55),
.B(n_136),
.CI(n_140),
.CON(n_166),
.SN(n_166)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_67),
.C(n_99),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_56),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_56),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_56),
.B(n_250),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_56),
.B(n_191),
.C(n_444),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_56),
.A2(n_152),
.B1(n_191),
.B2(n_328),
.Y(n_451)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_63),
.A2(n_64),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_63),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_63),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_63),
.B(n_379),
.C(n_382),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_63),
.B(n_319),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_63),
.B(n_190),
.Y(n_396)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_64),
.B(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_64),
.Y(n_370)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2x2_ASAP7_75t_L g154 ( 
.A(n_68),
.B(n_99),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_68),
.B(n_160),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_91),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_69),
.B(n_228),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_78),
.Y(n_69)
);

NAND2x1_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g255 ( 
.A1(n_70),
.A2(n_78),
.B1(n_229),
.B2(n_256),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_75),
.Y(n_381)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_76),
.Y(n_292)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_85),
.B2(n_88),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_90),
.Y(n_234)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_90),
.Y(n_259)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_90),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_91),
.A2(n_178),
.B1(n_179),
.B2(n_190),
.Y(n_177)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_98),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_107),
.B1(n_129),
.B2(n_130),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_100),
.A2(n_107),
.B1(n_129),
.B2(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

AOI22x1_ASAP7_75t_L g250 ( 
.A1(n_107),
.A2(n_129),
.B1(n_161),
.B2(n_251),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_107),
.A2(n_129),
.B(n_161),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_120),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_128),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_129),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_138),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_143),
.B1(n_192),
.B2(n_198),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_167),
.B(n_469),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_166),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_149),
.B(n_166),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.C(n_158),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_151),
.B1(n_155),
.B2(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_152),
.B(n_249),
.C(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_159),
.C(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_155),
.A2(n_156),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_155),
.B(n_427),
.C(n_432),
.Y(n_426)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_174),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_157),
.B(n_432),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_157),
.B(n_250),
.C(n_278),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_166),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_272),
.B(n_466),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_237),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_169),
.A2(n_467),
.B(n_468),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_170),
.B(n_172),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_199),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_176),
.A2(n_177),
.B(n_191),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_178),
.A2(n_179),
.B1(n_190),
.B2(n_228),
.Y(n_227)
);

AO22x2_ASAP7_75t_L g364 ( 
.A1(n_178),
.A2(n_190),
.B1(n_228),
.B2(n_365),
.Y(n_364)
);

BUFx2_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_183),
.Y(n_231)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_191),
.B(n_283),
.C(n_285),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_191),
.A2(n_324),
.B1(n_325),
.B2(n_328),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_191),
.Y(n_328)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_200),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_225),
.B(n_235),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_202),
.B1(n_235),
.B2(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_201),
.A2(n_202),
.B1(n_227),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_212),
.Y(n_202)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_212),
.B(n_294),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_213),
.A2(n_262),
.B1(n_269),
.B2(n_270),
.Y(n_261)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_214),
.B(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_214),
.A2(n_288),
.B1(n_294),
.B2(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_216),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_221),
.Y(n_385)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_244),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_227),
.Y(n_425)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_238),
.B(n_242),
.Y(n_467)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_248),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_243),
.A2(n_246),
.B1(n_247),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_243),
.Y(n_419)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_248),
.B(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_250),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_249),
.A2(n_250),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_R g408 ( 
.A(n_249),
.B(n_364),
.C(n_366),
.Y(n_408)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_253),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_254),
.A2(n_255),
.B1(n_368),
.B2(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_254),
.A2(n_255),
.B1(n_329),
.B2(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_254),
.A2(n_255),
.B1(n_261),
.B2(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_255),
.B(n_322),
.C(n_329),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_255),
.B(n_316),
.C(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_256),
.Y(n_365)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_261),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_262),
.A2(n_293),
.B(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_267),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_268),
.Y(n_394)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AO221x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_415),
.B1(n_459),
.B2(n_464),
.C(n_465),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_358),
.B(n_414),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_321),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_275),
.B(n_321),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_276),
.B(n_282),
.C(n_299),
.Y(n_456)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_299),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_285),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_285),
.B(n_389),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B(n_293),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_315),
.B2(n_316),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_301),
.B(n_315),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_305),
.B1(n_310),
.B2(n_314),
.Y(n_301)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_315),
.A2(n_316),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_396),
.Y(n_397)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_322),
.A2(n_323),
.B1(n_410),
.B2(n_412),
.Y(n_409)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_327),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_357),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_330),
.B(n_357),
.Y(n_366)
);

OAI32xp33_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_333),
.A3(n_336),
.B1(n_342),
.B2(n_349),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_407),
.B(n_413),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_371),
.B(n_406),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_367),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_367),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_366),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_363),
.A2(n_364),
.B1(n_375),
.B2(n_386),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_363),
.A2(n_364),
.B1(n_428),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_386),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_364),
.B(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

AOI21x1_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_399),
.B(n_405),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_387),
.B(n_398),
.Y(n_372)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_395),
.B(n_397),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_SL g405 ( 
.A(n_400),
.B(n_401),
.Y(n_405)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_409),
.Y(n_413)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_410),
.Y(n_412)
);

NOR3xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_433),
.C(n_445),
.Y(n_415)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_416),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_420),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_420),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.C(n_426),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_422),
.B1(n_424),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_435),
.Y(n_434)
);

XNOR2x1_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_433),
.A2(n_460),
.B(n_461),
.C(n_463),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_437),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.C(n_442),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_440),
.Y(n_448)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_444),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_455),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_449),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_454),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_458),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_454),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_457),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);


endmodule