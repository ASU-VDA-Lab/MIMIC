module fake_ariane_503_n_1005 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1005);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1005;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_516;
wire n_307;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_906;
wire n_690;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_953;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_770;
wire n_928;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_429;
wire n_365;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_861;
wire n_780;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_658;
wire n_705;
wire n_630;
wire n_617;
wire n_570;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_527;
wire n_290;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_967;
wire n_999;
wire n_998;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_548;
wire n_289;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

BUFx10_ASAP7_75t_L g195 ( 
.A(n_3),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_95),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_91),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_43),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_84),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_189),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_142),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_34),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_62),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_72),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_140),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_69),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_115),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_181),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g227 ( 
.A(n_105),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_111),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_188),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_124),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_112),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_161),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_61),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_108),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_48),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_113),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_100),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_10),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_136),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_98),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_190),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_16),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_23),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_169),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_52),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_102),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_153),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_128),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_81),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_0),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_90),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_180),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_94),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_127),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_155),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_55),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_13),
.Y(n_269)
);

BUFx2_ASAP7_75t_R g270 ( 
.A(n_8),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_18),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_0),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_184),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

BUFx2_ASAP7_75t_SL g278 ( 
.A(n_41),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_179),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_5),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_58),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_50),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_70),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_86),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_165),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_75),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_156),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_160),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_154),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_167),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_150),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_76),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_74),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_141),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_3),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_9),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_79),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_60),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_175),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_12),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_109),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_214),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_195),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_266),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_211),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_205),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_195),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_225),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_233),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_218),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_219),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_220),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_224),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_238),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_250),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_203),
.Y(n_339)
);

INVxp33_ASAP7_75t_SL g340 ( 
.A(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_252),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_273),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_275),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_277),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_296),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_294),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_264),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_265),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_284),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_297),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_198),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_196),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_212),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_209),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_280),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_199),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_200),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_278),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_201),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_202),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_204),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_197),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_206),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_207),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_197),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_270),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_208),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_210),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_213),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_215),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_216),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_197),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_217),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_221),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_222),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_197),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_223),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_292),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_226),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_229),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_377),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_230),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_372),
.A2(n_232),
.B(n_231),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_235),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_227),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_326),
.A2(n_311),
.B1(n_308),
.B2(n_237),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_332),
.B(n_246),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_239),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_387),
.Y(n_405)
);

AND2x6_ASAP7_75t_L g406 ( 
.A(n_364),
.B(n_246),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_240),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_345),
.A2(n_274),
.B1(n_306),
.B2(n_244),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_333),
.B(n_246),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_246),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_331),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_363),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_316),
.B(n_241),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_339),
.B(n_245),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_338),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_247),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_317),
.B(n_249),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_314),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_343),
.B(n_283),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_347),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_351),
.B(n_283),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_362),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_353),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_356),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_329),
.Y(n_450)
);

AND2x2_ASAP7_75t_SL g451 ( 
.A(n_319),
.B(n_283),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_451),
.B(n_373),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_426),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_438),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_329),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_320),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_450),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_450),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_393),
.B(n_360),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_420),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_414),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_R g465 ( 
.A(n_425),
.B(n_388),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_342),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_444),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_R g468 ( 
.A(n_427),
.B(n_388),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_392),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_392),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_409),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_409),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_393),
.B(n_366),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_R g476 ( 
.A(n_429),
.B(n_344),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_397),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_416),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_439),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_439),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_373),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_398),
.B(n_369),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_441),
.B(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_441),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_401),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_426),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_426),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_426),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_446),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_446),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_446),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_434),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_328),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_446),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_398),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_R g501 ( 
.A(n_435),
.B(n_371),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_412),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_412),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_432),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_R g506 ( 
.A(n_442),
.B(n_383),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_443),
.B(n_385),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_436),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_395),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_404),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_418),
.B(n_362),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_403),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_400),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_448),
.B(n_346),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_400),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_402),
.B(n_355),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_418),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_407),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_R g520 ( 
.A(n_423),
.B(n_348),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_407),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_418),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_407),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_407),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_480),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

INVx4_ASAP7_75t_SL g527 ( 
.A(n_496),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_454),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_482),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_403),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_482),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_464),
.A2(n_396),
.B1(n_348),
.B2(n_422),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_498),
.B(n_503),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_509),
.B(n_510),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_504),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_496),
.B(n_424),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_455),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_500),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_463),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_505),
.A2(n_340),
.B1(n_447),
.B2(n_433),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_494),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_466),
.B(n_327),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_459),
.B(n_365),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_457),
.B(n_376),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_462),
.B(n_340),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_493),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_460),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_515),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_493),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_467),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_452),
.B(n_449),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_496),
.B(n_449),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_489),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_461),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_518),
.B(n_402),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_491),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_471),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_473),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_514),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_478),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

AND2x4_ASAP7_75t_SL g570 ( 
.A(n_499),
.B(n_325),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_483),
.B(n_440),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_469),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_475),
.B(n_440),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_511),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_492),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_472),
.B(n_430),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_497),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_513),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_519),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_474),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_479),
.B(n_430),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_508),
.A2(n_447),
.B1(n_433),
.B2(n_431),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_522),
.B(n_365),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_495),
.B(n_445),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_521),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_520),
.B(n_324),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_512),
.A2(n_488),
.B1(n_477),
.B2(n_396),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_520),
.B(n_325),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_481),
.B(n_431),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_445),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_517),
.B(n_402),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_484),
.B(n_419),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_468),
.B(n_501),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_523),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_524),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_527),
.B(n_506),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_525),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_573),
.B(n_408),
.Y(n_602)
);

OR2x6_ASAP7_75t_SL g603 ( 
.A(n_551),
.B(n_507),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_555),
.Y(n_604)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_527),
.B(n_421),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_528),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_534),
.B(n_476),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_561),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_531),
.B(n_422),
.Y(n_612)
);

AND3x4_ASAP7_75t_L g613 ( 
.A(n_575),
.B(n_408),
.C(n_1),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_565),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_564),
.B(n_413),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_526),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_531),
.B(n_422),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_526),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_529),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_571),
.A2(n_413),
.B1(n_359),
.B2(n_358),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_545),
.B(n_413),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_588),
.B(n_357),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_539),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_549),
.A2(n_251),
.B1(n_258),
.B2(n_254),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_565),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_566),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_541),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_540),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_566),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_540),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_544),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_568),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_570),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_536),
.B(n_530),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_591),
.A2(n_396),
.B1(n_406),
.B2(n_422),
.Y(n_639)
);

AND2x4_ASAP7_75t_L g640 ( 
.A(n_564),
.B(n_406),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_537),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_562),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_544),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_592),
.B(n_1),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_538),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_574),
.A2(n_406),
.B1(n_415),
.B2(n_307),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_557),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_596),
.B(n_415),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_564),
.B(n_406),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_283),
.Y(n_652)
);

NOR2x1p5_ASAP7_75t_L g653 ( 
.A(n_548),
.B(n_256),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_558),
.B(n_305),
.Y(n_654)
);

OAI221xp5_ASAP7_75t_L g655 ( 
.A1(n_589),
.A2(n_542),
.B1(n_584),
.B2(n_574),
.C(n_594),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_552),
.B(n_406),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_552),
.B(n_257),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_587),
.B(n_2),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_554),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_623),
.B(n_587),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_610),
.B(n_576),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_638),
.B(n_597),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_642),
.Y(n_663)
);

NOR2xp67_ASAP7_75t_L g664 ( 
.A(n_604),
.B(n_567),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_SL g665 ( 
.A1(n_654),
.A2(n_582),
.B(n_597),
.C(n_572),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_602),
.A2(n_638),
.B(n_641),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_621),
.B(n_579),
.Y(n_667)
);

NOR2x1_ASAP7_75t_L g668 ( 
.A(n_624),
.B(n_558),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_645),
.A2(n_586),
.B(n_598),
.C(n_580),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_629),
.B(n_576),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_602),
.A2(n_546),
.B(n_550),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_609),
.B(n_579),
.Y(n_672)
);

CKINVDCx6p67_ASAP7_75t_R g673 ( 
.A(n_603),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_605),
.A2(n_585),
.B1(n_590),
.B2(n_533),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_654),
.A2(n_550),
.B(n_546),
.C(n_560),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_611),
.B(n_614),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_625),
.A2(n_577),
.B1(n_583),
.B2(n_539),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g678 ( 
.A1(n_656),
.A2(n_593),
.B(n_535),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_643),
.A2(n_599),
.B(n_553),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_627),
.B(n_577),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_604),
.B(n_576),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_657),
.A2(n_553),
.B(n_560),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_608),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_628),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_655),
.B(n_595),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_645),
.A2(n_563),
.B(n_583),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_615),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_631),
.B(n_646),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_608),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_657),
.A2(n_553),
.B(n_578),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_620),
.A2(n_578),
.B(n_556),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_647),
.B(n_581),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_608),
.Y(n_693)
);

BUFx12f_ASAP7_75t_L g694 ( 
.A(n_636),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_615),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_606),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_655),
.B(n_556),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_633),
.A2(n_543),
.B1(n_528),
.B2(n_307),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_635),
.B(n_528),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_640),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_620),
.A2(n_543),
.B(n_262),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_637),
.B(n_543),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_626),
.B(n_4),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_601),
.A2(n_616),
.B(n_607),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_658),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_650),
.B(n_7),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_618),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_658),
.A2(n_634),
.B1(n_632),
.B2(n_644),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_619),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_626),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_630),
.A2(n_289),
.B(n_263),
.C(n_303),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_660),
.B(n_649),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_663),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_SL g714 ( 
.A(n_705),
.B(n_600),
.C(n_613),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_662),
.B(n_649),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_685),
.A2(n_600),
.B1(n_653),
.B2(n_612),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_SL g717 ( 
.A(n_661),
.B(n_267),
.C(n_260),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_676),
.B(n_606),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_703),
.B(n_640),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_680),
.B(n_697),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_710),
.B(n_651),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_669),
.A2(n_652),
.B(n_612),
.C(n_617),
.Y(n_722)
);

BUFx4f_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_694),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_667),
.B(n_651),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_666),
.A2(n_656),
.B(n_639),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_691),
.A2(n_648),
.B(n_659),
.C(n_622),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_670),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_686),
.B(n_652),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_671),
.A2(n_617),
.B(n_648),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_SL g731 ( 
.A(n_700),
.B(n_268),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_696),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_677),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_689),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_684),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_707),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_708),
.B(n_291),
.C(n_281),
.Y(n_737)
);

O2A1O1Ixp5_ASAP7_75t_L g738 ( 
.A1(n_675),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_738)
);

O2A1O1Ixp5_ASAP7_75t_SL g739 ( 
.A1(n_681),
.A2(n_307),
.B(n_305),
.C(n_300),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_687),
.B(n_276),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_689),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_695),
.A2(n_295),
.B1(n_285),
.B2(n_299),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_696),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_696),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_672),
.B(n_282),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_683),
.B(n_693),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_700),
.B(n_21),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_706),
.A2(n_298),
.B1(n_290),
.B2(n_307),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_692),
.B(n_683),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_682),
.A2(n_305),
.B(n_103),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_683),
.B(n_11),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_674),
.A2(n_709),
.B1(n_688),
.B2(n_699),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_702),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_693),
.B(n_12),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_678),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_665),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_700),
.B(n_15),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_723),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_713),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_732),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_736),
.Y(n_761)
);

INVx5_ASAP7_75t_SL g762 ( 
.A(n_713),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_741),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_734),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_734),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_735),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_740),
.Y(n_767)
);

INVx6_ASAP7_75t_SL g768 ( 
.A(n_747),
.Y(n_768)
);

INVx5_ASAP7_75t_L g769 ( 
.A(n_732),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_747),
.B(n_693),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_753),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_755),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_746),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_712),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_732),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_715),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_743),
.Y(n_777)
);

BUFx2_ASAP7_75t_SL g778 ( 
.A(n_724),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_729),
.B(n_668),
.Y(n_779)
);

BUFx2_ASAP7_75t_SL g780 ( 
.A(n_743),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_744),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_720),
.B(n_704),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_721),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_716),
.B(n_690),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_719),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_718),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_725),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_726),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_749),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_728),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_733),
.A2(n_752),
.B1(n_745),
.B2(n_748),
.Y(n_792)
);

BUFx12f_ASAP7_75t_L g793 ( 
.A(n_751),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_714),
.Y(n_794)
);

BUFx4f_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

CKINVDCx6p67_ASAP7_75t_R g796 ( 
.A(n_757),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_754),
.Y(n_797)
);

INVx5_ASAP7_75t_L g798 ( 
.A(n_722),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_727),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_737),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_738),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_742),
.B(n_664),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_750),
.Y(n_803)
);

BUFx12f_ASAP7_75t_L g804 ( 
.A(n_756),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_730),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_739),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_712),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_732),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_755),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_791),
.B(n_679),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_807),
.B(n_18),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_794),
.B(n_19),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_773),
.B(n_701),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_766),
.Y(n_814)
);

AO21x2_ASAP7_75t_L g815 ( 
.A1(n_806),
.A2(n_711),
.B(n_698),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_790),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_784),
.A2(n_305),
.B(n_22),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_761),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_771),
.Y(n_819)
);

OA21x2_ASAP7_75t_L g820 ( 
.A1(n_788),
.A2(n_19),
.B(n_193),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_789),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_788),
.A2(n_24),
.B(n_25),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_782),
.A2(n_27),
.B(n_28),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_798),
.A2(n_29),
.B(n_30),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_792),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_776),
.B(n_36),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_804),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_827)
);

AO21x2_ASAP7_75t_L g828 ( 
.A1(n_782),
.A2(n_40),
.B(n_42),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_802),
.A2(n_795),
.B(n_798),
.C(n_800),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_L g830 ( 
.A(n_791),
.B(n_44),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_787),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_760),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_758),
.B(n_45),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_795),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_834)
);

OA21x2_ASAP7_75t_L g835 ( 
.A1(n_799),
.A2(n_192),
.B(n_54),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_798),
.A2(n_51),
.B(n_56),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_57),
.Y(n_837)
);

AOI21xp33_ASAP7_75t_L g838 ( 
.A1(n_801),
.A2(n_59),
.B(n_63),
.Y(n_838)
);

OAI21x1_ASAP7_75t_L g839 ( 
.A1(n_805),
.A2(n_64),
.B(n_65),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_772),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_774),
.B(n_66),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_772),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_803),
.A2(n_67),
.B(n_68),
.C(n_71),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_769),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_796),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_845)
);

AOI21xp33_ASAP7_75t_L g846 ( 
.A1(n_786),
.A2(n_82),
.B(n_83),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_785),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_783),
.B(n_85),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_809),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_779),
.A2(n_87),
.B(n_89),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_825),
.A2(n_800),
.B1(n_793),
.B2(n_787),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_814),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_821),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_827),
.A2(n_797),
.B1(n_800),
.B2(n_768),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_815),
.A2(n_787),
.B1(n_786),
.B2(n_783),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_832),
.Y(n_856)
);

BUFx2_ASAP7_75t_SL g857 ( 
.A(n_844),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_814),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_847),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_818),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_820),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_819),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_840),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_840),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_842),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_811),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_844),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_842),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_849),
.Y(n_869)
);

AO21x1_ASAP7_75t_SL g870 ( 
.A1(n_849),
.A2(n_768),
.B(n_779),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_843),
.A2(n_770),
.B(n_763),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_831),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_810),
.A2(n_775),
.B(n_777),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_816),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_848),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_820),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_832),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_828),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_837),
.Y(n_879)
);

AO31x2_ASAP7_75t_L g880 ( 
.A1(n_876),
.A2(n_829),
.A3(n_836),
.B(n_824),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_866),
.A2(n_812),
.B1(n_835),
.B2(n_813),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_853),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_853),
.B(n_758),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_859),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_R g885 ( 
.A(n_856),
.B(n_767),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_859),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_SL g887 ( 
.A(n_867),
.B(n_781),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_856),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_858),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_R g890 ( 
.A(n_861),
.B(n_835),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_877),
.B(n_813),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_858),
.B(n_809),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_879),
.B(n_826),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_877),
.B(n_762),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_862),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_874),
.B(n_762),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_851),
.A2(n_834),
.B1(n_845),
.B2(n_830),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_875),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_889),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_892),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_898),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_886),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_893),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_895),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_884),
.B(n_852),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_888),
.B(n_863),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_891),
.B(n_868),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_891),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_882),
.B(n_869),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_894),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_880),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_911),
.A2(n_881),
.B(n_897),
.C(n_883),
.Y(n_912)
);

AOI21xp33_ASAP7_75t_L g913 ( 
.A1(n_911),
.A2(n_890),
.B(n_881),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_904),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_908),
.A2(n_861),
.B(n_873),
.Y(n_915)
);

NAND4xp25_ASAP7_75t_L g916 ( 
.A(n_909),
.B(n_883),
.C(n_887),
.D(n_896),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_902),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_L g918 ( 
.A1(n_912),
.A2(n_902),
.B1(n_910),
.B2(n_908),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_917),
.B(n_910),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_916),
.Y(n_920)
);

OAI221xp5_ASAP7_75t_L g921 ( 
.A1(n_913),
.A2(n_903),
.B1(n_890),
.B2(n_900),
.C(n_871),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_914),
.B(n_901),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_919),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_920),
.B(n_906),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_922),
.B(n_907),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_918),
.B(n_905),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_921),
.B(n_905),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_923),
.B(n_899),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_923),
.B(n_915),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_925),
.B(n_885),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_928),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_929),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_930),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_929),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_933),
.B(n_924),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_931),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_934),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_932),
.B(n_927),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_934),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_933),
.B(n_924),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_933),
.Y(n_941)
);

OAI211xp5_ASAP7_75t_SL g942 ( 
.A1(n_935),
.A2(n_926),
.B(n_885),
.C(n_854),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_939),
.Y(n_943)
);

OR4x1_ASAP7_75t_L g944 ( 
.A(n_937),
.B(n_936),
.C(n_940),
.D(n_941),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_938),
.A2(n_759),
.B1(n_778),
.B2(n_861),
.Y(n_945)
);

AOI21xp33_ASAP7_75t_L g946 ( 
.A1(n_941),
.A2(n_878),
.B(n_841),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_941),
.B(n_764),
.Y(n_947)
);

AOI21xp33_ASAP7_75t_SL g948 ( 
.A1(n_935),
.A2(n_765),
.B(n_770),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_939),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_941),
.B(n_904),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_943),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_949),
.B(n_864),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_947),
.B(n_864),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_945),
.B(n_867),
.Y(n_954)
);

NOR2x1_ASAP7_75t_L g955 ( 
.A(n_942),
.B(n_833),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_950),
.B(n_867),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_944),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_957),
.B(n_951),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_956),
.B(n_948),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_952),
.B(n_946),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_954),
.B(n_955),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_953),
.B(n_865),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_951),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_951),
.Y(n_965)
);

AOI211x1_ASAP7_75t_L g966 ( 
.A1(n_959),
.A2(n_873),
.B(n_846),
.C(n_838),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_958),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_964),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_961),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_963),
.A2(n_878),
.B1(n_855),
.B2(n_780),
.Y(n_970)
);

OAI211xp5_ASAP7_75t_L g971 ( 
.A1(n_965),
.A2(n_781),
.B(n_822),
.C(n_839),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_960),
.B(n_850),
.C(n_823),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_962),
.B(n_865),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_SL g974 ( 
.A(n_967),
.B(n_857),
.C(n_93),
.Y(n_974)
);

AOI221xp5_ASAP7_75t_L g975 ( 
.A1(n_968),
.A2(n_872),
.B1(n_760),
.B2(n_808),
.C(n_862),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_969),
.A2(n_817),
.B(n_872),
.C(n_880),
.Y(n_976)
);

NAND4xp25_ASAP7_75t_L g977 ( 
.A(n_966),
.B(n_857),
.C(n_870),
.D(n_769),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_L g978 ( 
.A(n_971),
.B(n_92),
.C(n_96),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_978),
.A2(n_974),
.B1(n_976),
.B2(n_975),
.C(n_973),
.Y(n_979)
);

OAI21xp33_ASAP7_75t_SL g980 ( 
.A1(n_977),
.A2(n_970),
.B(n_972),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_974),
.A2(n_769),
.B1(n_808),
.B2(n_760),
.Y(n_981)
);

OAI221xp5_ASAP7_75t_SL g982 ( 
.A1(n_978),
.A2(n_870),
.B1(n_880),
.B2(n_860),
.C(n_808),
.Y(n_982)
);

OAI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_982),
.A2(n_860),
.B1(n_880),
.B2(n_104),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_979),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_984),
.B(n_980),
.Y(n_985)
);

NAND5xp2_ASAP7_75t_L g986 ( 
.A(n_983),
.B(n_981),
.C(n_101),
.D(n_106),
.E(n_110),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_985),
.Y(n_987)
);

NOR2xp67_ASAP7_75t_L g988 ( 
.A(n_986),
.B(n_99),
.Y(n_988)
);

AND4x1_ASAP7_75t_L g989 ( 
.A(n_987),
.B(n_114),
.C(n_116),
.D(n_117),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_988),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_990),
.Y(n_991)
);

NAND4xp25_ASAP7_75t_L g992 ( 
.A(n_989),
.B(n_118),
.C(n_119),
.D(n_120),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_991),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_992),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_993),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_SL g996 ( 
.A1(n_994),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_993),
.B(n_129),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_995),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_997),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_999),
.A2(n_996),
.B1(n_134),
.B2(n_135),
.Y(n_1000)
);

XNOR2xp5_ASAP7_75t_L g1001 ( 
.A(n_1000),
.B(n_998),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_SL g1002 ( 
.A1(n_1001),
.A2(n_133),
.B1(n_138),
.B2(n_139),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_1002),
.B(n_143),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_1003),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_1004)
);

AOI211xp5_ASAP7_75t_L g1005 ( 
.A1(n_1004),
.A2(n_148),
.B(n_149),
.C(n_152),
.Y(n_1005)
);


endmodule