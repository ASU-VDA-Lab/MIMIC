module fake_jpeg_16115_n_159 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_159);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_1),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_50),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_33),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_37),
.Y(n_69)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_55),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_69),
.Y(n_77)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_34),
.B1(n_20),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_65),
.B1(n_32),
.B2(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_72),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_20),
.B1(n_28),
.B2(n_34),
.Y(n_65)
);

OA22x2_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_71),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_36),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_53),
.B1(n_49),
.B2(n_62),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_17),
.A3(n_14),
.B1(n_23),
.B2(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_43),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_47),
.C(n_46),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_47),
.C(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_35),
.B1(n_49),
.B2(n_23),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_72),
.B1(n_14),
.B2(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_21),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_104),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_70),
.B(n_71),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_57),
.B(n_66),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_58),
.B1(n_54),
.B2(n_53),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_100),
.B1(n_82),
.B2(n_83),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_66),
.B(n_57),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_74),
.A2(n_25),
.B1(n_24),
.B2(n_15),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_25),
.B(n_24),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_86),
.B(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_81),
.C(n_76),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_115),
.C(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_117),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_77),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_98),
.B1(n_79),
.B2(n_29),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_95),
.B(n_102),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_91),
.C(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_22),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_124),
.C(n_116),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_131),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_97),
.A3(n_98),
.B1(n_100),
.B2(n_85),
.C1(n_87),
.C2(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_130),
.B1(n_132),
.B2(n_109),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_98),
.B(n_4),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_18),
.C(n_29),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_120),
.C(n_115),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_29),
.B1(n_22),
.B2(n_18),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_136),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_140),
.C(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_146),
.Y(n_147)
);

OR2x6_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_108),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_134),
.B(n_127),
.C(n_22),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_9),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_145),
.B(n_137),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_149),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_141),
.B(n_9),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_151),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_8),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_147),
.B(n_10),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_155),
.A2(n_156),
.B(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_10),
.Y(n_156)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_11),
.A3(n_12),
.B1(n_6),
.B2(n_3),
.C(n_5),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_3),
.Y(n_159)
);


endmodule