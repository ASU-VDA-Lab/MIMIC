module real_jpeg_31725_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_0),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_91),
.B1(n_92),
.B2(n_97),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_1),
.A2(n_91),
.B1(n_302),
.B2(n_307),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_1),
.A2(n_91),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_1),
.A2(n_91),
.B1(n_444),
.B2(n_450),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_3),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_3),
.A2(n_162),
.B1(n_249),
.B2(n_252),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_3),
.A2(n_162),
.B1(n_378),
.B2(n_382),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_3),
.A2(n_162),
.B1(n_425),
.B2(n_430),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_4),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_4),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_5),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_128),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_5),
.A2(n_128),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_5),
.A2(n_128),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_6),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g341 ( 
.A(n_6),
.B(n_99),
.Y(n_341)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_6),
.A2(n_349),
.A3(n_352),
.B1(n_356),
.B2(n_362),
.Y(n_348)
);

OAI32xp33_ASAP7_75t_L g400 ( 
.A1(n_6),
.A2(n_349),
.A3(n_352),
.B1(n_356),
.B2(n_362),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_6),
.A2(n_298),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

OAI21xp33_ASAP7_75t_L g489 ( 
.A1(n_6),
.A2(n_189),
.B(n_435),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_7),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_7),
.A2(n_196),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_7),
.A2(n_196),
.B1(n_332),
.B2(n_336),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_8),
.A2(n_39),
.B1(n_229),
.B2(n_234),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_11),
.Y(n_449)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_12),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_12),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_14),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_15),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_15),
.Y(n_184)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_16),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_16),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_16),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_17),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_18),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_18),
.A2(n_55),
.B1(n_267),
.B2(n_271),
.Y(n_266)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_313),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_274),
.B(n_312),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_24),
.B(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_174),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_88),
.C(n_131),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2x1_ASAP7_75t_L g276 ( 
.A(n_28),
.B(n_277),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_62),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_29),
.B(n_62),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_37),
.B1(n_48),
.B2(n_54),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_30),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_30),
.B(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_30),
.A2(n_442),
.B1(n_453),
.B2(n_455),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_33),
.Y(n_188)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_33),
.Y(n_209)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_33),
.Y(n_335)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_34),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_36),
.Y(n_258)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_38),
.A2(n_189),
.B1(n_331),
.B2(n_337),
.Y(n_330)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_43),
.Y(n_183)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_43),
.Y(n_429)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_46),
.Y(n_336)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_48),
.B(n_372),
.Y(n_435)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_53),
.Y(n_180)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_53),
.Y(n_339)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_54),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_57),
.Y(n_374)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_60),
.Y(n_373)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.A3(n_71),
.B1(n_76),
.B2(n_81),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_101),
.B1(n_105),
.B2(n_107),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_76),
.A2(n_112),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_78),
.Y(n_251)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_80),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_84),
.Y(n_357)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_88),
.B(n_131),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_111),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.Y(n_89)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_90),
.A2(n_99),
.B1(n_112),
.B2(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2x1_ASAP7_75t_SL g292 ( 
.A(n_99),
.B(n_123),
.Y(n_292)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_104),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_149),
.B1(n_152),
.B2(n_155),
.Y(n_148)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_123),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_115),
.Y(n_253)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_158),
.B(n_166),
.Y(n_131)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_132),
.A2(n_240),
.B1(n_241),
.B2(n_246),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_132),
.A2(n_166),
.B(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_133),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_133),
.B(n_168),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_148),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_142),
.B2(n_146),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_139),
.Y(n_236)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_140),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_141),
.Y(n_367)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_145),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_151),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_158),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_167),
.Y(n_311)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_173),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_173),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_254),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_238),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_177),
.B(n_191),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_189),
.B2(n_190),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_181),
.A2(n_189),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_188),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_189),
.A2(n_424),
.B(n_435),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_202),
.B1(n_228),
.B2(n_237),
.Y(n_191)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_201),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_201),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_201),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_201),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_202),
.A2(n_228),
.B1(n_237),
.B2(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_202),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_SL g376 ( 
.A1(n_202),
.A2(n_377),
.B(n_385),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_202),
.A2(n_237),
.B1(n_377),
.B2(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_202),
.A2(n_402),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_217),
.Y(n_202)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_203),
.Y(n_290)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_208),
.B1(n_210),
.B2(n_214),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_210),
.Y(n_468)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_213),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_215),
.Y(n_460)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_216),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_224),
.B2(n_226),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_233),
.Y(n_466)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_247),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_246),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_246),
.B(n_298),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_275),
.A2(n_276),
.B1(n_317),
.B2(n_319),
.Y(n_316)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_281),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_291),
.C(n_299),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_299),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_289),
.B2(n_290),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_283),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_284),
.B(n_290),
.Y(n_385)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_284),
.Y(n_420)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_290),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_298),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_298),
.B(n_463),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_SL g479 ( 
.A1(n_298),
.A2(n_462),
.B(n_480),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_298),
.B(n_419),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_298),
.B(n_492),
.Y(n_491)
);

AOI22x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_310),
.B2(n_311),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_342),
.B(n_510),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_316),
.B(n_320),
.Y(n_510)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.C(n_324),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_321),
.B(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_323),
.B(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.C(n_340),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_388),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B(n_329),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_330),
.A2(n_340),
.B1(n_341),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_369),
.B(n_371),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx12f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_392),
.B(n_508),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_390),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_346),
.B(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_375),
.C(n_386),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_375),
.B1(n_376),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_368),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_366),
.Y(n_482)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_368),
.B(n_400),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_369),
.A2(n_371),
.B(n_443),
.Y(n_487)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_380),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_385),
.B(n_478),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

AOI21x1_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_436),
.B(n_507),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_414),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_398),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.C(n_407),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_407),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_415),
.Y(n_505)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.C(n_423),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_418),
.B(n_422),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_423),
.B(n_500),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_424),
.Y(n_455)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_503),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_498),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_483),
.B(n_497),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_456),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_456),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_454),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_477),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_457),
.B(n_477),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_461),
.B1(n_467),
.B2(n_469),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_460),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_474),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_488),
.B(n_496),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_486),
.B(n_487),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_501),
.Y(n_498)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_499),
.Y(n_506)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_503)
);


endmodule