module real_jpeg_1119_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_68),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g211 ( 
.A1(n_1),
.A2(n_43),
.B1(n_46),
.B2(n_68),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_2),
.B(n_55),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_2),
.B(n_81),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_2),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_2),
.A2(n_55),
.B(n_184),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_27),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_2),
.A2(n_34),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_2),
.B(n_43),
.C(n_45),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_2),
.B(n_99),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_2),
.B(n_41),
.Y(n_275)
);

BUFx4f_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_4),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_194),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_194),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_4),
.A2(n_43),
.B1(n_46),
.B2(n_194),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_63),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_5),
.A2(n_43),
.B1(n_46),
.B2(n_63),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_36),
.B1(n_55),
.B2(n_56),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_36),
.B1(n_43),
.B2(n_46),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_9),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_110),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_110),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_9),
.A2(n_43),
.B1(n_46),
.B2(n_110),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_10),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_149),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_149),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_13),
.A2(n_43),
.B1(n_46),
.B2(n_149),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_14),
.A2(n_55),
.B1(n_56),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_14),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_175),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_14),
.A2(n_43),
.B1(n_46),
.B2(n_175),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_16),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_16),
.A2(n_43),
.B1(n_46),
.B2(n_65),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_74),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.C(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_22),
.A2(n_66),
.B1(n_118),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_22),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_50),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_40),
.C(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_26),
.A2(n_37),
.B1(n_115),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_26),
.A2(n_37),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_26),
.A2(n_37),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_26),
.A2(n_37),
.B1(n_190),
.B2(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_26),
.A2(n_37),
.B1(n_205),
.B2(n_252),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_27),
.A2(n_72),
.B(n_77),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_27),
.A2(n_71),
.B1(n_72),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_27),
.A2(n_72),
.B1(n_145),
.B2(n_172),
.Y(n_171)
);

AO22x2_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_29),
.B1(n_44),
.B2(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_28),
.B(n_31),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_29),
.A2(n_30),
.A3(n_34),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_29),
.B(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_33),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_34),
.B1(n_58),
.B2(n_60),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_33),
.B(n_58),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_33),
.B(n_220),
.Y(n_219)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_34),
.A2(n_56),
.A3(n_60),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_66),
.C(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_40),
.A2(n_50),
.B1(n_70),
.B2(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_49),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_47),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_106),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_41),
.A2(n_47),
.B1(n_105),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_41),
.A2(n_47),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_41),
.A2(n_47),
.B1(n_216),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_41),
.A2(n_47),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_41),
.A2(n_47),
.B1(n_243),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_42),
.A2(n_142),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_42),
.A2(n_168),
.B1(n_215),
.B2(n_255),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_43),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_43),
.B(n_271),
.Y(n_270)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_47),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_61),
.B1(n_62),
.B2(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_52),
.A2(n_61),
.B1(n_67),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_52),
.A2(n_61),
.B1(n_109),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_52),
.A2(n_61),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_52),
.A2(n_61),
.B1(n_193),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_53),
.A2(n_81),
.B1(n_148),
.B2(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_69),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_155),
.B(n_310),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_150),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_124),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_91),
.B(n_124),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_111),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_92),
.B(n_117),
.C(n_122),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_107),
.B(n_108),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_94),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_107),
.B1(n_108),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_95),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_101),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_96),
.A2(n_98),
.B1(n_138),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_96),
.A2(n_98),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_96),
.A2(n_98),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_99),
.B1(n_102),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_97),
.A2(n_99),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_97),
.A2(n_99),
.B1(n_187),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_97),
.A2(n_99),
.B1(n_224),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_97),
.A2(n_99),
.B1(n_220),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_97),
.A2(n_99),
.B1(n_273),
.B2(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_117),
.B1(n_122),
.B2(n_123),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_113),
.B(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_132),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.C(n_146),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_134),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_146),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_150),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_151),
.B(n_154),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_176),
.B(n_309),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_157),
.B(n_159),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.C(n_173),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_166),
.B(n_169),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_173),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_199),
.B(n_308),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_197),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_178),
.B(n_197),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_196),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_196),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_181),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.C(n_192),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_182),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_186),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_189),
.B(n_192),
.Y(n_299)
);

AOI31xp33_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_293),
.A3(n_302),
.B(n_305),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_238),
.B(n_292),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_226),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_202),
.B(n_226),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_213),
.C(n_217),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_203),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_213),
.B(n_217),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_303),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.CI(n_229),
.CON(n_226),
.SN(n_226)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_233),
.C(n_237),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_287),
.B(n_291),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_256),
.B(n_286),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_245),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_267),
.B(n_285),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_279),
.B(n_284),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B(n_278),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);


endmodule