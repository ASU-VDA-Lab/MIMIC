module real_aes_10068_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1699;
wire n_1023;
wire n_730;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_1691;
wire n_640;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AO221x1_ASAP7_75t_L g1502 ( .A1(n_0), .A2(n_134), .B1(n_1458), .B2(n_1503), .C(n_1505), .Y(n_1502) );
INVxp67_ASAP7_75t_SL g1368 ( .A(n_1), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_1), .A2(n_10), .B1(n_498), .B2(n_1384), .Y(n_1383) );
INVxp33_ASAP7_75t_L g664 ( .A(n_2), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_2), .A2(n_633), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g1406 ( .A(n_3), .Y(n_1406) );
AOI22xp5_ASAP7_75t_L g1491 ( .A1(n_4), .A2(n_122), .B1(n_1458), .B2(n_1462), .Y(n_1491) );
INVx1_ASAP7_75t_L g1173 ( .A(n_5), .Y(n_1173) );
AOI22xp33_ASAP7_75t_SL g974 ( .A1(n_6), .A2(n_17), .B1(n_654), .B2(n_731), .Y(n_974) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_6), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_7), .A2(n_167), .B1(n_520), .B2(n_822), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_7), .A2(n_167), .B1(n_433), .B2(n_441), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_8), .A2(n_224), .B1(n_538), .B2(n_802), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_8), .A2(n_224), .B1(n_520), .B2(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1360 ( .A(n_9), .Y(n_1360) );
INVx1_ASAP7_75t_L g1367 ( .A(n_10), .Y(n_1367) );
OAI22xp5_ASAP7_75t_L g1743 ( .A1(n_11), .A2(n_99), .B1(n_418), .B2(n_423), .Y(n_1743) );
INVx1_ASAP7_75t_L g1777 ( .A(n_11), .Y(n_1777) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_12), .A2(n_283), .B1(n_617), .B2(n_618), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_12), .A2(n_283), .B1(n_642), .B2(n_643), .Y(n_641) );
INVxp33_ASAP7_75t_SL g970 ( .A(n_13), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_13), .A2(n_308), .B1(n_617), .B2(n_984), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_14), .Y(n_886) );
INVx1_ASAP7_75t_L g1018 ( .A(n_15), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_15), .A2(n_70), .B1(n_502), .B2(n_871), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g966 ( .A(n_16), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_16), .A2(n_218), .B1(n_462), .B2(n_997), .Y(n_996) );
INVxp67_ASAP7_75t_SL g1002 ( .A(n_17), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_18), .A2(n_217), .B1(n_844), .B2(n_1324), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_18), .A2(n_217), .B1(n_519), .B2(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g612 ( .A(n_19), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_19), .A2(n_60), .B1(n_623), .B2(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g1359 ( .A(n_20), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_20), .A2(n_66), .B1(n_871), .B2(n_1194), .Y(n_1386) );
INVx1_ASAP7_75t_L g1506 ( .A(n_21), .Y(n_1506) );
INVxp33_ASAP7_75t_SL g599 ( .A(n_22), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_22), .A2(n_103), .B1(n_650), .B2(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g1317 ( .A(n_23), .Y(n_1317) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_23), .A2(n_235), .B1(n_1082), .B2(n_1184), .Y(n_1345) );
INVx1_ASAP7_75t_L g1136 ( .A(n_24), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_24), .A2(n_313), .B1(n_418), .B2(n_423), .Y(n_1150) );
XOR2x2_ASAP7_75t_L g957 ( .A(n_25), .B(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g1268 ( .A(n_26), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_27), .A2(n_78), .B1(n_787), .B2(n_790), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_27), .A2(n_78), .B1(n_811), .B2(n_814), .Y(n_810) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_28), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_28), .A2(n_214), .B1(n_729), .B2(n_731), .Y(n_1209) );
AOI22xp33_ASAP7_75t_SL g1028 ( .A1(n_29), .A2(n_247), .B1(n_538), .B2(n_802), .Y(n_1028) );
AOI22xp33_ASAP7_75t_SL g1039 ( .A1(n_29), .A2(n_247), .B1(n_552), .B2(n_556), .Y(n_1039) );
INVx1_ASAP7_75t_L g763 ( .A(n_30), .Y(n_763) );
INVx1_ASAP7_75t_L g1704 ( .A(n_31), .Y(n_1704) );
AOI22xp33_ASAP7_75t_SL g1717 ( .A1(n_31), .A2(n_197), .B1(n_822), .B2(n_823), .Y(n_1717) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_32), .Y(n_940) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_33), .A2(n_87), .B1(n_844), .B2(n_1092), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_33), .A2(n_87), .B1(n_729), .B2(n_745), .Y(n_1106) );
INVx1_ASAP7_75t_L g1262 ( .A(n_34), .Y(n_1262) );
INVx1_ASAP7_75t_L g1007 ( .A(n_35), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g1044 ( .A1(n_35), .A2(n_157), .B1(n_822), .B2(n_823), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_36), .Y(n_941) );
INVx1_ASAP7_75t_L g896 ( .A(n_37), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_37), .A2(n_184), .B1(n_433), .B2(n_441), .Y(n_942) );
INVx1_ASAP7_75t_L g595 ( .A(n_38), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g1742 ( .A(n_39), .B(n_841), .Y(n_1742) );
INVx1_ASAP7_75t_L g1775 ( .A(n_39), .Y(n_1775) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_40), .A2(n_339), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
INVxp67_ASAP7_75t_SL g1348 ( .A(n_40), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_41), .A2(n_116), .B1(n_479), .B2(n_484), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_41), .A2(n_116), .B1(n_729), .B2(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g350 ( .A(n_42), .Y(n_350) );
XNOR2xp5_ASAP7_75t_L g876 ( .A(n_43), .B(n_877), .Y(n_876) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_44), .A2(n_226), .B1(n_844), .B2(n_845), .C(n_846), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_44), .A2(n_226), .B1(n_822), .B2(n_823), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_45), .A2(n_64), .B1(n_359), .B2(n_470), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_45), .A2(n_332), .B1(n_418), .B2(n_423), .Y(n_583) );
XNOR2xp5_ASAP7_75t_L g1398 ( .A(n_46), .B(n_1399), .Y(n_1398) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_47), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_47), .A2(n_190), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_48), .A2(n_143), .B1(n_1458), .B2(n_1462), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1224 ( .A1(n_49), .A2(n_119), .B1(n_418), .B2(n_840), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1240 ( .A1(n_49), .A2(n_119), .B1(n_617), .B2(n_621), .Y(n_1240) );
AOI22xp33_ASAP7_75t_SL g1321 ( .A1(n_50), .A2(n_187), .B1(n_794), .B2(n_1322), .Y(n_1321) );
AOI22xp33_ASAP7_75t_SL g1335 ( .A1(n_50), .A2(n_187), .B1(n_652), .B2(n_1336), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_51), .A2(n_333), .B1(n_1097), .B2(n_1238), .Y(n_1237) );
AOI22xp33_ASAP7_75t_SL g1248 ( .A1(n_51), .A2(n_227), .B1(n_643), .B2(n_1249), .Y(n_1248) );
INVxp33_ASAP7_75t_L g1087 ( .A(n_52), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_52), .A2(n_280), .B1(n_514), .B2(n_1105), .Y(n_1108) );
INVxp67_ASAP7_75t_SL g610 ( .A(n_53), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_53), .A2(n_279), .B1(n_617), .B2(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g1401 ( .A1(n_54), .A2(n_329), .B1(n_418), .B2(n_840), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g1416 ( .A1(n_54), .A2(n_239), .B1(n_799), .B2(n_984), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_55), .A2(n_298), .B1(n_538), .B2(n_539), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_55), .A2(n_298), .B1(n_518), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g1708 ( .A1(n_56), .A2(n_192), .B1(n_541), .B2(n_871), .Y(n_1708) );
AOI22xp33_ASAP7_75t_L g1713 ( .A1(n_56), .A2(n_192), .B1(n_527), .B2(n_550), .Y(n_1713) );
INVxp33_ASAP7_75t_SL g1174 ( .A(n_57), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_57), .A2(n_195), .B1(n_498), .B2(n_499), .Y(n_1192) );
INVxp33_ASAP7_75t_SL g1189 ( .A(n_58), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_58), .A2(n_74), .B1(n_779), .B2(n_1204), .Y(n_1208) );
AO221x2_ASAP7_75t_L g1589 ( .A1(n_59), .A2(n_260), .B1(n_1503), .B2(n_1590), .C(n_1592), .Y(n_1589) );
INVxp33_ASAP7_75t_SL g605 ( .A(n_60), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_61), .A2(n_84), .B1(n_433), .B2(n_441), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_61), .A2(n_84), .B1(n_518), .B2(n_519), .Y(n_529) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_62), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_62), .A2(n_72), .B1(n_820), .B2(n_823), .Y(n_819) );
INVxp33_ASAP7_75t_SL g1231 ( .A(n_63), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_63), .A2(n_160), .B1(n_642), .B2(n_643), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_64), .A2(n_180), .B1(n_559), .B2(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g864 ( .A(n_65), .Y(n_864) );
INVx1_ASAP7_75t_L g1362 ( .A(n_66), .Y(n_1362) );
INVx1_ASAP7_75t_L g1371 ( .A(n_67), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_67), .A2(n_245), .B1(n_514), .B2(n_827), .Y(n_1394) );
OAI211xp5_ASAP7_75t_L g833 ( .A1(n_68), .A2(n_413), .B(n_834), .C(n_836), .Y(n_833) );
INVx1_ASAP7_75t_L g856 ( .A(n_68), .Y(n_856) );
INVx1_ASAP7_75t_L g1010 ( .A(n_69), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_69), .A2(n_169), .B1(n_900), .B2(n_1042), .Y(n_1041) );
OAI211xp5_ASAP7_75t_L g1049 ( .A1(n_69), .A2(n_453), .B(n_1050), .C(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1022 ( .A(n_70), .Y(n_1022) );
OAI211xp5_ASAP7_75t_L g1055 ( .A1(n_70), .A2(n_413), .B(n_1056), .C(n_1058), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1465 ( .A1(n_71), .A2(n_291), .B1(n_1458), .B2(n_1462), .Y(n_1465) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_72), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g1490 ( .A1(n_73), .A2(n_324), .B1(n_1446), .B2(n_1454), .Y(n_1490) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_74), .Y(n_1182) );
INVx1_ASAP7_75t_L g1260 ( .A(n_75), .Y(n_1260) );
INVx1_ASAP7_75t_L g1019 ( .A(n_76), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_76), .A2(n_318), .B1(n_498), .B2(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g570 ( .A(n_77), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_79), .Y(n_1154) );
AO22x1_ASAP7_75t_L g1468 ( .A1(n_80), .A2(n_244), .B1(n_1462), .B2(n_1469), .Y(n_1468) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_81), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_81), .A2(n_264), .B1(n_729), .B2(n_745), .Y(n_744) );
XOR2xp5_ASAP7_75t_L g1212 ( .A(n_82), .B(n_1213), .Y(n_1212) );
AO22x1_ASAP7_75t_L g1470 ( .A1(n_82), .A2(n_242), .B1(n_1446), .B2(n_1454), .Y(n_1470) );
INVx1_ASAP7_75t_L g1219 ( .A(n_83), .Y(n_1219) );
OAI222xp33_ASAP7_75t_L g1228 ( .A1(n_83), .A2(n_177), .B1(n_262), .B2(n_704), .C1(n_765), .C2(n_1082), .Y(n_1228) );
OAI21xp33_ASAP7_75t_SL g1217 ( .A1(n_85), .A2(n_883), .B(n_1218), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_85), .A2(n_293), .B1(n_499), .B2(n_1242), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_86), .A2(n_95), .B1(n_503), .B2(n_1200), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_86), .A2(n_95), .B1(n_779), .B2(n_1204), .Y(n_1203) );
BUFx2_ASAP7_75t_L g430 ( .A(n_88), .Y(n_430) );
BUFx2_ASAP7_75t_L g473 ( .A(n_88), .Y(n_473) );
INVx1_ASAP7_75t_L g509 ( .A(n_88), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_89), .A2(n_184), .B1(n_898), .B2(n_900), .Y(n_897) );
OAI211xp5_ASAP7_75t_L g935 ( .A1(n_89), .A2(n_453), .B(n_936), .C(n_939), .Y(n_935) );
INVx1_ASAP7_75t_L g1315 ( .A(n_90), .Y(n_1315) );
AOI22xp33_ASAP7_75t_SL g1327 ( .A1(n_90), .A2(n_191), .B1(n_794), .B2(n_1328), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_91), .A2(n_241), .B1(n_636), .B2(n_639), .Y(n_973) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_91), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g1412 ( .A1(n_92), .A2(n_230), .B1(n_794), .B2(n_1413), .Y(n_1412) );
AOI22xp33_ASAP7_75t_SL g1419 ( .A1(n_92), .A2(n_230), .B1(n_652), .B2(n_1251), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_93), .A2(n_336), .B1(n_729), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_93), .A2(n_336), .B1(n_617), .B2(n_627), .Y(n_987) );
INVx1_ASAP7_75t_L g1176 ( .A(n_94), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_94), .A2(n_114), .B1(n_491), .B2(n_1194), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_96), .A2(n_311), .B1(n_491), .B2(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_96), .A2(n_311), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_97), .A2(n_272), .B1(n_639), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_97), .A2(n_272), .B1(n_623), .B2(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1690 ( .A(n_98), .Y(n_1690) );
AOI22xp33_ASAP7_75t_L g1710 ( .A1(n_98), .A2(n_340), .B1(n_789), .B2(n_802), .Y(n_1710) );
INVx1_ASAP7_75t_L g1738 ( .A(n_99), .Y(n_1738) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_100), .A2(n_269), .B1(n_498), .B2(n_1197), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_100), .A2(n_269), .B1(n_557), .B2(n_1206), .Y(n_1205) );
XNOR2xp5_ASAP7_75t_L g374 ( .A(n_101), .B(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_102), .A2(n_301), .B1(n_491), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_102), .A2(n_301), .B1(n_561), .B2(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g594 ( .A(n_103), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_104), .Y(n_1011) );
OAI22xp33_ASAP7_75t_L g839 ( .A1(n_105), .A2(n_240), .B1(n_840), .B2(n_841), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g851 ( .A1(n_105), .A2(n_240), .B1(n_787), .B2(n_800), .C(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g931 ( .A(n_106), .Y(n_931) );
OAI211xp5_ASAP7_75t_SL g946 ( .A1(n_106), .A2(n_674), .B(n_947), .C(n_949), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_107), .A2(n_227), .B1(n_989), .B2(n_1235), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_107), .A2(n_333), .B1(n_1245), .B2(n_1247), .Y(n_1244) );
INVx1_ASAP7_75t_L g1293 ( .A(n_108), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1694 ( .A1(n_109), .A2(n_117), .B1(n_1365), .B2(n_1695), .Y(n_1694) );
OAI22xp5_ASAP7_75t_L g1699 ( .A1(n_109), .A2(n_117), .B1(n_462), .B2(n_997), .Y(n_1699) );
AO221x1_ASAP7_75t_L g1475 ( .A1(n_110), .A2(n_126), .B1(n_1458), .B2(n_1462), .C(n_1476), .Y(n_1475) );
AO221x1_ASAP7_75t_L g1483 ( .A1(n_111), .A2(n_305), .B1(n_1458), .B2(n_1462), .C(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g584 ( .A(n_112), .Y(n_584) );
INVx1_ASAP7_75t_L g847 ( .A(n_113), .Y(n_847) );
INVxp33_ASAP7_75t_SL g1170 ( .A(n_114), .Y(n_1170) );
INVx1_ASAP7_75t_L g1287 ( .A(n_115), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_118), .A2(n_151), .B1(n_487), .B2(n_1030), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_118), .A2(n_151), .B1(n_514), .B2(n_827), .Y(n_1038) );
INVx1_ASAP7_75t_L g1272 ( .A(n_120), .Y(n_1272) );
OAI22xp33_ASAP7_75t_SL g1299 ( .A1(n_120), .A2(n_216), .B1(n_359), .B2(n_433), .Y(n_1299) );
INVx1_ASAP7_75t_L g1480 ( .A(n_121), .Y(n_1480) );
AOI22xp33_ASAP7_75t_L g1723 ( .A1(n_122), .A2(n_1724), .B1(n_1729), .B2(n_1784), .Y(n_1723) );
OA22x2_ASAP7_75t_L g1731 ( .A1(n_122), .A2(n_1732), .B1(n_1782), .B2(n_1783), .Y(n_1731) );
INVxp67_ASAP7_75t_SL g1783 ( .A(n_122), .Y(n_1783) );
AOI22xp33_ASAP7_75t_L g1424 ( .A1(n_123), .A2(n_222), .B1(n_1339), .B2(n_1425), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g1433 ( .A1(n_123), .A2(n_222), .B1(n_433), .B2(n_441), .Y(n_1433) );
INVx1_ASAP7_75t_L g838 ( .A(n_124), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_125), .A2(n_148), .B1(n_1446), .B2(n_1454), .Y(n_1445) );
INVxp33_ASAP7_75t_SL g1084 ( .A(n_127), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_127), .A2(n_215), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
XOR2xp5_ASAP7_75t_L g1119 ( .A(n_128), .B(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1593 ( .A(n_129), .Y(n_1593) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_130), .A2(n_239), .B1(n_423), .B2(n_841), .Y(n_1402) );
INVxp33_ASAP7_75t_SL g1432 ( .A(n_130), .Y(n_1432) );
INVxp33_ASAP7_75t_L g772 ( .A(n_131), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_131), .A2(n_183), .B1(n_794), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_132), .A2(n_287), .B1(n_632), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_132), .A2(n_287), .B1(n_636), .B2(n_1105), .Y(n_1104) );
INVxp33_ASAP7_75t_SL g1070 ( .A(n_133), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_133), .A2(n_330), .B1(n_1097), .B2(n_1099), .Y(n_1096) );
INVx1_ASAP7_75t_L g1283 ( .A(n_135), .Y(n_1283) );
OAI22xp33_ASAP7_75t_L g1289 ( .A1(n_135), .A2(n_142), .B1(n_418), .B2(n_840), .Y(n_1289) );
INVx1_ASAP7_75t_L g758 ( .A(n_136), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_137), .A2(n_207), .B1(n_888), .B2(n_890), .Y(n_887) );
INVx1_ASAP7_75t_L g915 ( .A(n_137), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g1739 ( .A(n_138), .Y(n_1739) );
INVx1_ASAP7_75t_L g1134 ( .A(n_139), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_139), .A2(n_281), .B1(n_840), .B2(n_841), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_140), .A2(n_587), .B1(n_658), .B2(n_659), .Y(n_586) );
INVxp67_ASAP7_75t_L g658 ( .A(n_140), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_141), .A2(n_181), .B1(n_359), .B2(n_470), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g1250 ( .A1(n_141), .A2(n_262), .B1(n_1247), .B2(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1286 ( .A(n_142), .Y(n_1286) );
INVx1_ASAP7_75t_L g1450 ( .A(n_144), .Y(n_1450) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_145), .A2(n_448), .B(n_453), .C(n_460), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_145), .A2(n_250), .B1(n_515), .B2(n_527), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g1688 ( .A(n_146), .Y(n_1688) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_147), .A2(n_223), .B1(n_477), .B2(n_482), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_147), .A2(n_223), .B1(n_518), .B2(n_519), .Y(n_517) );
XOR2x2_ASAP7_75t_L g1305 ( .A(n_148), .B(n_1306), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_149), .A2(n_236), .B1(n_1030), .B2(n_1194), .Y(n_1381) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_149), .A2(n_236), .B1(n_900), .B2(n_1389), .Y(n_1388) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_150), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g1485 ( .A(n_152), .Y(n_1485) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_153), .Y(n_761) );
INVx1_ASAP7_75t_L g1076 ( .A(n_154), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_154), .A2(n_277), .B1(n_765), .B2(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1146 ( .A(n_155), .Y(n_1146) );
OAI22xp33_ASAP7_75t_SL g1161 ( .A1(n_155), .A2(n_164), .B1(n_359), .B2(n_433), .Y(n_1161) );
INVxp33_ASAP7_75t_SL g961 ( .A(n_156), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_156), .A2(n_162), .B1(n_621), .B2(n_623), .Y(n_985) );
INVx1_ASAP7_75t_L g1008 ( .A(n_157), .Y(n_1008) );
INVx1_ASAP7_75t_L g1451 ( .A(n_158), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_158), .B(n_1449), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_159), .Y(n_1012) );
INVxp33_ASAP7_75t_L g1230 ( .A(n_160), .Y(n_1230) );
INVx2_ASAP7_75t_L g362 ( .A(n_161), .Y(n_362) );
INVxp67_ASAP7_75t_SL g964 ( .A(n_162), .Y(n_964) );
INVxp33_ASAP7_75t_L g1069 ( .A(n_163), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_163), .A2(n_320), .B1(n_624), .B2(n_1102), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_164), .A2(n_276), .B1(n_518), .B2(n_520), .Y(n_1148) );
AOI22xp33_ASAP7_75t_SL g1337 ( .A1(n_165), .A2(n_295), .B1(n_779), .B2(n_808), .Y(n_1337) );
INVxp33_ASAP7_75t_SL g1350 ( .A(n_165), .Y(n_1350) );
CKINVDCx5p33_ASAP7_75t_R g1754 ( .A(n_166), .Y(n_1754) );
BUFx3_ASAP7_75t_L g384 ( .A(n_168), .Y(n_384) );
INVx1_ASAP7_75t_L g411 ( .A(n_168), .Y(n_411) );
INVx1_ASAP7_75t_L g1014 ( .A(n_169), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g1747 ( .A(n_170), .Y(n_1747) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_171), .A2(n_175), .B1(n_652), .B2(n_1336), .Y(n_1423) );
INVx1_ASAP7_75t_L g1431 ( .A(n_171), .Y(n_1431) );
INVx1_ASAP7_75t_L g671 ( .A(n_172), .Y(n_671) );
INVx1_ASAP7_75t_L g668 ( .A(n_173), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g1707 ( .A1(n_174), .A2(n_229), .B1(n_538), .B2(n_802), .Y(n_1707) );
AOI22xp33_ASAP7_75t_SL g1714 ( .A1(n_174), .A2(n_229), .B1(n_520), .B2(n_822), .Y(n_1714) );
INVx1_ASAP7_75t_L g1429 ( .A(n_175), .Y(n_1429) );
CKINVDCx5p33_ASAP7_75t_R g1740 ( .A(n_176), .Y(n_1740) );
INVx1_ASAP7_75t_L g1220 ( .A(n_177), .Y(n_1220) );
INVx1_ASAP7_75t_L g1687 ( .A(n_178), .Y(n_1687) );
AOI22xp33_ASAP7_75t_L g1711 ( .A1(n_178), .A2(n_296), .B1(n_541), .B2(n_871), .Y(n_1711) );
INVxp33_ASAP7_75t_L g767 ( .A(n_179), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_179), .A2(n_234), .B1(n_808), .B2(n_825), .Y(n_824) );
OAI211xp5_ASAP7_75t_SL g565 ( .A1(n_180), .A2(n_453), .B(n_566), .C(n_569), .Y(n_565) );
INVx1_ASAP7_75t_L g1222 ( .A(n_181), .Y(n_1222) );
INVxp33_ASAP7_75t_L g666 ( .A(n_182), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_182), .A2(n_288), .B1(n_477), .B2(n_499), .C(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g777 ( .A(n_183), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_185), .A2(n_314), .B1(n_799), .B2(n_1410), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_185), .A2(n_314), .B1(n_1245), .B2(n_1340), .Y(n_1420) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_186), .A2(n_332), .B1(n_487), .B2(n_491), .Y(n_545) );
INVx1_ASAP7_75t_L g576 ( .A(n_186), .Y(n_576) );
INVx1_ASAP7_75t_L g1507 ( .A(n_188), .Y(n_1507) );
INVx1_ASAP7_75t_L g395 ( .A(n_189), .Y(n_395) );
INVx1_ASAP7_75t_L g412 ( .A(n_190), .Y(n_412) );
INVxp33_ASAP7_75t_SL g1309 ( .A(n_191), .Y(n_1309) );
INVx1_ASAP7_75t_L g1273 ( .A(n_193), .Y(n_1273) );
OAI211xp5_ASAP7_75t_SL g1297 ( .A1(n_193), .A2(n_448), .B(n_453), .C(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1595 ( .A(n_194), .Y(n_1595) );
INVxp33_ASAP7_75t_SL g1171 ( .A(n_195), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_196), .A2(n_278), .B1(n_418), .B2(n_423), .Y(n_832) );
INVx1_ASAP7_75t_L g873 ( .A(n_196), .Y(n_873) );
INVx1_ASAP7_75t_L g1702 ( .A(n_197), .Y(n_1702) );
INVx1_ASAP7_75t_L g428 ( .A(n_198), .Y(n_428) );
INVx1_ASAP7_75t_L g571 ( .A(n_199), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_200), .A2(n_203), .B1(n_621), .B2(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_200), .A2(n_203), .B1(n_636), .B2(n_639), .Y(n_635) );
INVxp67_ASAP7_75t_L g1377 ( .A(n_201), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_201), .A2(n_282), .B1(n_822), .B2(n_823), .Y(n_1395) );
CKINVDCx5p33_ASAP7_75t_R g1758 ( .A(n_202), .Y(n_1758) );
INVxp67_ASAP7_75t_SL g1130 ( .A(n_204), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_204), .A2(n_319), .B1(n_520), .B2(n_556), .Y(n_1143) );
INVx1_ASAP7_75t_L g926 ( .A(n_205), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_205), .A2(n_209), .B1(n_418), .B2(n_840), .Y(n_944) );
INVx1_ASAP7_75t_L g1477 ( .A(n_206), .Y(n_1477) );
INVx1_ASAP7_75t_L g908 ( .A(n_207), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g1466 ( .A1(n_208), .A2(n_343), .B1(n_1446), .B2(n_1454), .Y(n_1466) );
INVx1_ASAP7_75t_L g922 ( .A(n_209), .Y(n_922) );
CKINVDCx14_ASAP7_75t_R g829 ( .A(n_210), .Y(n_829) );
INVx1_ASAP7_75t_L g837 ( .A(n_211), .Y(n_837) );
INVx1_ASAP7_75t_L g1312 ( .A(n_212), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_213), .A2(n_290), .B1(n_556), .B2(n_557), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_213), .A2(n_290), .B1(n_433), .B2(n_441), .Y(n_564) );
INVxp33_ASAP7_75t_L g1186 ( .A(n_214), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g1085 ( .A(n_215), .Y(n_1085) );
INVx1_ASAP7_75t_L g1275 ( .A(n_216), .Y(n_1275) );
INVxp67_ASAP7_75t_SL g967 ( .A(n_218), .Y(n_967) );
INVx1_ASAP7_75t_L g1126 ( .A(n_219), .Y(n_1126) );
INVx1_ASAP7_75t_L g969 ( .A(n_220), .Y(n_969) );
INVx1_ASAP7_75t_L g386 ( .A(n_221), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_225), .A2(n_256), .B1(n_487), .B2(n_491), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_225), .A2(n_256), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g849 ( .A(n_228), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_231), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g1735 ( .A1(n_232), .A2(n_253), .B1(n_433), .B2(n_441), .Y(n_1735) );
INVx1_ASAP7_75t_L g1765 ( .A(n_232), .Y(n_1765) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_233), .A2(n_266), .B1(n_538), .B2(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g582 ( .A(n_233), .Y(n_582) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_234), .Y(n_762) );
INVx1_ASAP7_75t_L g1318 ( .A(n_235), .Y(n_1318) );
OAI211xp5_ASAP7_75t_L g1736 ( .A1(n_237), .A2(n_453), .B(n_930), .C(n_1737), .Y(n_1736) );
INVx1_ASAP7_75t_L g1762 ( .A(n_237), .Y(n_1762) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_238), .Y(n_700) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_241), .Y(n_999) );
INVx1_ASAP7_75t_L g1276 ( .A(n_243), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_243), .A2(n_252), .B1(n_441), .B2(n_470), .Y(n_1296) );
INVxp33_ASAP7_75t_L g1374 ( .A(n_245), .Y(n_1374) );
BUFx3_ASAP7_75t_L g385 ( .A(n_246), .Y(n_385) );
INVx1_ASAP7_75t_L g404 ( .A(n_246), .Y(n_404) );
INVx1_ASAP7_75t_L g865 ( .A(n_248), .Y(n_865) );
INVxp67_ASAP7_75t_SL g1313 ( .A(n_249), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1326 ( .A1(n_249), .A2(n_257), .B1(n_787), .B2(n_845), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_250), .A2(n_317), .B1(n_359), .B2(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g894 ( .A(n_251), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_251), .A2(n_307), .B1(n_359), .B2(n_470), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_252), .A2(n_259), .B1(n_423), .B2(n_841), .Y(n_1290) );
INVx1_ASAP7_75t_L g1764 ( .A(n_253), .Y(n_1764) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_254), .Y(n_358) );
INVx1_ASAP7_75t_L g511 ( .A(n_254), .Y(n_511) );
AND2x2_ASAP7_75t_L g680 ( .A(n_254), .B(n_437), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_254), .B(n_323), .Y(n_694) );
INVx1_ASAP7_75t_L g673 ( .A(n_255), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_255), .A2(n_342), .B1(n_688), .B2(n_695), .C(n_697), .Y(n_687) );
INVxp33_ASAP7_75t_SL g1310 ( .A(n_257), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1155 ( .A(n_258), .Y(n_1155) );
INVx1_ASAP7_75t_L g1284 ( .A(n_259), .Y(n_1284) );
XNOR2xp5_ASAP7_75t_L g1255 ( .A(n_261), .B(n_1256), .Y(n_1255) );
INVx2_ASAP7_75t_L g390 ( .A(n_263), .Y(n_390) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_264), .Y(n_681) );
INVx1_ASAP7_75t_L g1355 ( .A(n_265), .Y(n_1355) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_266), .Y(n_581) );
INVx1_ASAP7_75t_L g1072 ( .A(n_267), .Y(n_1072) );
INVx1_ASAP7_75t_L g1178 ( .A(n_268), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_268), .A2(n_303), .B1(n_997), .B2(n_1184), .Y(n_1183) );
INVxp33_ASAP7_75t_SL g590 ( .A(n_270), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_270), .A2(n_273), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g1294 ( .A(n_271), .Y(n_1294) );
INVxp33_ASAP7_75t_SL g592 ( .A(n_273), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_274), .A2(n_413), .B(n_742), .C(n_1404), .Y(n_1403) );
AOI22xp33_ASAP7_75t_SL g1417 ( .A1(n_274), .A2(n_329), .B1(n_621), .B2(n_1413), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g1751 ( .A(n_275), .Y(n_1751) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_276), .A2(n_313), .B1(n_441), .B2(n_470), .Y(n_1158) );
INVx1_ASAP7_75t_L g1077 ( .A(n_277), .Y(n_1077) );
INVx1_ASAP7_75t_L g853 ( .A(n_278), .Y(n_853) );
INVxp33_ASAP7_75t_SL g608 ( .A(n_279), .Y(n_608) );
INVxp67_ASAP7_75t_SL g1080 ( .A(n_280), .Y(n_1080) );
INVx1_ASAP7_75t_L g1132 ( .A(n_281), .Y(n_1132) );
INVx1_ASAP7_75t_L g1375 ( .A(n_282), .Y(n_1375) );
AO22x2_ASAP7_75t_L g1003 ( .A1(n_284), .A2(n_1004), .B1(n_1045), .B2(n_1046), .Y(n_1003) );
INVxp67_ASAP7_75t_L g1045 ( .A(n_284), .Y(n_1045) );
CKINVDCx5p33_ASAP7_75t_R g1759 ( .A(n_285), .Y(n_1759) );
INVx1_ASAP7_75t_L g1147 ( .A(n_286), .Y(n_1147) );
OAI211xp5_ASAP7_75t_SL g1159 ( .A1(n_286), .A2(n_448), .B(n_453), .C(n_1160), .Y(n_1159) );
INVxp67_ASAP7_75t_SL g669 ( .A(n_288), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_289), .A2(n_321), .B1(n_1364), .B2(n_1365), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_289), .A2(n_321), .B1(n_997), .B2(n_1184), .Y(n_1372) );
INVx1_ASAP7_75t_L g1701 ( .A(n_292), .Y(n_1701) );
AOI22xp33_ASAP7_75t_L g1716 ( .A1(n_292), .A2(n_326), .B1(n_527), .B2(n_827), .Y(n_1716) );
INVxp67_ASAP7_75t_SL g1223 ( .A(n_293), .Y(n_1223) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_294), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_295), .Y(n_1344) );
INVx1_ASAP7_75t_L g1693 ( .A(n_296), .Y(n_1693) );
INVx1_ASAP7_75t_L g754 ( .A(n_297), .Y(n_754) );
INVx1_ASAP7_75t_L g596 ( .A(n_299), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_300), .A2(n_317), .B1(n_418), .B2(n_423), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_300), .A2(n_331), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g1265 ( .A(n_302), .Y(n_1265) );
INVx1_ASAP7_75t_L g1177 ( .A(n_303), .Y(n_1177) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_304), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_304), .A2(n_325), .B1(n_799), .B2(n_800), .Y(n_798) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_306), .B(n_350), .Y(n_1453) );
AND3x2_ASAP7_75t_L g1461 ( .A(n_306), .B(n_350), .C(n_1450), .Y(n_1461) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_307), .A2(n_335), .B1(n_423), .B2(n_841), .Y(n_945) );
INVxp33_ASAP7_75t_SL g962 ( .A(n_308), .Y(n_962) );
INVx2_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
XOR2xp5_ASAP7_75t_L g1681 ( .A(n_310), .B(n_1682), .Y(n_1681) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_312), .A2(n_505), .B(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_312), .Y(n_727) );
INVx1_ASAP7_75t_L g713 ( .A(n_315), .Y(n_713) );
INVx1_ASAP7_75t_L g601 ( .A(n_316), .Y(n_601) );
INVx1_ASAP7_75t_L g1024 ( .A(n_318), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1128 ( .A(n_319), .Y(n_1128) );
INVxp67_ASAP7_75t_SL g1075 ( .A(n_320), .Y(n_1075) );
INVx1_ASAP7_75t_L g1125 ( .A(n_322), .Y(n_1125) );
INVx1_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
INVx2_ASAP7_75t_L g437 ( .A(n_323), .Y(n_437) );
INVxp67_ASAP7_75t_SL g775 ( .A(n_325), .Y(n_775) );
INVx1_ASAP7_75t_L g1698 ( .A(n_326), .Y(n_1698) );
INVx1_ASAP7_75t_L g711 ( .A(n_327), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g1734 ( .A(n_328), .Y(n_1734) );
INVxp33_ASAP7_75t_L g1073 ( .A(n_330), .Y(n_1073) );
INVx1_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g1744 ( .A1(n_334), .A2(n_413), .B(n_834), .C(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1780 ( .A(n_334), .Y(n_1780) );
INVx1_ASAP7_75t_L g929 ( .A(n_335), .Y(n_929) );
INVx1_ASAP7_75t_L g1405 ( .A(n_337), .Y(n_1405) );
XOR2x2_ASAP7_75t_L g1166 ( .A(n_338), .B(n_1167), .Y(n_1166) );
INVxp33_ASAP7_75t_SL g1347 ( .A(n_339), .Y(n_1347) );
INVx1_ASAP7_75t_L g1691 ( .A(n_340), .Y(n_1691) );
INVx1_ASAP7_75t_L g1138 ( .A(n_341), .Y(n_1138) );
INVx1_ASAP7_75t_L g672 ( .A(n_342), .Y(n_672) );
AO22x1_ASAP7_75t_L g1064 ( .A1(n_343), .A2(n_1065), .B1(n_1066), .B2(n_1112), .Y(n_1064) );
INVxp67_ASAP7_75t_L g1065 ( .A(n_343), .Y(n_1065) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_366), .B(n_1437), .Y(n_344) );
BUFx12f_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
AND2x4_ASAP7_75t_L g1728 ( .A(n_348), .B(n_354), .Y(n_1728) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_SL g1722 ( .A(n_349), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_349), .B(n_351), .Y(n_1789) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_351), .B(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x6_ASAP7_75t_L g472 ( .A(n_356), .B(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_356), .B(n_473), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g495 ( .A(n_357), .B(n_365), .Y(n_495) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g906 ( .A(n_358), .B(n_436), .Y(n_906) );
INVx8_ASAP7_75t_L g600 ( .A(n_359), .Y(n_600) );
OR2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
OR2x6_ASAP7_75t_L g470 ( .A(n_360), .B(n_435), .Y(n_470) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_360), .A2(n_495), .B(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_360), .Y(n_848) );
INVx2_ASAP7_75t_SL g855 ( .A(n_360), .Y(n_855) );
INVx2_ASAP7_75t_SL g918 ( .A(n_360), .Y(n_918) );
BUFx6f_ASAP7_75t_L g1124 ( .A(n_360), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx2_ASAP7_75t_L g440 ( .A(n_362), .Y(n_440) );
AND2x4_ASAP7_75t_L g445 ( .A(n_362), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g452 ( .A(n_362), .Y(n_452) );
INVx1_ASAP7_75t_L g459 ( .A(n_362), .Y(n_459) );
AND2x2_ASAP7_75t_L g490 ( .A(n_362), .B(n_363), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_363), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g446 ( .A(n_363), .Y(n_446) );
INVx1_ASAP7_75t_L g451 ( .A(n_363), .Y(n_451) );
INVx1_ASAP7_75t_L g464 ( .A(n_363), .Y(n_464) );
INVx1_ASAP7_75t_L g481 ( .A(n_363), .Y(n_481) );
AND2x4_ASAP7_75t_L g463 ( .A(n_364), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g997 ( .A(n_365), .B(n_467), .Y(n_997) );
OR2x2_ASAP7_75t_L g1082 ( .A(n_365), .B(n_467), .Y(n_1082) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_1303), .B2(n_1304), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_951), .B1(n_952), .B2(n_1302), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_875), .B2(n_950), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_370), .A2(n_371), .B1(n_875), .B2(n_950), .Y(n_1302) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
XOR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_751), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_585), .B1(n_749), .B2(n_750), .Y(n_372) );
INVx2_ASAP7_75t_L g749 ( .A(n_373), .Y(n_749) );
XOR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_533), .Y(n_373) );
NAND3x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_431), .C(n_474), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_417), .B(n_426), .Y(n_376) );
NAND3xp33_ASAP7_75t_SL g377 ( .A(n_378), .B(n_400), .C(n_413), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_386), .B2(n_387), .C1(n_395), .C2(n_396), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g577 ( .A(n_381), .Y(n_577) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g516 ( .A(n_382), .Y(n_516) );
BUFx3_ASAP7_75t_L g652 ( .A(n_382), .Y(n_652) );
BUFx4f_ASAP7_75t_L g779 ( .A(n_382), .Y(n_779) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_382), .Y(n_827) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g398 ( .A(n_384), .Y(n_398) );
AND2x4_ASAP7_75t_L g403 ( .A(n_384), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g394 ( .A(n_385), .Y(n_394) );
AND2x4_ASAP7_75t_L g410 ( .A(n_385), .B(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_386), .A2(n_395), .B1(n_461), .B2(n_465), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g611 ( .A1(n_387), .A2(n_396), .B1(n_561), .B2(n_595), .C1(n_596), .C2(n_612), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_387), .A2(n_396), .B1(n_652), .B2(n_671), .C1(n_672), .C2(n_673), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g963 ( .A1(n_387), .A2(n_396), .B1(n_964), .B2(n_965), .C1(n_966), .C2(n_967), .Y(n_963) );
AOI222xp33_ASAP7_75t_L g1074 ( .A1(n_387), .A2(n_396), .B1(n_827), .B2(n_1075), .C1(n_1076), .C2(n_1077), .Y(n_1074) );
AOI222xp33_ASAP7_75t_L g1175 ( .A1(n_387), .A2(n_396), .B1(n_639), .B2(n_1176), .C1(n_1177), .C2(n_1178), .Y(n_1175) );
AOI322xp5_ASAP7_75t_L g1745 ( .A1(n_387), .A2(n_396), .A3(n_518), .B1(n_1739), .B2(n_1740), .C1(n_1746), .C2(n_1747), .Y(n_1745) );
AND2x2_ASAP7_75t_SL g387 ( .A(n_388), .B(n_391), .Y(n_387) );
AND2x4_ASAP7_75t_L g424 ( .A(n_388), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g781 ( .A(n_388), .B(n_391), .Y(n_781) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g399 ( .A(n_390), .Y(n_399) );
INVx1_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
AND2x2_ASAP7_75t_L g524 ( .A(n_390), .B(n_428), .Y(n_524) );
INVx2_ASAP7_75t_L g532 ( .A(n_390), .Y(n_532) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g579 ( .A(n_392), .Y(n_579) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g425 ( .A(n_394), .B(n_398), .Y(n_425) );
AOI222xp33_ASAP7_75t_L g575 ( .A1(n_396), .A2(n_570), .B1(n_571), .B2(n_576), .C1(n_577), .C2(n_578), .Y(n_575) );
AOI222xp33_ASAP7_75t_L g776 ( .A1(n_396), .A2(n_761), .B1(n_763), .B2(n_777), .C1(n_778), .C2(n_780), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_396), .A2(n_781), .B1(n_837), .B2(n_838), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_396), .A2(n_781), .B1(n_940), .B2(n_941), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g1020 ( .A1(n_396), .A2(n_780), .B1(n_1011), .B2(n_1012), .C1(n_1021), .C2(n_1022), .Y(n_1020) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_396), .A2(n_781), .B1(n_1011), .B2(n_1012), .Y(n_1058) );
AOI222xp33_ASAP7_75t_L g1152 ( .A1(n_396), .A2(n_578), .B1(n_1138), .B2(n_1153), .C1(n_1154), .C2(n_1155), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_396), .A2(n_578), .B1(n_1219), .B2(n_1220), .Y(n_1218) );
AOI222xp33_ASAP7_75t_L g1292 ( .A1(n_396), .A2(n_578), .B1(n_1105), .B2(n_1287), .C1(n_1293), .C2(n_1294), .Y(n_1292) );
AOI222xp33_ASAP7_75t_L g1314 ( .A1(n_396), .A2(n_780), .B1(n_1315), .B2(n_1316), .C1(n_1317), .C2(n_1318), .Y(n_1314) );
INVx3_ASAP7_75t_L g1365 ( .A(n_396), .Y(n_1365) );
AOI22xp33_ASAP7_75t_SL g1404 ( .A1(n_396), .A2(n_781), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
AND2x6_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_399), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_405), .B1(n_406), .B2(n_412), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_401), .A2(n_406), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_401), .A2(n_605), .B1(n_606), .B2(n_608), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_401), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_401), .A2(n_606), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx6p67_ASAP7_75t_R g840 ( .A(n_401), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_401), .A2(n_414), .B1(n_606), .B2(n_961), .C(n_962), .Y(n_960) );
AOI22xp5_ASAP7_75t_SL g1017 ( .A1(n_401), .A2(n_665), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_401), .A2(n_665), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_401), .A2(n_606), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_401), .A2(n_665), .B1(n_1309), .B2(n_1310), .Y(n_1308) );
AOI22xp5_ASAP7_75t_L g1366 ( .A1(n_401), .A2(n_406), .B1(n_1367), .B2(n_1368), .Y(n_1366) );
AOI22xp5_ASAP7_75t_L g1689 ( .A1(n_401), .A2(n_406), .B1(n_1690), .B2(n_1691), .Y(n_1689) );
AND2x6_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g415 ( .A(n_402), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_402), .Y(n_419) );
AND2x2_ASAP7_75t_L g835 ( .A(n_402), .B(n_550), .Y(n_835) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_403), .Y(n_518) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_403), .Y(n_556) );
BUFx2_ASAP7_75t_L g642 ( .A(n_403), .Y(n_642) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_403), .Y(n_730) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_403), .Y(n_813) );
BUFx3_ASAP7_75t_L g822 ( .A(n_403), .Y(n_822) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_403), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1206 ( .A(n_403), .Y(n_1206) );
INVx2_ASAP7_75t_SL g1392 ( .A(n_403), .Y(n_1392) );
INVx1_ASAP7_75t_L g422 ( .A(n_404), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_406), .A2(n_424), .B1(n_601), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_406), .A2(n_424), .B1(n_668), .B2(n_669), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_406), .A2(n_424), .B1(n_758), .B2(n_775), .Y(n_774) );
INVx4_ASAP7_75t_L g841 ( .A(n_406), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_406), .A2(n_424), .B1(n_969), .B2(n_970), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g1023 ( .A1(n_406), .A2(n_424), .B1(n_1015), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_406), .A2(n_424), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_406), .A2(n_424), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_406), .A2(n_424), .B1(n_1222), .B2(n_1223), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_406), .A2(n_424), .B1(n_1312), .B2(n_1313), .Y(n_1311) );
AND2x6_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
AND2x4_ASAP7_75t_L g606 ( .A(n_407), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g665 ( .A(n_407), .B(n_607), .Y(n_665) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g578 ( .A(n_408), .B(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_409), .Y(n_557) );
INVx1_ASAP7_75t_L g746 ( .A(n_409), .Y(n_746) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_409), .Y(n_823) );
INVx2_ASAP7_75t_L g891 ( .A(n_409), .Y(n_891) );
INVx1_ASAP7_75t_L g981 ( .A(n_409), .Y(n_981) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_410), .Y(n_520) );
INVx1_ASAP7_75t_L g553 ( .A(n_410), .Y(n_553) );
INVx1_ASAP7_75t_L g644 ( .A(n_410), .Y(n_644) );
INVx2_ASAP7_75t_L g734 ( .A(n_410), .Y(n_734) );
INVx1_ASAP7_75t_L g421 ( .A(n_411), .Y(n_421) );
NAND3xp33_ASAP7_75t_SL g574 ( .A(n_413), .B(n_575), .C(n_580), .Y(n_574) );
NAND4xp25_ASAP7_75t_SL g603 ( .A(n_413), .B(n_604), .C(n_609), .D(n_611), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g1151 ( .A(n_413), .B(n_1152), .Y(n_1151) );
NAND4xp25_ASAP7_75t_L g1168 ( .A(n_413), .B(n_1169), .C(n_1172), .D(n_1175), .Y(n_1168) );
NAND2xp5_ASAP7_75t_SL g1291 ( .A(n_413), .B(n_1292), .Y(n_1291) );
CKINVDCx8_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
INVx5_ASAP7_75t_L g674 ( .A(n_414), .Y(n_674) );
NOR2xp33_ASAP7_75t_SL g1216 ( .A(n_414), .B(n_1217), .Y(n_1216) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_416), .Y(n_550) );
INVx2_ASAP7_75t_L g562 ( .A(n_416), .Y(n_562) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_416), .Y(n_640) );
INVx1_ASAP7_75t_L g901 ( .A(n_416), .Y(n_901) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g1746 ( .A(n_419), .Y(n_1746) );
INVx1_ASAP7_75t_L g724 ( .A(n_420), .Y(n_724) );
INVx2_ASAP7_75t_L g740 ( .A(n_420), .Y(n_740) );
BUFx2_ASAP7_75t_L g882 ( .A(n_420), .Y(n_882) );
INVx1_ASAP7_75t_L g1267 ( .A(n_420), .Y(n_1267) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AND2x2_ASAP7_75t_L g726 ( .A(n_421), .B(n_422), .Y(n_726) );
INVx4_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_SL g1358 ( .A1(n_424), .A2(n_606), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
AOI22xp5_ASAP7_75t_SL g1686 ( .A1(n_424), .A2(n_665), .B1(n_1687), .B2(n_1688), .Y(n_1686) );
BUFx2_ASAP7_75t_L g514 ( .A(n_425), .Y(n_514) );
INVx2_ASAP7_75t_L g528 ( .A(n_425), .Y(n_528) );
INVx6_ASAP7_75t_L g560 ( .A(n_425), .Y(n_560) );
OAI21xp5_ASAP7_75t_SL g573 ( .A1(n_426), .A2(n_574), .B(n_583), .Y(n_573) );
OAI31xp33_ASAP7_75t_L g831 ( .A1(n_426), .A2(n_832), .A3(n_833), .B(n_839), .Y(n_831) );
OAI31xp33_ASAP7_75t_SL g1149 ( .A1(n_426), .A2(n_1150), .A3(n_1151), .B(n_1156), .Y(n_1149) );
OAI31xp33_ASAP7_75t_L g1288 ( .A1(n_426), .A2(n_1289), .A3(n_1290), .B(n_1291), .Y(n_1288) );
AOI211xp5_ASAP7_75t_L g1356 ( .A1(n_426), .A2(n_1357), .B(n_1369), .C(n_1378), .Y(n_1356) );
OAI31xp33_ASAP7_75t_L g1400 ( .A1(n_426), .A2(n_1401), .A3(n_1402), .B(n_1403), .Y(n_1400) );
AOI211xp5_ASAP7_75t_L g1684 ( .A1(n_426), .A2(n_1685), .B(n_1696), .C(n_1705), .Y(n_1684) );
OAI31xp33_ASAP7_75t_SL g1741 ( .A1(n_426), .A2(n_1742), .A3(n_1743), .B(n_1744), .Y(n_1741) );
AND2x4_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
AND2x4_ASAP7_75t_L g613 ( .A(n_427), .B(n_429), .Y(n_613) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g531 ( .A(n_428), .B(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g494 ( .A(n_430), .Y(n_494) );
OR2x6_ASAP7_75t_L g905 ( .A(n_430), .B(n_906), .Y(n_905) );
OAI31xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_447), .A3(n_469), .B(n_471), .Y(n_431) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_438), .Y(n_433) );
AOI322xp5_ASAP7_75t_L g1737 ( .A1(n_434), .A2(n_463), .A3(n_541), .B1(n_597), .B2(n_1738), .C1(n_1739), .C2(n_1740), .Y(n_1737) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g442 ( .A(n_435), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g591 ( .A(n_435), .B(n_479), .Y(n_591) );
AND2x4_ASAP7_75t_L g768 ( .A(n_435), .B(n_443), .Y(n_768) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
INVx2_ASAP7_75t_L g1770 ( .A(n_438), .Y(n_1770) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g911 ( .A(n_439), .Y(n_911) );
INVx1_ASAP7_75t_L g925 ( .A(n_439), .Y(n_925) );
AND2x4_ASAP7_75t_L g479 ( .A(n_440), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g696 ( .A(n_440), .Y(n_696) );
INVx5_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_442), .A2(n_590), .B1(n_591), .B2(n_592), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_442), .A2(n_591), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_442), .A2(n_591), .B1(n_1347), .B2(n_1348), .Y(n_1346) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_442), .A2(n_1088), .B1(n_1360), .B2(n_1377), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g1703 ( .A1(n_442), .A2(n_1088), .B1(n_1688), .B2(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g1385 ( .A(n_444), .Y(n_1385) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
INVx1_ASAP7_75t_L g630 ( .A(n_445), .Y(n_630) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_445), .Y(n_802) );
AND2x4_ASAP7_75t_L g458 ( .A(n_446), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g930 ( .A(n_449), .Y(n_930) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g568 ( .A(n_450), .Y(n_568) );
INVx3_ASAP7_75t_L g704 ( .A(n_450), .Y(n_704) );
INVx2_ASAP7_75t_L g1137 ( .A(n_450), .Y(n_1137) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_451), .B(n_452), .Y(n_938) );
INVx1_ASAP7_75t_L g467 ( .A(n_452), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g588 ( .A(n_453), .B(n_589), .C(n_593), .D(n_598), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g756 ( .A(n_453), .B(n_757), .C(n_760), .D(n_766), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_453), .B(n_869), .C(n_872), .Y(n_868) );
NAND4xp25_ASAP7_75t_L g1005 ( .A(n_453), .B(n_1006), .C(n_1009), .D(n_1013), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1427 ( .A(n_453), .B(n_1428), .C(n_1430), .Y(n_1427) );
CKINVDCx11_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g994 ( .A1(n_454), .A2(n_491), .B(n_995), .C(n_996), .Y(n_994) );
AOI211xp5_ASAP7_75t_L g1079 ( .A1(n_454), .A2(n_623), .B(n_1080), .C(n_1081), .Y(n_1079) );
AOI211xp5_ASAP7_75t_L g1180 ( .A1(n_454), .A2(n_1181), .B(n_1182), .C(n_1183), .Y(n_1180) );
NOR3xp33_ASAP7_75t_L g1226 ( .A(n_454), .B(n_1227), .C(n_1228), .Y(n_1226) );
AOI211xp5_ASAP7_75t_SL g1343 ( .A1(n_454), .A2(n_1030), .B(n_1344), .C(n_1345), .Y(n_1343) );
AOI211xp5_ASAP7_75t_L g1370 ( .A1(n_454), .A2(n_870), .B(n_1371), .C(n_1372), .Y(n_1370) );
AOI211xp5_ASAP7_75t_L g1697 ( .A1(n_454), .A2(n_1413), .B(n_1698), .C(n_1699), .Y(n_1697) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp67_ASAP7_75t_L g468 ( .A(n_456), .Y(n_468) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_457), .B(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g492 ( .A(n_458), .Y(n_492) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_458), .Y(n_505) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_458), .Y(n_624) );
BUFx3_ASAP7_75t_L g871 ( .A(n_458), .Y(n_871) );
INVx1_ASAP7_75t_L g1031 ( .A(n_458), .Y(n_1031) );
BUFx2_ASAP7_75t_L g1330 ( .A(n_458), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_461), .A2(n_465), .B1(n_1011), .B2(n_1012), .Y(n_1051) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_463), .A2(n_465), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_463), .A2(n_505), .B1(n_594), .B2(n_595), .C1(n_596), .C2(n_597), .Y(n_593) );
INVx2_ASAP7_75t_L g765 ( .A(n_463), .Y(n_765) );
AOI222xp33_ASAP7_75t_L g869 ( .A1(n_463), .A2(n_465), .B1(n_837), .B2(n_838), .C1(n_865), .C2(n_870), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_463), .A2(n_465), .B1(n_940), .B2(n_941), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_463), .A2(n_465), .B1(n_1154), .B2(n_1155), .Y(n_1160) );
INVx2_ASAP7_75t_L g1184 ( .A(n_463), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_463), .A2(n_465), .B1(n_1293), .B2(n_1294), .Y(n_1298) );
AOI222xp33_ASAP7_75t_L g1428 ( .A1(n_463), .A2(n_505), .B1(n_597), .B2(n_1405), .C1(n_1406), .C2(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g690 ( .A(n_464), .Y(n_690) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_465), .A2(n_623), .B1(n_761), .B2(n_762), .C1(n_763), .C2(n_764), .Y(n_760) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
AND2x4_ASAP7_75t_L g597 ( .A(n_466), .B(n_468), .Y(n_597) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g602 ( .A(n_470), .Y(n_602) );
INVx5_ASAP7_75t_L g1088 ( .A(n_470), .Y(n_1088) );
OAI31xp33_ASAP7_75t_SL g563 ( .A1(n_471), .A2(n_564), .A3(n_565), .B(n_572), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_471), .A2(n_588), .B1(n_603), .B2(n_613), .C(n_614), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_471), .A2(n_756), .B1(n_770), .B2(n_782), .C(n_784), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g867 ( .A1(n_471), .A2(n_868), .B(n_874), .Y(n_867) );
OAI31xp33_ASAP7_75t_SL g933 ( .A1(n_471), .A2(n_934), .A3(n_935), .B(n_942), .Y(n_933) );
AOI221x1_ASAP7_75t_L g1004 ( .A1(n_471), .A2(n_675), .B1(n_1005), .B2(n_1016), .C(n_1025), .Y(n_1004) );
OAI31xp33_ASAP7_75t_L g1047 ( .A1(n_471), .A2(n_1048), .A3(n_1049), .B(n_1052), .Y(n_1047) );
OAI31xp33_ASAP7_75t_SL g1157 ( .A1(n_471), .A2(n_1158), .A3(n_1159), .B(n_1161), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_471), .A2(n_613), .B1(n_1168), .B2(n_1179), .C(n_1190), .Y(n_1167) );
OAI31xp33_ASAP7_75t_SL g1295 ( .A1(n_471), .A2(n_1296), .A3(n_1297), .B(n_1299), .Y(n_1295) );
OAI21xp5_ASAP7_75t_L g1426 ( .A1(n_471), .A2(n_1427), .B(n_1433), .Y(n_1426) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
AOI31xp33_ASAP7_75t_SL g993 ( .A1(n_472), .A2(n_994), .A3(n_998), .B(n_1000), .Y(n_993) );
AOI31xp33_ASAP7_75t_L g1078 ( .A1(n_472), .A2(n_1079), .A3(n_1083), .B(n_1086), .Y(n_1078) );
AOI31xp33_ASAP7_75t_L g1342 ( .A1(n_472), .A2(n_1343), .A3(n_1346), .B(n_1349), .Y(n_1342) );
AND2x4_ASAP7_75t_L g530 ( .A(n_473), .B(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g657 ( .A(n_473), .B(n_531), .Y(n_657) );
AND4x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_496), .C(n_512), .D(n_525), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .C(n_493), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g617 ( .A(n_478), .Y(n_617) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_479), .Y(n_498) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
AND2x2_ASAP7_75t_L g679 ( .A(n_479), .B(n_680), .Y(n_679) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_479), .Y(n_789) );
BUFx2_ASAP7_75t_L g799 ( .A(n_479), .Y(n_799) );
BUFx2_ASAP7_75t_L g844 ( .A(n_479), .Y(n_844) );
INVx1_ASAP7_75t_L g1098 ( .A(n_479), .Y(n_1098) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g928 ( .A(n_482), .Y(n_928) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g619 ( .A(n_484), .Y(n_619) );
INVx1_ASAP7_75t_L g914 ( .A(n_484), .Y(n_914) );
INVx2_ASAP7_75t_L g1100 ( .A(n_484), .Y(n_1100) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_485), .Y(n_500) );
INVx3_ASAP7_75t_L g792 ( .A(n_485), .Y(n_792) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
INVx2_ASAP7_75t_L g1194 ( .A(n_488), .Y(n_1194) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g502 ( .A(n_489), .Y(n_502) );
AND2x4_ASAP7_75t_L g714 ( .A(n_489), .B(n_680), .Y(n_714) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g622 ( .A(n_490), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g1009 ( .A1(n_491), .A2(n_597), .B1(n_764), .B2(n_1010), .C1(n_1011), .C2(n_1012), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1181 ( .A(n_491), .Y(n_1181) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g712 ( .A(n_492), .B(n_683), .Y(n_712) );
INVx1_ASAP7_75t_L g1236 ( .A(n_492), .Y(n_1236) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_493), .B(n_537), .C(n_540), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g615 ( .A(n_493), .B(n_616), .C(n_620), .Y(n_615) );
INVx2_ASAP7_75t_L g796 ( .A(n_493), .Y(n_796) );
BUFx3_ASAP7_75t_L g850 ( .A(n_493), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g1027 ( .A(n_493), .B(n_1028), .C(n_1029), .Y(n_1027) );
NAND3xp33_ASAP7_75t_L g1090 ( .A(n_493), .B(n_1091), .C(n_1093), .Y(n_1090) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_493), .B(n_1196), .C(n_1199), .Y(n_1195) );
NAND3xp33_ASAP7_75t_L g1379 ( .A(n_493), .B(n_1380), .C(n_1381), .Y(n_1379) );
NAND3xp33_ASAP7_75t_L g1706 ( .A(n_493), .B(n_1707), .C(n_1708), .Y(n_1706) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OR2x2_ASAP7_75t_L g522 ( .A(n_494), .B(n_523), .Y(n_522) );
OR2x6_ASAP7_75t_L g646 ( .A(n_494), .B(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g720 ( .A(n_494), .Y(n_720) );
OR2x2_ASAP7_75t_L g858 ( .A(n_494), .B(n_647), .Y(n_858) );
AND2x4_ASAP7_75t_L g992 ( .A(n_494), .B(n_495), .Y(n_992) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_494), .B(n_707), .Y(n_1036) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .C(n_506), .Y(n_496) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g539 ( .A(n_500), .Y(n_539) );
INVx2_ASAP7_75t_L g544 ( .A(n_500), .Y(n_544) );
INVx3_ASAP7_75t_L g1034 ( .A(n_500), .Y(n_1034) );
INVx2_ASAP7_75t_SL g1774 ( .A(n_500), .Y(n_1774) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g1413 ( .A(n_504), .Y(n_1413) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_505), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_505), .Y(n_1242) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_506), .B(n_626), .C(n_631), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g797 ( .A(n_506), .B(n_798), .C(n_803), .Y(n_797) );
CKINVDCx8_ASAP7_75t_R g932 ( .A(n_506), .Y(n_932) );
NAND3xp33_ASAP7_75t_L g982 ( .A(n_506), .B(n_983), .C(n_985), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_506), .B(n_1096), .C(n_1101), .Y(n_1095) );
NAND3xp33_ASAP7_75t_L g1191 ( .A(n_506), .B(n_1192), .C(n_1193), .Y(n_1191) );
NAND3xp33_ASAP7_75t_L g1415 ( .A(n_506), .B(n_1416), .C(n_1417), .Y(n_1415) );
INVx5_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx6_ASAP7_75t_L g546 ( .A(n_507), .Y(n_546) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g707 ( .A(n_510), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .C(n_521), .Y(n_512) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g1153 ( .A(n_516), .Y(n_1153) );
INVx1_ASAP7_75t_L g1247 ( .A(n_516), .Y(n_1247) );
BUFx3_ASAP7_75t_L g654 ( .A(n_518), .Y(n_654) );
INVx2_ASAP7_75t_L g1334 ( .A(n_518), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g655 ( .A(n_520), .Y(n_655) );
INVx1_ASAP7_75t_L g1263 ( .A(n_520), .Y(n_1263) );
INVx1_ASAP7_75t_L g1341 ( .A(n_520), .Y(n_1341) );
NAND3xp33_ASAP7_75t_L g547 ( .A(n_521), .B(n_548), .C(n_551), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g1037 ( .A(n_521), .B(n_1038), .C(n_1039), .Y(n_1037) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_521), .B(n_1104), .C(n_1106), .Y(n_1103) );
NAND3xp33_ASAP7_75t_L g1202 ( .A(n_521), .B(n_1203), .C(n_1205), .Y(n_1202) );
NAND3xp33_ASAP7_75t_L g1387 ( .A(n_521), .B(n_1388), .C(n_1390), .Y(n_1387) );
NAND3xp33_ASAP7_75t_L g1712 ( .A(n_521), .B(n_1713), .C(n_1714), .Y(n_1712) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g1140 ( .A1(n_522), .A2(n_818), .B1(n_1141), .B2(n_1144), .Y(n_1140) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g647 ( .A(n_524), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .C(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g549 ( .A(n_528), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_530), .B(n_555), .C(n_558), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g1040 ( .A(n_530), .B(n_1041), .C(n_1044), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1107 ( .A(n_530), .B(n_1108), .C(n_1109), .Y(n_1107) );
NAND3xp33_ASAP7_75t_L g1207 ( .A(n_530), .B(n_1208), .C(n_1209), .Y(n_1207) );
INVx1_ASAP7_75t_L g1277 ( .A(n_530), .Y(n_1277) );
NAND3xp33_ASAP7_75t_L g1393 ( .A(n_530), .B(n_1394), .C(n_1395), .Y(n_1393) );
NAND3xp33_ASAP7_75t_L g1715 ( .A(n_530), .B(n_1716), .C(n_1717), .Y(n_1715) );
XOR2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_584), .Y(n_533) );
NAND3xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_563), .C(n_573), .Y(n_534) );
AND4x1_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .C(n_547), .D(n_554), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .C(n_546), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_546), .A2(n_843), .B1(n_850), .B2(n_851), .C(n_857), .Y(n_842) );
AOI33xp33_ASAP7_75t_L g1233 ( .A1(n_546), .A2(n_992), .A3(n_1234), .B1(n_1237), .B2(n_1240), .B3(n_1241), .Y(n_1233) );
AOI33xp33_ASAP7_75t_L g1320 ( .A1(n_546), .A2(n_992), .A3(n_1321), .B1(n_1323), .B2(n_1326), .B3(n_1327), .Y(n_1320) );
INVx2_ASAP7_75t_L g1781 ( .A(n_546), .Y(n_1781) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_550), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_550), .Y(n_1316) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g899 ( .A(n_556), .Y(n_899) );
INVx2_ASAP7_75t_L g1246 ( .A(n_556), .Y(n_1246) );
INVx1_ASAP7_75t_L g895 ( .A(n_557), .Y(n_895) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g607 ( .A(n_560), .Y(n_607) );
INVx2_ASAP7_75t_SL g638 ( .A(n_560), .Y(n_638) );
INVx2_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
INVx2_ASAP7_75t_L g809 ( .A(n_560), .Y(n_809) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_560), .Y(n_978) );
BUFx6f_ASAP7_75t_L g1043 ( .A(n_560), .Y(n_1043) );
INVx1_ASAP7_75t_L g1389 ( .A(n_560), .Y(n_1389) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g1105 ( .A(n_562), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1767 ( .A1(n_566), .A2(n_1124), .B1(n_1758), .B2(n_1759), .Y(n_1767) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x6_ASAP7_75t_L g709 ( .A(n_568), .B(n_692), .Y(n_709) );
INVx2_ASAP7_75t_L g1364 ( .A(n_578), .Y(n_1364) );
INVx1_ASAP7_75t_L g1695 ( .A(n_578), .Y(n_1695) );
OAI22xp33_ASAP7_75t_L g1484 ( .A1(n_584), .A2(n_1478), .B1(n_1481), .B2(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g750 ( .A(n_585), .Y(n_750) );
XNOR2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_660), .Y(n_585) );
INVx1_ASAP7_75t_L g659 ( .A(n_587), .Y(n_659) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_591), .A2(n_602), .B1(n_758), .B2(n_759), .Y(n_757) );
AOI22xp5_ASAP7_75t_SL g1000 ( .A1(n_591), .A2(n_768), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_591), .A2(n_768), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_591), .A2(n_768), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_591), .A2(n_768), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
AOI22xp33_ASAP7_75t_SL g1373 ( .A1(n_591), .A2(n_600), .B1(n_1374), .B2(n_1375), .Y(n_1373) );
AOI22xp33_ASAP7_75t_L g1700 ( .A1(n_591), .A2(n_600), .B1(n_1701), .B2(n_1702), .Y(n_1700) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_600), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_600), .A2(n_602), .B1(n_864), .B2(n_873), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_600), .A2(n_602), .B1(n_969), .B2(n_999), .Y(n_998) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_600), .A2(n_602), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_600), .A2(n_1072), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_600), .A2(n_1088), .B1(n_1173), .B2(n_1189), .Y(n_1188) );
AOI22xp33_ASAP7_75t_SL g1349 ( .A1(n_600), .A2(n_602), .B1(n_1312), .B2(n_1350), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1430 ( .A1(n_600), .A2(n_602), .B1(n_1431), .B2(n_1432), .Y(n_1430) );
AOI211xp5_ASAP7_75t_L g1733 ( .A1(n_600), .A2(n_1734), .B(n_1735), .C(n_1736), .Y(n_1733) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_613), .Y(n_675) );
INVx1_ASAP7_75t_L g783 ( .A(n_613), .Y(n_783) );
OAI31xp33_ASAP7_75t_SL g943 ( .A1(n_613), .A2(n_944), .A3(n_945), .B(n_946), .Y(n_943) );
OAI21xp5_ASAP7_75t_L g1214 ( .A1(n_613), .A2(n_1215), .B(n_1224), .Y(n_1214) );
NAND4xp25_ASAP7_75t_SL g614 ( .A(n_615), .B(n_625), .C(n_634), .D(n_648), .Y(n_614) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g1092 ( .A(n_619), .Y(n_1092) );
BUFx3_ASAP7_75t_L g794 ( .A(n_621), .Y(n_794) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g633 ( .A(n_622), .Y(n_633) );
INVx2_ASAP7_75t_SL g991 ( .A(n_622), .Y(n_991) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g805 ( .A(n_624), .Y(n_805) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g1239 ( .A(n_629), .Y(n_1239) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g685 ( .A(n_630), .Y(n_685) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_633), .B(n_717), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_641), .C(n_645), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g814 ( .A(n_644), .Y(n_814) );
INVx1_ASAP7_75t_L g1425 ( .A(n_644), .Y(n_1425) );
NAND3xp33_ASAP7_75t_L g975 ( .A(n_645), .B(n_976), .C(n_979), .Y(n_975) );
AOI33xp33_ASAP7_75t_L g1331 ( .A1(n_645), .A2(n_656), .A3(n_1332), .B1(n_1335), .B2(n_1337), .B3(n_1338), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g736 ( .A(n_646), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_646), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_646), .A2(n_818), .B1(n_880), .B2(n_892), .Y(n_879) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .C(n_656), .Y(n_648) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g1422 ( .A(n_656), .B(n_1423), .C(n_1424), .Y(n_1422) );
BUFx4f_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx4f_ASAP7_75t_L g748 ( .A(n_657), .Y(n_748) );
INVx4_ASAP7_75t_L g818 ( .A(n_657), .Y(n_818) );
AOI221x1_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_675), .B1(n_676), .B2(n_718), .C(n_721), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .C(n_670), .D(n_674), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_668), .A2(n_711), .B1(n_712), .B2(n_713), .C1(n_714), .C2(n_715), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g703 ( .A1(n_671), .A2(n_704), .B(n_705), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_674), .B(n_771), .C(n_774), .D(n_776), .Y(n_770) );
NAND4xp25_ASAP7_75t_L g1016 ( .A(n_674), .B(n_1017), .C(n_1020), .D(n_1023), .Y(n_1016) );
NAND4xp25_ASAP7_75t_SL g1067 ( .A(n_674), .B(n_1068), .C(n_1071), .D(n_1074), .Y(n_1067) );
NAND4xp25_ASAP7_75t_SL g1307 ( .A(n_674), .B(n_1308), .C(n_1311), .D(n_1314), .Y(n_1307) );
NAND4xp25_ASAP7_75t_L g1357 ( .A(n_674), .B(n_1358), .C(n_1361), .D(n_1366), .Y(n_1357) );
NAND4xp25_ASAP7_75t_L g1685 ( .A(n_674), .B(n_1686), .C(n_1689), .D(n_1692), .Y(n_1685) );
OAI31xp33_ASAP7_75t_L g1053 ( .A1(n_675), .A2(n_1054), .A3(n_1055), .B(n_1059), .Y(n_1053) );
AOI211xp5_ASAP7_75t_L g1066 ( .A1(n_675), .A2(n_1067), .B(n_1078), .C(n_1089), .Y(n_1066) );
AOI211xp5_ASAP7_75t_SL g1306 ( .A1(n_675), .A2(n_1307), .B(n_1319), .C(n_1342), .Y(n_1306) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_686), .C(n_710), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_681), .B2(n_682), .Y(n_677) );
INVx2_ASAP7_75t_L g684 ( .A(n_680), .Y(n_684) );
AND2x4_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g1198 ( .A(n_685), .Y(n_1198) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_702), .C(n_708), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x6_ASAP7_75t_L g695 ( .A(n_692), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g717 ( .A(n_692), .Y(n_717) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g722 ( .A1(n_700), .A2(n_723), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g846 ( .A1(n_704), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_846) );
OAI22xp33_ASAP7_75t_SL g852 ( .A1(n_704), .A2(n_853), .B1(n_854), .B2(n_856), .Y(n_852) );
INVx1_ASAP7_75t_L g920 ( .A(n_704), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g1285 ( .A1(n_704), .A2(n_917), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI221xp5_ASAP7_75t_SL g737 ( .A1(n_711), .A2(n_713), .B1(n_738), .B2(n_741), .C(n_744), .Y(n_737) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx8_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_735), .B1(n_737), .B2(n_747), .Y(n_721) );
BUFx2_ASAP7_75t_L g893 ( .A(n_723), .Y(n_893) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
BUFx3_ASAP7_75t_L g861 ( .A(n_725), .Y(n_861) );
INVx1_ASAP7_75t_L g948 ( .A(n_725), .Y(n_948) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g743 ( .A(n_726), .Y(n_743) );
INVx1_ASAP7_75t_L g885 ( .A(n_726), .Y(n_885) );
INVx1_ASAP7_75t_L g1057 ( .A(n_726), .Y(n_1057) );
BUFx4f_ASAP7_75t_L g1270 ( .A(n_726), .Y(n_1270) );
BUFx4f_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g1261 ( .A(n_730), .Y(n_1261) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g1111 ( .A(n_732), .Y(n_1111) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g1756 ( .A(n_734), .Y(n_1756) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI33xp33_ASAP7_75t_L g1243 ( .A1(n_736), .A2(n_748), .A3(n_1244), .B1(n_1248), .B2(n_1250), .B3(n_1252), .Y(n_1243) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g860 ( .A(n_740), .Y(n_860) );
INVx2_ASAP7_75t_L g1142 ( .A(n_740), .Y(n_1142) );
INVx2_ASAP7_75t_L g1145 ( .A(n_740), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_742), .A2(n_1145), .B1(n_1146), .B2(n_1147), .C(n_1148), .Y(n_1144) );
INVx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g1763 ( .A1(n_746), .A2(n_1392), .B1(n_1764), .B2(n_1765), .Y(n_1763) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g972 ( .A(n_748), .B(n_973), .C(n_974), .Y(n_972) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
XNOR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_828), .Y(n_752) );
XNOR2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
BUFx4f_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI31xp33_ASAP7_75t_L g959 ( .A1(n_783), .A2(n_960), .A3(n_963), .B(n_968), .Y(n_959) );
NAND4xp25_ASAP7_75t_L g784 ( .A(n_785), .B(n_797), .C(n_806), .D(n_816), .Y(n_784) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_793), .C(n_795), .Y(n_785) );
INVx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx3_ASAP7_75t_L g984 ( .A(n_792), .Y(n_984) );
INVx2_ASAP7_75t_L g1133 ( .A(n_792), .Y(n_1133) );
INVx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVxp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
BUFx3_ASAP7_75t_L g845 ( .A(n_802), .Y(n_845) );
INVx2_ASAP7_75t_SL g1325 ( .A(n_802), .Y(n_1325) );
INVx4_ASAP7_75t_L g1411 ( .A(n_802), .Y(n_1411) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_SL g1322 ( .A(n_805), .Y(n_1322) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_810), .C(n_815), .Y(n_806) );
BUFx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1274 ( .A1(n_812), .A2(n_891), .B1(n_1275), .B2(n_1276), .Y(n_1274) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_SL g889 ( .A(n_813), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .C(n_824), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI22xp5_ASAP7_75t_SL g857 ( .A1(n_818), .A2(n_858), .B1(n_859), .B2(n_863), .Y(n_857) );
OAI33xp33_ASAP7_75t_L g1749 ( .A1(n_818), .A2(n_858), .A3(n_1750), .B1(n_1757), .B2(n_1761), .B3(n_1763), .Y(n_1749) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
BUFx2_ASAP7_75t_SL g965 ( .A(n_827), .Y(n_965) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND3x1_ASAP7_75t_SL g830 ( .A(n_831), .B(n_842), .C(n_867), .Y(n_830) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g1361 ( .A1(n_835), .A2(n_1362), .B(n_1363), .Y(n_1361) );
AOI21xp5_ASAP7_75t_L g1692 ( .A1(n_835), .A2(n_1693), .B(n_1694), .Y(n_1692) );
OAI221xp5_ASAP7_75t_L g859 ( .A1(n_847), .A2(n_849), .B1(n_860), .B2(n_861), .C(n_862), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g1135 ( .A1(n_848), .A2(n_1136), .B1(n_1137), .B2(n_1138), .Y(n_1135) );
INVx3_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI33xp33_ASAP7_75t_L g1258 ( .A1(n_858), .A2(n_1259), .A3(n_1264), .B1(n_1271), .B2(n_1274), .B3(n_1277), .Y(n_1258) );
INVx1_ASAP7_75t_SL g1421 ( .A(n_858), .Y(n_1421) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_860), .A2(n_861), .B1(n_864), .B2(n_865), .C(n_866), .Y(n_863) );
OAI22xp33_ASAP7_75t_SL g1757 ( .A1(n_860), .A2(n_1758), .B1(n_1759), .B2(n_1760), .Y(n_1757) );
OAI22xp33_ASAP7_75t_L g1761 ( .A1(n_860), .A2(n_861), .B1(n_1734), .B2(n_1762), .Y(n_1761) );
BUFx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g950 ( .A(n_875), .Y(n_950) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_933), .C(n_943), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_902), .Y(n_878) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_882), .B1(n_883), .B2(n_886), .C(n_887), .Y(n_880) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_881), .A2(n_886), .B1(n_917), .B2(n_919), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_883), .A2(n_1125), .B1(n_1126), .B2(n_1142), .C(n_1143), .Y(n_1141) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
BUFx2_ASAP7_75t_L g1760 ( .A(n_885), .Y(n_1760) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B1(n_895), .B2(n_896), .C(n_897), .Y(n_892) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI33xp33_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_907), .A3(n_916), .B1(n_921), .B2(n_927), .B3(n_932), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI33xp33_ASAP7_75t_L g1122 ( .A1(n_905), .A2(n_1123), .A3(n_1127), .B1(n_1131), .B2(n_1135), .B3(n_1139), .Y(n_1122) );
OAI33xp33_ASAP7_75t_L g1278 ( .A1(n_905), .A2(n_1139), .A3(n_1279), .B1(n_1280), .B2(n_1281), .B3(n_1285), .Y(n_1278) );
OAI33xp33_ASAP7_75t_L g1766 ( .A1(n_905), .A2(n_1767), .A3(n_1768), .B1(n_1771), .B2(n_1776), .B3(n_1781), .Y(n_1766) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_909), .B1(n_912), .B2(n_915), .Y(n_907) );
INVx2_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx2_ASAP7_75t_SL g1772 ( .A(n_910), .Y(n_1772) );
BUFx3_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
OAI22xp33_ASAP7_75t_SL g1127 ( .A1(n_914), .A2(n_1128), .B1(n_1129), .B2(n_1130), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g921 ( .A1(n_917), .A2(n_922), .B1(n_923), .B2(n_926), .Y(n_921) );
OAI22xp33_ASAP7_75t_L g1279 ( .A1(n_917), .A2(n_937), .B1(n_1265), .B2(n_1268), .Y(n_1279) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g1050 ( .A(n_920), .Y(n_1050) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
HB1xp67_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g1129 ( .A(n_925), .Y(n_1129) );
INVx1_ASAP7_75t_L g1282 ( .A(n_925), .Y(n_1282) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_927) );
BUFx3_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
OAI22xp33_ASAP7_75t_L g1123 ( .A1(n_937), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1123) );
INVx2_ASAP7_75t_L g1779 ( .A(n_937), .Y(n_1779) );
BUFx6f_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
XNOR2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_1162), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_1114), .B2(n_1117), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_1062), .B1(n_1063), .B2(n_1113), .Y(n_955) );
INVx1_ASAP7_75t_L g1113 ( .A(n_956), .Y(n_1113) );
OAI22x1_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_1003), .B1(n_1060), .B2(n_1061), .Y(n_956) );
INVx2_ASAP7_75t_L g1060 ( .A(n_957), .Y(n_1060) );
NOR3xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_971), .C(n_993), .Y(n_958) );
NAND4xp25_ASAP7_75t_L g971 ( .A(n_972), .B(n_975), .C(n_982), .D(n_986), .Y(n_971) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g1336 ( .A(n_978), .Y(n_1336) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND3xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .C(n_992), .Y(n_986) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_991), .Y(n_1102) );
INVx1_ASAP7_75t_L g1201 ( .A(n_991), .Y(n_1201) );
BUFx2_ASAP7_75t_L g1414 ( .A(n_992), .Y(n_1414) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1003), .Y(n_1061) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1006), .Y(n_1052) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1013), .Y(n_1048) );
INVxp67_ASAP7_75t_L g1054 ( .A(n_1017), .Y(n_1054) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_1023), .Y(n_1059) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_1026), .B(n_1047), .C(n_1053), .Y(n_1046) );
AND4x1_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1032), .C(n_1037), .D(n_1040), .Y(n_1026) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
NAND3xp33_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1035), .C(n_1036), .Y(n_1032) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1036), .Y(n_1139) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_1036), .B(n_1383), .C(n_1386), .Y(n_1382) );
NAND3xp33_ASAP7_75t_L g1709 ( .A(n_1036), .B(n_1710), .C(n_1711), .Y(n_1709) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1043), .Y(n_1204) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1043), .Y(n_1249) );
INVx4_ASAP7_75t_L g1251 ( .A(n_1043), .Y(n_1251) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1066), .Y(n_1112) );
NAND4xp25_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1095), .C(n_1103), .D(n_1107), .Y(n_1089) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1149), .C(n_1157), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1140), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1776 ( .A1(n_1124), .A2(n_1777), .B1(n_1778), .B2(n_1780), .Y(n_1776) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_1129), .A2(n_1132), .B1(n_1133), .B2(n_1134), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1280 ( .A1(n_1129), .A2(n_1133), .B1(n_1260), .B2(n_1262), .Y(n_1280) );
OAI22xp33_ASAP7_75t_L g1281 ( .A1(n_1133), .A2(n_1282), .B1(n_1283), .B2(n_1284), .Y(n_1281) );
XNOR2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1210), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
NAND3xp33_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1185), .C(n_1188), .Y(n_1179) );
NAND4xp25_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1195), .C(n_1202), .D(n_1207), .Y(n_1190) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1768 ( .A1(n_1198), .A2(n_1751), .B1(n_1754), .B2(n_1769), .Y(n_1768) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AOI22xp5_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1253), .B1(n_1300), .B2(n_1301), .Y(n_1210) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1211), .Y(n_1300) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
NAND4xp25_ASAP7_75t_L g1213 ( .A(n_1214), .B(n_1225), .C(n_1233), .D(n_1243), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1221), .Y(n_1215) );
AO21x1_ASAP7_75t_SL g1225 ( .A1(n_1226), .A2(n_1229), .B(n_1232), .Y(n_1225) );
AOI31xp33_ASAP7_75t_L g1369 ( .A1(n_1232), .A2(n_1370), .A3(n_1373), .B(n_1376), .Y(n_1369) );
AOI31xp33_ASAP7_75t_L g1696 ( .A1(n_1232), .A2(n_1697), .A3(n_1700), .B(n_1703), .Y(n_1696) );
OAI211xp5_ASAP7_75t_L g1732 ( .A1(n_1232), .A2(n_1733), .B(n_1741), .C(n_1748), .Y(n_1732) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1253), .Y(n_1301) );
INVx2_ASAP7_75t_SL g1253 ( .A(n_1254), .Y(n_1253) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
NAND3xp33_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1288), .C(n_1295), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1278), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_1260), .A2(n_1261), .B1(n_1262), .B2(n_1263), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1266), .B1(n_1268), .B2(n_1269), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_1266), .A2(n_1269), .B1(n_1272), .B2(n_1273), .Y(n_1271) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_1305), .A2(n_1351), .B1(n_1435), .B2(n_1436), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1435 ( .A(n_1305), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1331), .Y(n_1319) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_1334), .Y(n_1339) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1334), .Y(n_1753) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1351), .Y(n_1436) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1396), .B1(n_1397), .B2(n_1434), .Y(n_1351) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1352), .Y(n_1434) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
HB1xp67_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
XNOR2xp5_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1356), .Y(n_1354) );
NAND4xp25_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1382), .C(n_1387), .D(n_1393), .Y(n_1378) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
INVx2_ASAP7_75t_SL g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
NAND3x1_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1407), .C(n_1426), .Y(n_1399) );
AND4x1_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1415), .C(n_1418), .D(n_1422), .Y(n_1407) );
NAND3xp33_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1412), .C(n_1414), .Y(n_1408) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
NAND3xp33_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1420), .C(n_1421), .Y(n_1418) );
OAI221xp5_ASAP7_75t_SL g1437 ( .A1(n_1438), .A2(n_1679), .B1(n_1681), .B2(n_1718), .C(n_1723), .Y(n_1437) );
AND5x1_ASAP7_75t_L g1438 ( .A(n_1439), .B(n_1598), .C(n_1645), .D(n_1658), .E(n_1672), .Y(n_1438) );
OAI31xp33_ASAP7_75t_SL g1439 ( .A1(n_1440), .A2(n_1524), .A3(n_1559), .B(n_1588), .Y(n_1439) );
OAI322xp33_ASAP7_75t_L g1440 ( .A1(n_1441), .A2(n_1471), .A3(n_1488), .B1(n_1492), .B2(n_1498), .C1(n_1511), .C2(n_1513), .Y(n_1440) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
A2O1A1Ixp33_ASAP7_75t_L g1619 ( .A1(n_1442), .A2(n_1500), .B(n_1556), .C(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1463), .Y(n_1442) );
NOR2xp33_ASAP7_75t_L g1551 ( .A(n_1443), .B(n_1536), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1443), .B(n_1488), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1443), .B(n_1531), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1443), .B(n_1509), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1443), .B(n_1464), .Y(n_1671) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1443), .Y(n_1677) );
INVx4_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
INVx3_ASAP7_75t_L g1494 ( .A(n_1444), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1444), .B(n_1533), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1444), .B(n_1531), .Y(n_1568) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1444), .B(n_1539), .Y(n_1625) );
NOR3xp33_ASAP7_75t_L g1631 ( .A(n_1444), .B(n_1497), .C(n_1588), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1444), .B(n_1509), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1662 ( .A(n_1444), .B(n_1464), .Y(n_1662) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1444), .B(n_1486), .Y(n_1673) );
AND2x4_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1457), .Y(n_1444) );
AND2x4_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1452), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1479 ( .A(n_1448), .B(n_1453), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1451), .Y(n_1448) );
HB1xp67_ASAP7_75t_L g1787 ( .A(n_1449), .Y(n_1787) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1451), .Y(n_1460) );
AND2x4_ASAP7_75t_L g1454 ( .A(n_1452), .B(n_1455), .Y(n_1454) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1481 ( .A(n_1453), .B(n_1456), .Y(n_1481) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1458), .Y(n_1591) );
BUFx3_ASAP7_75t_L g1680 ( .A(n_1458), .Y(n_1680) );
AND2x4_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1461), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1459), .B(n_1461), .Y(n_1469) );
HB1xp67_ASAP7_75t_L g1788 ( .A(n_1459), .Y(n_1788) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
AND2x4_ASAP7_75t_L g1462 ( .A(n_1460), .B(n_1461), .Y(n_1462) );
INVx2_ASAP7_75t_L g1504 ( .A(n_1462), .Y(n_1504) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1463), .Y(n_1557) );
AOI22xp33_ASAP7_75t_L g1612 ( .A1(n_1463), .A2(n_1613), .B1(n_1615), .B2(n_1618), .Y(n_1612) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1463), .B(n_1501), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1467), .Y(n_1463) );
INVx1_ASAP7_75t_SL g1510 ( .A(n_1464), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g1518 ( .A(n_1464), .Y(n_1518) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1464), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1464), .B(n_1519), .Y(n_1555) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1464), .Y(n_1582) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1464), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1465), .B(n_1466), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1467), .B(n_1510), .Y(n_1509) );
CKINVDCx6p67_ASAP7_75t_R g1519 ( .A(n_1467), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1541 ( .A(n_1467), .B(n_1536), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g1577 ( .A(n_1467), .Y(n_1577) );
AOI221xp5_ASAP7_75t_L g1645 ( .A1(n_1467), .A2(n_1602), .B1(n_1646), .B2(n_1648), .C(n_1650), .Y(n_1645) );
OR2x6_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1470), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1486), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1473), .B(n_1489), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1473), .B(n_1488), .Y(n_1558) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1473), .B(n_1561), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1473), .B(n_1554), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1482), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1474), .B(n_1483), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1474), .B(n_1488), .Y(n_1548) );
INVx2_ASAP7_75t_L g1638 ( .A(n_1474), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1474), .B(n_1533), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1678 ( .A(n_1474), .B(n_1533), .Y(n_1678) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1475), .B(n_1483), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1475), .B(n_1482), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1476 ( .A1(n_1477), .A2(n_1478), .B1(n_1480), .B2(n_1481), .Y(n_1476) );
OAI22xp33_ASAP7_75t_L g1505 ( .A1(n_1478), .A2(n_1506), .B1(n_1507), .B2(n_1508), .Y(n_1505) );
BUFx3_ASAP7_75t_L g1594 ( .A(n_1478), .Y(n_1594) );
BUFx6f_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g1508 ( .A(n_1481), .Y(n_1508) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1481), .Y(n_1597) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1483), .Y(n_1497) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1487), .B(n_1489), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1487), .B(n_1532), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1487), .B(n_1488), .Y(n_1603) );
NOR2x1_ASAP7_75t_L g1496 ( .A(n_1488), .B(n_1497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1537 ( .A(n_1488), .B(n_1538), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1488), .B(n_1567), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1621 ( .A(n_1488), .B(n_1497), .Y(n_1621) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
BUFx3_ASAP7_75t_L g1533 ( .A(n_1489), .Y(n_1533) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1489), .B(n_1580), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1489), .B(n_1497), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1489), .B(n_1531), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1491), .Y(n_1489) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
NOR2xp33_ASAP7_75t_L g1493 ( .A(n_1494), .B(n_1495), .Y(n_1493) );
INVx2_ASAP7_75t_L g1516 ( .A(n_1494), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1494), .B(n_1539), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_1494), .B(n_1548), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1494), .B(n_1512), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1494), .B(n_1576), .Y(n_1575) );
OAI21xp5_ASAP7_75t_SL g1611 ( .A1(n_1494), .A2(n_1612), .B(n_1619), .Y(n_1611) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
OAI21xp33_ASAP7_75t_L g1549 ( .A1(n_1497), .A2(n_1550), .B(n_1552), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1497), .B(n_1533), .Y(n_1628) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1500), .B(n_1509), .Y(n_1499) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx2_ASAP7_75t_L g1523 ( .A(n_1501), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1501), .B(n_1589), .Y(n_1644) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVx2_ASAP7_75t_SL g1536 ( .A(n_1502), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1502), .B(n_1519), .Y(n_1545) );
OR2x2_ASAP7_75t_L g1587 ( .A(n_1502), .B(n_1522), .Y(n_1587) );
INVx2_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1510), .B(n_1545), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_1511), .B(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
NOR2xp33_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1520), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
NAND2xp5_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1517), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1516), .B(n_1603), .Y(n_1602) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_1516), .B(n_1628), .Y(n_1627) );
A2O1A1Ixp33_ASAP7_75t_L g1659 ( .A1(n_1516), .A2(n_1614), .B(n_1635), .C(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1517), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1519), .Y(n_1517) );
INVx3_ASAP7_75t_L g1522 ( .A(n_1518), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1518), .B(n_1535), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1518), .B(n_1602), .Y(n_1601) );
NOR2xp33_ASAP7_75t_L g1605 ( .A(n_1518), .B(n_1606), .Y(n_1605) );
OAI32xp33_ASAP7_75t_L g1654 ( .A1(n_1518), .A2(n_1586), .A3(n_1603), .B1(n_1609), .B2(n_1655), .Y(n_1654) );
AND2x4_ASAP7_75t_SL g1535 ( .A(n_1519), .B(n_1536), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1571 ( .A(n_1519), .B(n_1536), .Y(n_1571) );
NOR2xp33_ASAP7_75t_L g1615 ( .A(n_1519), .B(n_1616), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1519), .B(n_1617), .Y(n_1636) );
NAND3xp33_ASAP7_75t_L g1660 ( .A(n_1519), .B(n_1620), .C(n_1661), .Y(n_1660) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
OAI322xp33_ASAP7_75t_L g1665 ( .A1(n_1521), .A2(n_1534), .A3(n_1584), .B1(n_1587), .B2(n_1616), .C1(n_1666), .C2(n_1668), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1521 ( .A(n_1522), .B(n_1523), .Y(n_1521) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_1522), .B(n_1565), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1522), .B(n_1536), .Y(n_1647) );
OR2x2_ASAP7_75t_L g1649 ( .A(n_1522), .B(n_1530), .Y(n_1649) );
AOI21xp5_ASAP7_75t_L g1675 ( .A1(n_1522), .A2(n_1669), .B(n_1676), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1523), .B(n_1589), .Y(n_1657) );
OAI221xp5_ASAP7_75t_SL g1524 ( .A1(n_1525), .A2(n_1534), .B1(n_1537), .B2(n_1540), .C(n_1542), .Y(n_1524) );
INVxp67_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1529), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1532), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1531), .B(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1531), .Y(n_1580) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1532), .B(n_1539), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1533), .B(n_1609), .Y(n_1608) );
OR2x2_ASAP7_75t_L g1629 ( .A(n_1533), .B(n_1625), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1626 ( .A(n_1534), .B(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1581 ( .A(n_1541), .B(n_1582), .Y(n_1581) );
AOI21xp5_ASAP7_75t_L g1623 ( .A1(n_1541), .A2(n_1624), .B(n_1626), .Y(n_1623) );
AOI221xp5_ASAP7_75t_L g1542 ( .A1(n_1543), .A2(n_1546), .B1(n_1549), .B2(n_1555), .C(n_1556), .Y(n_1542) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1545), .Y(n_1610) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1555), .Y(n_1664) );
NOR2xp33_ASAP7_75t_L g1556 ( .A(n_1557), .B(n_1558), .Y(n_1556) );
NOR2xp33_ASAP7_75t_L g1663 ( .A(n_1558), .B(n_1664), .Y(n_1663) );
NAND4xp25_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1563), .C(n_1569), .D(n_1574), .Y(n_1559) );
O2A1O1Ixp33_ASAP7_75t_L g1672 ( .A1(n_1561), .A2(n_1566), .B(n_1673), .C(n_1674), .Y(n_1672) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1572), .Y(n_1569) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
AOI221xp5_ASAP7_75t_L g1574 ( .A1(n_1575), .A2(n_1577), .B1(n_1578), .B2(n_1581), .C(n_1583), .Y(n_1574) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1576), .Y(n_1606) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
AOI21xp33_ASAP7_75t_L g1583 ( .A1(n_1584), .A2(n_1585), .B(n_1587), .Y(n_1583) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
OAI221xp5_ASAP7_75t_SL g1622 ( .A1(n_1587), .A2(n_1616), .B1(n_1623), .B2(n_1629), .C(n_1630), .Y(n_1622) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
BUFx3_ASAP7_75t_L g1617 ( .A(n_1589), .Y(n_1617) );
O2A1O1Ixp33_ASAP7_75t_L g1658 ( .A1(n_1589), .A2(n_1659), .B(n_1663), .C(n_1665), .Y(n_1658) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
OAI22xp33_ASAP7_75t_L g1592 ( .A1(n_1593), .A2(n_1594), .B1(n_1595), .B2(n_1596), .Y(n_1592) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NOR5xp2_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1611), .C(n_1622), .D(n_1633), .E(n_1637), .Y(n_1598) );
AOI31xp33_ASAP7_75t_L g1599 ( .A1(n_1600), .A2(n_1604), .A3(n_1607), .B(n_1610), .Y(n_1599) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1603), .Y(n_1614) );
OAI21xp33_ASAP7_75t_L g1630 ( .A1(n_1603), .A2(n_1631), .B(n_1632), .Y(n_1630) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
AOI31xp33_ASAP7_75t_L g1633 ( .A1(n_1607), .A2(n_1634), .A3(n_1635), .B(n_1636), .Y(n_1633) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx2_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1632), .Y(n_1634) );
O2A1O1Ixp33_ASAP7_75t_L g1637 ( .A1(n_1638), .A2(n_1639), .B(n_1641), .C(n_1643), .Y(n_1637) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
OAI22xp5_ASAP7_75t_L g1674 ( .A1(n_1641), .A2(n_1643), .B1(n_1664), .B2(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
O2A1O1Ixp33_ASAP7_75t_SL g1650 ( .A1(n_1651), .A2(n_1653), .B(n_1654), .C(n_1657), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
NOR2xp33_ASAP7_75t_L g1669 ( .A(n_1652), .B(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVxp67_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1678), .Y(n_1676) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
HB1xp67_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
NAND4xp25_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1709), .C(n_1712), .D(n_1715), .Y(n_1705) );
CKINVDCx14_ASAP7_75t_R g1718 ( .A(n_1719), .Y(n_1718) );
INVx2_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
CKINVDCx5p33_ASAP7_75t_R g1720 ( .A(n_1721), .Y(n_1720) );
A2O1A1Ixp33_ASAP7_75t_L g1785 ( .A1(n_1722), .A2(n_1786), .B(n_1788), .C(n_1789), .Y(n_1785) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
HB1xp67_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1732), .Y(n_1782) );
OAI22xp5_ASAP7_75t_L g1771 ( .A1(n_1747), .A2(n_1772), .B1(n_1773), .B2(n_1775), .Y(n_1771) );
NOR2xp33_ASAP7_75t_L g1748 ( .A(n_1749), .B(n_1766), .Y(n_1748) );
OAI22xp5_ASAP7_75t_L g1750 ( .A1(n_1751), .A2(n_1752), .B1(n_1754), .B2(n_1755), .Y(n_1750) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
INVx2_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
INVx2_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
HB1xp67_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
endmodule