module fake_ariane_2081_n_1144 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_115, n_133, n_66, n_205, n_236, n_265, n_71, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_122, n_257, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1144);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_257;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1144;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_679;
wire n_643;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_1138;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_779;
wire n_731;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_557;
wire n_405;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_320;
wire n_559;
wire n_309;
wire n_331;
wire n_1134;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_721;
wire n_600;
wire n_433;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_839;
wire n_928;
wire n_821;
wire n_1099;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_677;
wire n_439;
wire n_604;
wire n_614;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_671;
wire n_303;
wire n_442;
wire n_777;
wire n_929;
wire n_538;
wire n_352;
wire n_899;
wire n_920;
wire n_1080;
wire n_576;
wire n_843;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_654;
wire n_455;
wire n_429;
wire n_365;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_1142;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_683;
wire n_601;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_708;
wire n_308;
wire n_551;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_626;
wire n_430;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_697;
wire n_274;
wire n_622;
wire n_437;
wire n_999;
wire n_998;
wire n_967;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_170),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_43),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_117),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_87),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_184),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_94),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_83),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_194),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_85),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_82),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_219),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_188),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_158),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_63),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_129),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_149),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_227),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_45),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_134),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_92),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_18),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_105),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_98),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_106),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_151),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_110),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_116),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_137),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_192),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_118),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_32),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_216),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_247),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_99),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_139),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_16),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_204),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_69),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_225),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_182),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_28),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_211),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_100),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_51),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_201),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_84),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_91),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_73),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_220),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_208),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_28),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_7),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_233),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_193),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_86),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_168),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_125),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_115),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_251),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_228),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_250),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_29),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_239),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_130),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_205),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_126),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_243),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_101),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_218),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_169),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_199),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_212),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_127),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_196),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_232),
.B(n_200),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_157),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_62),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_50),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_187),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_47),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_238),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_133),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_76),
.B(n_68),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_226),
.B(n_198),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_13),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_95),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_135),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_236),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_222),
.B(n_190),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_131),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_35),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_240),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_160),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_148),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_42),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_244),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_177),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_155),
.B(n_52),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_96),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_65),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_136),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_3),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_223),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_61),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_39),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_167),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_54),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_260),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_40),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_230),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_113),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_123),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_77),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_255),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_6),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_37),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_145),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_27),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_17),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_107),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_197),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_64),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_44),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_153),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_71),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_17),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_215),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_4),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_21),
.B(n_72),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_150),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_112),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_234),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_5),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_224),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_121),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_241),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_14),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_8),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_90),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_11),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_138),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_56),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_66),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_265),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_38),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_74),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_210),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_256),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_237),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_207),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_124),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_162),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_178),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_154),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_249),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_252),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_97),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_102),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_412),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_299),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_299),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_337),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_342),
.B(n_0),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_299),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_299),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_2),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_351),
.B(n_6),
.Y(n_453)
);

OAI22x1_ASAP7_75t_SL g454 ( 
.A1(n_323),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_454)
);

OA21x2_ASAP7_75t_L g455 ( 
.A1(n_266),
.A2(n_9),
.B(n_11),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_349),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_424),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_267),
.A2(n_159),
.B(n_261),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_290),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_280),
.A2(n_338),
.B1(n_341),
.B2(n_322),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_326),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_333),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_300),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_280),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_386),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_274),
.A2(n_152),
.B(n_259),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_334),
.Y(n_468)
);

CKINVDCx11_ASAP7_75t_R g469 ( 
.A(n_403),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_322),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_270),
.B(n_12),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_284),
.Y(n_472)
);

AND2x2_ASAP7_75t_SL g473 ( 
.A(n_348),
.B(n_15),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_410),
.Y(n_474)
);

OA21x2_ASAP7_75t_L g475 ( 
.A1(n_271),
.A2(n_15),
.B(n_16),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_272),
.B(n_18),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_338),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_275),
.B(n_30),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_378),
.B(n_284),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_345),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_369),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_304),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_319),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_273),
.B(n_19),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_334),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_319),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_347),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_347),
.Y(n_489)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_403),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_311),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_286),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_341),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_301),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_279),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_316),
.B(n_20),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_282),
.B(n_22),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_287),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_321),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_383),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_281),
.A2(n_166),
.B(n_258),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_294),
.A2(n_165),
.B(n_257),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_288),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_343),
.B(n_22),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_289),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_293),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_298),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_305),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_307),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_308),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_310),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_315),
.B(n_23),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_317),
.B(n_23),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

BUFx8_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_343),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_335),
.B(n_24),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_417),
.B(n_25),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_318),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_320),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_324),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_325),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_327),
.Y(n_528)
);

NOR2x1_ASAP7_75t_L g529 ( 
.A(n_328),
.B(n_31),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_268),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_329),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_330),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_336),
.B(n_26),
.Y(n_533)
);

BUFx8_ASAP7_75t_L g534 ( 
.A(n_440),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_344),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_346),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_350),
.B(n_27),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_361),
.B(n_29),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_355),
.A2(n_362),
.B(n_356),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_364),
.Y(n_540)
);

BUFx8_ASAP7_75t_L g541 ( 
.A(n_418),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_374),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_277),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_375),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_459),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_444),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_461),
.Y(n_548)
);

AO21x2_ASAP7_75t_L g549 ( 
.A1(n_471),
.A2(n_413),
.B(n_381),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_444),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_443),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

AO21x2_ASAP7_75t_L g554 ( 
.A1(n_471),
.A2(n_485),
.B(n_476),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_452),
.B(n_380),
.Y(n_555)
);

CKINVDCx6p67_ASAP7_75t_R g556 ( 
.A(n_469),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_476),
.B(n_358),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_464),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_543),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_487),
.B(n_379),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_487),
.B(n_384),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_445),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_472),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_486),
.B(n_358),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_506),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_448),
.B(n_276),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_446),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_456),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_530),
.B(n_385),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_457),
.B(n_306),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_450),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_506),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_450),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_470),
.A2(n_359),
.B1(n_373),
.B2(n_391),
.Y(n_578)
);

CKINVDCx6p67_ASAP7_75t_R g579 ( 
.A(n_469),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_511),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_511),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_452),
.B(n_380),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_453),
.B(n_420),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_451),
.Y(n_586)
);

AND3x2_ASAP7_75t_L g587 ( 
.A(n_507),
.B(n_382),
.C(n_434),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_453),
.B(n_387),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_466),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_494),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_466),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_493),
.B(n_388),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_520),
.B(n_414),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_501),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_493),
.B(n_389),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_492),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_465),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_492),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_502),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_484),
.B(n_406),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_479),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_502),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_512),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_507),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_538),
.B(n_435),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_539),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_496),
.B(n_394),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_457),
.B(n_398),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_479),
.A2(n_442),
.B1(n_414),
.B2(n_269),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_539),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_512),
.Y(n_618)
);

CKINVDCx6p67_ASAP7_75t_R g619 ( 
.A(n_490),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_442),
.Y(n_620)
);

AOI21x1_ASAP7_75t_L g621 ( 
.A1(n_529),
.A2(n_401),
.B(n_400),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_483),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_515),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_515),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_515),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_535),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_538),
.B(n_485),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_554),
.B(n_497),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_564),
.B(n_449),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_567),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_566),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_603),
.B(n_473),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_554),
.B(n_509),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_602),
.B(n_508),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_617),
.B(n_513),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_566),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_569),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_617),
.B(n_526),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_590),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_589),
.B(n_508),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_570),
.B(n_530),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_589),
.B(n_519),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_595),
.B(n_519),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_589),
.B(n_534),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_571),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_623),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_555),
.B(n_489),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_599),
.B(n_468),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_589),
.B(n_536),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_591),
.B(n_460),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_612),
.B(n_460),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_542),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_623),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_559),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_627),
.B(n_534),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_593),
.B(n_500),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_555),
.B(n_516),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_624),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_548),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_585),
.B(n_510),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_550),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_607),
.B(n_496),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_624),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_583),
.B(n_522),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_514),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_622),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_596),
.B(n_524),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_583),
.B(n_522),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_573),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_627),
.B(n_585),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_596),
.B(n_518),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_574),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_611),
.B(n_518),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_611),
.B(n_518),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_560),
.B(n_491),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_608),
.B(n_531),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_581),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_552),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_610),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_620),
.B(n_486),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_SL g684 ( 
.A(n_562),
.B(n_283),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_565),
.B(n_495),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_578),
.A2(n_470),
.B1(n_447),
.B2(n_520),
.C(n_454),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_615),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_619),
.B(n_527),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_558),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_610),
.B(n_525),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

BUFx8_ASAP7_75t_L g692 ( 
.A(n_556),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_549),
.B(n_528),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_579),
.Y(n_694)
);

AO221x1_ASAP7_75t_L g695 ( 
.A1(n_578),
.A2(n_447),
.B1(n_454),
.B2(n_477),
.C(n_540),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_549),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_SL g697 ( 
.A(n_608),
.B(n_516),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_587),
.A2(n_523),
.B1(n_521),
.B2(n_498),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_584),
.B(n_527),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_605),
.B(n_533),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_557),
.B(n_532),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_587),
.B(n_517),
.C(n_499),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_609),
.B(n_533),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_557),
.B(n_535),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_618),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_625),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_590),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_621),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_626),
.B(n_541),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_630),
.B(n_371),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_702),
.A2(n_499),
.B(n_517),
.C(n_537),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_660),
.A2(n_537),
.B(n_467),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_636),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_658),
.B(n_477),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_651),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_628),
.A2(n_504),
.B(n_458),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_648),
.B(n_541),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_628),
.A2(n_505),
.B(n_529),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_642),
.B(n_535),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_640),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_650),
.A2(n_478),
.B(n_427),
.C(n_411),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_683),
.B(n_578),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_698),
.B(n_544),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_633),
.A2(n_368),
.B(n_367),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_673),
.B(n_544),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_659),
.B(n_544),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_654),
.B(n_594),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_638),
.B(n_278),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_689),
.B(n_594),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_640),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_640),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_633),
.A2(n_368),
.B(n_367),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_662),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_663),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_674),
.A2(n_677),
.B(n_676),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_695),
.A2(n_594),
.B1(n_475),
.B2(n_455),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_659),
.B(n_540),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_668),
.A2(n_474),
.B(n_481),
.C(n_405),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_668),
.A2(n_478),
.B(n_475),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_687),
.B(n_463),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_649),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_670),
.B(n_285),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_670),
.B(n_291),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_708),
.A2(n_382),
.B(n_455),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_686),
.A2(n_426),
.B(n_407),
.C(n_409),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_664),
.A2(n_423),
.B1(n_430),
.B2(n_436),
.Y(n_746)
);

AOI33xp33_ASAP7_75t_L g747 ( 
.A1(n_681),
.A2(n_482),
.A3(n_463),
.B1(n_480),
.B2(n_439),
.B3(n_604),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_635),
.A2(n_639),
.B(n_701),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_632),
.A2(n_416),
.B1(n_295),
.B2(n_296),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_635),
.A2(n_547),
.B(n_545),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_639),
.A2(n_547),
.B(n_545),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_641),
.B(n_480),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_701),
.A2(n_703),
.B(n_700),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_708),
.A2(n_553),
.B(n_551),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_682),
.A2(n_553),
.B(n_551),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_667),
.A2(n_671),
.B(n_665),
.C(n_704),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_678),
.B(n_292),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_663),
.B(n_616),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_692),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_656),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_697),
.A2(n_397),
.B1(n_302),
.B2(n_303),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_690),
.A2(n_568),
.B(n_561),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_704),
.A2(n_568),
.B(n_561),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_637),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_691),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_693),
.A2(n_616),
.B1(n_614),
.B2(n_613),
.Y(n_767)
);

AOI21x1_ASAP7_75t_L g768 ( 
.A1(n_690),
.A2(n_575),
.B(n_572),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_652),
.A2(n_655),
.B(n_685),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_652),
.A2(n_575),
.B(n_572),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_669),
.B(n_297),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_655),
.A2(n_577),
.B(n_576),
.Y(n_772)
);

NAND2x1p5_ASAP7_75t_L g773 ( 
.A(n_657),
.B(n_576),
.Y(n_773)
);

BUFx12f_ASAP7_75t_L g774 ( 
.A(n_692),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_679),
.B(n_614),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_629),
.B(n_309),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_707),
.A2(n_580),
.B(n_577),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_706),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_693),
.A2(n_646),
.B(n_644),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_643),
.A2(n_586),
.B(n_580),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_679),
.B(n_586),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_SL g782 ( 
.A(n_694),
.B(n_312),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_684),
.B(n_313),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_647),
.A2(n_592),
.B(n_588),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_661),
.A2(n_592),
.B(n_588),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_716),
.A2(n_666),
.B(n_672),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_748),
.A2(n_680),
.B(n_675),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_724),
.A2(n_696),
.B1(n_634),
.B2(n_645),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_735),
.A2(n_705),
.B(n_331),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_737),
.B(n_709),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_732),
.A2(n_754),
.B(n_739),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_718),
.A2(n_598),
.B(n_597),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_712),
.A2(n_699),
.B(n_598),
.Y(n_793)
);

AO31x2_ASAP7_75t_L g794 ( 
.A1(n_779),
.A2(n_721),
.A3(n_711),
.B(n_763),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_745),
.A2(n_688),
.B(n_597),
.C(n_613),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_760),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_743),
.A2(n_392),
.B(n_332),
.Y(n_797)
);

AOI21x1_ASAP7_75t_L g798 ( 
.A1(n_768),
.A2(n_772),
.B(n_770),
.Y(n_798)
);

AOI21x1_ASAP7_75t_L g799 ( 
.A1(n_769),
.A2(n_606),
.B(n_604),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_714),
.A2(n_653),
.B1(n_390),
.B2(n_377),
.Y(n_800)
);

AND3x2_ASAP7_75t_L g801 ( 
.A(n_782),
.B(n_606),
.C(n_601),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_715),
.B(n_600),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_314),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_710),
.B(n_339),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_719),
.A2(n_393),
.B(n_352),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_726),
.A2(n_395),
.B(n_353),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_755),
.A2(n_396),
.B(n_354),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_717),
.A2(n_428),
.B(n_357),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_730),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_757),
.A2(n_601),
.B(n_600),
.C(n_419),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_713),
.A2(n_376),
.B1(n_441),
.B2(n_438),
.Y(n_811)
);

AO31x2_ASAP7_75t_L g812 ( 
.A1(n_750),
.A2(n_358),
.A3(n_590),
.B(n_36),
.Y(n_812)
);

O2A1O1Ixp5_ASAP7_75t_L g813 ( 
.A1(n_783),
.A2(n_358),
.B(n_437),
.C(n_433),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_740),
.B(n_733),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_744),
.A2(n_432),
.B(n_431),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_766),
.B(n_340),
.Y(n_816)
);

AOI21x1_ASAP7_75t_L g817 ( 
.A1(n_751),
.A2(n_358),
.B(n_590),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_776),
.A2(n_429),
.B(n_372),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_729),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_764),
.A2(n_358),
.B(n_34),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_756),
.A2(n_370),
.B(n_366),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_758),
.A2(n_365),
.B(n_363),
.Y(n_822)
);

O2A1O1Ixp5_ASAP7_75t_L g823 ( 
.A1(n_778),
.A2(n_360),
.B(n_46),
.C(n_48),
.Y(n_823)
);

AO22x2_ASAP7_75t_L g824 ( 
.A1(n_722),
.A2(n_33),
.B1(n_49),
.B2(n_53),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_734),
.B(n_55),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_727),
.B(n_57),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_741),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_771),
.A2(n_58),
.B(n_59),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_729),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_734),
.B(n_60),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_774),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_723),
.B(n_67),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_781),
.B(n_70),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_725),
.A2(n_75),
.B(n_78),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_730),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_762),
.A2(n_79),
.B(n_80),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_826),
.B(n_835),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_809),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_814),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_827),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_804),
.B(n_738),
.C(n_749),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_802),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_824),
.B(n_736),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_820),
.A2(n_785),
.B(n_777),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_809),
.Y(n_845)
);

HB1xp67_ASAP7_75t_SL g846 ( 
.A(n_819),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_829),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_831),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_836),
.A2(n_747),
.B(n_746),
.C(n_765),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_799),
.A2(n_784),
.B(n_780),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_835),
.B(n_759),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_809),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_798),
.A2(n_753),
.B(n_767),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_835),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_796),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_787),
.Y(n_856)
);

INVx6_ASAP7_75t_L g857 ( 
.A(n_830),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_791),
.A2(n_761),
.B(n_728),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_801),
.B(n_759),
.Y(n_859)
);

AO21x2_ASAP7_75t_L g860 ( 
.A1(n_810),
.A2(n_775),
.B(n_752),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_792),
.A2(n_720),
.B(n_765),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_786),
.A2(n_720),
.B(n_773),
.Y(n_862)
);

AOI22x1_ASAP7_75t_L g863 ( 
.A1(n_789),
.A2(n_731),
.B1(n_752),
.B2(n_775),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_795),
.B(n_731),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_815),
.A2(n_752),
.B(n_88),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_824),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_817),
.A2(n_81),
.B(n_89),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_800),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_794),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_794),
.Y(n_870)
);

AO21x2_ASAP7_75t_L g871 ( 
.A1(n_793),
.A2(n_93),
.B(n_103),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_869),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_851),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_851),
.B(n_833),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_869),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_870),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_840),
.Y(n_877)
);

AOI21x1_ASAP7_75t_L g878 ( 
.A1(n_856),
.A2(n_828),
.B(n_832),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_870),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_845),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_860),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_839),
.B(n_790),
.Y(n_882)
);

AOI21x1_ASAP7_75t_L g883 ( 
.A1(n_856),
.A2(n_807),
.B(n_803),
.Y(n_883)
);

INVx11_ASAP7_75t_L g884 ( 
.A(n_846),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_861),
.A2(n_823),
.B(n_834),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_861),
.A2(n_825),
.B(n_813),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_864),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_858),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_860),
.Y(n_889)
);

OAI22xp33_ASAP7_75t_L g890 ( 
.A1(n_868),
.A2(n_808),
.B1(n_788),
.B2(n_816),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_858),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_858),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_842),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_864),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_862),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_862),
.Y(n_896)
);

AOI21x1_ASAP7_75t_L g897 ( 
.A1(n_844),
.A2(n_806),
.B(n_805),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_837),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_860),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_838),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_847),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_844),
.A2(n_812),
.B(n_794),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_882),
.B(n_866),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_887),
.B(n_845),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_877),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_893),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_898),
.Y(n_907)
);

NAND2x1_ASAP7_75t_L g908 ( 
.A(n_887),
.B(n_894),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_882),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_901),
.B(n_838),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_898),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_887),
.B(n_845),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_898),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_876),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_872),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_876),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_900),
.B(n_848),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_900),
.B(n_851),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_872),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_873),
.B(n_855),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_894),
.B(n_845),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_873),
.B(n_855),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_890),
.B(n_843),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_879),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_874),
.A2(n_843),
.B1(n_841),
.B2(n_865),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_875),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_894),
.B(n_845),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_880),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_880),
.B(n_837),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_875),
.B(n_852),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_879),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_874),
.A2(n_857),
.B1(n_837),
.B2(n_818),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_888),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_881),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_881),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_880),
.B(n_852),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_874),
.B(n_854),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_926),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_910),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_926),
.B(n_889),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_924),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_909),
.B(n_857),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_915),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_908),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_906),
.B(n_889),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_919),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_905),
.B(n_899),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_931),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_924),
.B(n_899),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_914),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_920),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_904),
.B(n_895),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_903),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_904),
.B(n_902),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_904),
.B(n_902),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_934),
.B(n_892),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_923),
.B(n_857),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_914),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_934),
.B(n_892),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_916),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_912),
.B(n_895),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_916),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_912),
.B(n_896),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_912),
.B(n_896),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_922),
.B(n_857),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_918),
.B(n_852),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_933),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_917),
.B(n_852),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_933),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_921),
.B(n_888),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_930),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_935),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_928),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_927),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_954),
.B(n_935),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_971),
.B(n_921),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_954),
.B(n_921),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_955),
.B(n_936),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_953),
.B(n_925),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_939),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_971),
.B(n_891),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_955),
.B(n_929),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_938),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_956),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_973),
.B(n_925),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_939),
.B(n_891),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_941),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_951),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_943),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_940),
.B(n_928),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_951),
.B(n_932),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_974),
.B(n_937),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_952),
.B(n_907),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_961),
.B(n_937),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_961),
.B(n_812),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_968),
.B(n_884),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_963),
.B(n_812),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_974),
.B(n_907),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_963),
.B(n_883),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_964),
.B(n_883),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_940),
.B(n_911),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_941),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_943),
.B(n_911),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_946),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_964),
.B(n_871),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_978),
.B(n_972),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_1004),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_983),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_978),
.B(n_972),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_984),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1003),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_987),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_987),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1002),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1002),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_980),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_976),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_977),
.B(n_952),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_982),
.B(n_946),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_999),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_982),
.B(n_948),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_999),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_988),
.B(n_944),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_985),
.B(n_991),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_990),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1007),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1008),
.Y(n_1028)
);

OAI32xp33_ASAP7_75t_L g1029 ( 
.A1(n_1024),
.A2(n_985),
.A3(n_979),
.B1(n_1001),
.B2(n_998),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1012),
.B(n_975),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1009),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1011),
.B(n_975),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1011),
.B(n_948),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1021),
.B(n_1023),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_1017),
.A2(n_996),
.B(n_995),
.C(n_997),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_1017),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1026),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1013),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1025),
.A2(n_997),
.B1(n_995),
.B2(n_945),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1021),
.B(n_990),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1006),
.B(n_977),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1020),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1013),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1022),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1006),
.B(n_993),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_SL g1046 ( 
.A1(n_1036),
.A2(n_1023),
.B(n_1024),
.C(n_944),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_1033),
.B(n_1025),
.C(n_992),
.Y(n_1047)
);

OR2x2_ASAP7_75t_L g1048 ( 
.A(n_1032),
.B(n_1030),
.Y(n_1048)
);

OAI32xp33_ASAP7_75t_L g1049 ( 
.A1(n_1032),
.A2(n_1010),
.A3(n_1018),
.B1(n_1025),
.B2(n_966),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_1029),
.A2(n_1019),
.B(n_1005),
.C(n_957),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1035),
.A2(n_1039),
.B1(n_1044),
.B2(n_1042),
.Y(n_1051)
);

OAI211xp5_ASAP7_75t_SL g1052 ( 
.A1(n_1033),
.A2(n_944),
.B(n_965),
.C(n_797),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1031),
.B(n_1019),
.Y(n_1053)
);

OAI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_1037),
.A2(n_1019),
.B(n_1000),
.Y(n_1054)
);

INVxp33_ASAP7_75t_L g1055 ( 
.A(n_1045),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1027),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1041),
.A2(n_993),
.B1(n_973),
.B2(n_994),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1028),
.B(n_1000),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1040),
.B(n_884),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1038),
.A2(n_1005),
.B1(n_947),
.B2(n_945),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1034),
.B(n_993),
.Y(n_1061)
);

AOI322xp5_ASAP7_75t_L g1062 ( 
.A1(n_1034),
.A2(n_1015),
.A3(n_947),
.B1(n_849),
.B2(n_1016),
.C1(n_1014),
.C2(n_994),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1043),
.A2(n_959),
.B(n_956),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1056),
.B(n_1014),
.Y(n_1064)
);

AOI211xp5_ASAP7_75t_L g1065 ( 
.A1(n_1050),
.A2(n_942),
.B(n_811),
.C(n_849),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_1048),
.B(n_959),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1062),
.B(n_1063),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1059),
.B(n_973),
.Y(n_1068)
);

NAND3xp33_ASAP7_75t_L g1069 ( 
.A(n_1052),
.B(n_986),
.C(n_952),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1055),
.A2(n_986),
.B1(n_1016),
.B2(n_913),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_SL g1071 ( 
.A1(n_1051),
.A2(n_886),
.B(n_885),
.Y(n_1071)
);

AOI321xp33_ASAP7_75t_L g1072 ( 
.A1(n_1049),
.A2(n_970),
.A3(n_949),
.B1(n_960),
.B2(n_981),
.C(n_969),
.Y(n_1072)
);

AOI211x1_ASAP7_75t_L g1073 ( 
.A1(n_1047),
.A2(n_822),
.B(n_897),
.C(n_949),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_1053),
.B(n_913),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1054),
.A2(n_1060),
.B(n_1061),
.C(n_1058),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1046),
.B(n_897),
.C(n_854),
.Y(n_1076)
);

NAND3xp33_ASAP7_75t_L g1077 ( 
.A(n_1061),
.B(n_1057),
.C(n_913),
.Y(n_1077)
);

AOI211xp5_ASAP7_75t_L g1078 ( 
.A1(n_1050),
.A2(n_913),
.B(n_970),
.C(n_886),
.Y(n_1078)
);

CKINVDCx16_ASAP7_75t_R g1079 ( 
.A(n_1059),
.Y(n_1079)
);

OAI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1062),
.A2(n_854),
.B(n_863),
.C(n_885),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1050),
.A2(n_871),
.B(n_864),
.Y(n_1081)
);

AOI222xp33_ASAP7_75t_L g1082 ( 
.A1(n_1050),
.A2(n_960),
.B1(n_969),
.B2(n_962),
.C1(n_958),
.C2(n_950),
.Y(n_1082)
);

OAI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1050),
.A2(n_962),
.B1(n_958),
.B2(n_950),
.C(n_967),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1059),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1050),
.A2(n_871),
.B1(n_859),
.B2(n_852),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1067),
.A2(n_859),
.B(n_967),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_1073),
.B(n_821),
.C(n_859),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1078),
.A2(n_1080),
.B(n_1084),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_SL g1089 ( 
.A(n_1079),
.B(n_853),
.Y(n_1089)
);

NAND3x1_ASAP7_75t_L g1090 ( 
.A(n_1074),
.B(n_1076),
.C(n_1068),
.Y(n_1090)
);

NAND4xp25_ASAP7_75t_L g1091 ( 
.A(n_1077),
.B(n_104),
.C(n_108),
.D(n_109),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_1071),
.B(n_1069),
.C(n_1083),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1085),
.A2(n_853),
.B1(n_867),
.B2(n_850),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1066),
.B(n_867),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1064),
.B(n_878),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1070),
.Y(n_1096)
);

XNOR2x2_ASAP7_75t_L g1097 ( 
.A(n_1081),
.B(n_850),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1075),
.B(n_111),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1072),
.B(n_114),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_1098),
.B(n_1082),
.Y(n_1100)
);

NAND4xp75_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_1065),
.C(n_120),
.D(n_122),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1099),
.B(n_119),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1095),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1092),
.B(n_1096),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_L g1105 ( 
.A(n_1091),
.B(n_128),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_1087),
.B(n_878),
.C(n_140),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1094),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1089),
.B(n_262),
.C(n_141),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1086),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1097),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1093),
.B(n_132),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1090),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1095),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1095),
.Y(n_1114)
);

NOR2x1p5_ASAP7_75t_L g1115 ( 
.A(n_1104),
.B(n_147),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_1110),
.B(n_161),
.C(n_163),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_1107),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1112),
.B(n_164),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_SL g1119 ( 
.A(n_1101),
.B(n_171),
.C(n_172),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1109),
.B(n_173),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_L g1121 ( 
.A(n_1102),
.B(n_174),
.Y(n_1121)
);

AND3x1_ASAP7_75t_L g1122 ( 
.A(n_1100),
.B(n_175),
.C(n_176),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_L g1123 ( 
.A(n_1108),
.B(n_179),
.C(n_180),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1115),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1117),
.B(n_1114),
.Y(n_1125)
);

NOR2x1_ASAP7_75t_L g1126 ( 
.A(n_1116),
.B(n_1105),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_1120),
.B(n_1113),
.Y(n_1127)
);

XOR2xp5_ASAP7_75t_L g1128 ( 
.A(n_1122),
.B(n_1103),
.Y(n_1128)
);

NAND4xp75_ASAP7_75t_L g1129 ( 
.A(n_1121),
.B(n_1111),
.C(n_1106),
.D(n_185),
.Y(n_1129)
);

XNOR2xp5_ASAP7_75t_L g1130 ( 
.A(n_1119),
.B(n_181),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1127),
.B(n_1128),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1124),
.B(n_1118),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1125),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1126),
.A2(n_1123),
.B1(n_186),
.B2(n_189),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1130),
.Y(n_1135)
);

OA22x2_ASAP7_75t_L g1136 ( 
.A1(n_1135),
.A2(n_1131),
.B1(n_1132),
.B2(n_1133),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_1129),
.B1(n_191),
.B2(n_195),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1136),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1138),
.A2(n_1137),
.B(n_203),
.Y(n_1139)
);

AOI21xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1139),
.A2(n_202),
.B(n_206),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_SL g1141 ( 
.A(n_1140),
.B(n_213),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1141),
.A2(n_214),
.B(n_221),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1142),
.A2(n_229),
.B(n_235),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1143),
.A2(n_245),
.B(n_246),
.Y(n_1144)
);


endmodule