module fake_jpeg_12740_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_12),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_30),
.A2(n_22),
.B1(n_20),
.B2(n_16),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_13),
.B(n_10),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_36),
.B(n_22),
.C(n_16),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_39),
.Y(n_40)
);

AO22x2_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_21),
.B1(n_19),
.B2(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_36),
.B1(n_31),
.B2(n_33),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_13),
.C(n_10),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_38),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_35),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_44),
.B(n_42),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_9),
.C(n_44),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_48),
.B1(n_36),
.B2(n_46),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_36),
.B(n_1),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_0),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_0),
.C(n_2),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_3),
.Y(n_59)
);


endmodule