module real_aes_17167_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_855, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_855;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g845 ( .A(n_0), .B(n_846), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_1), .A2(n_3), .B1(n_132), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_2), .A2(n_47), .B1(n_139), .B2(n_245), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_4), .A2(n_28), .B1(n_210), .B2(n_245), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_5), .A2(n_18), .B1(n_129), .B2(n_178), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_6), .A2(n_105), .B1(n_839), .B2(n_852), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_7), .A2(n_64), .B1(n_157), .B2(n_212), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_8), .A2(n_20), .B1(n_139), .B2(n_161), .Y(n_555) );
INVx1_ASAP7_75t_L g846 ( .A(n_9), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_10), .A2(n_39), .B1(n_477), .B2(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_10), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_11), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_12), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g155 ( .A1(n_13), .A2(n_21), .B1(n_156), .B2(n_159), .Y(n_155) );
OR2x2_ASAP7_75t_L g475 ( .A(n_14), .B(n_44), .Y(n_475) );
BUFx2_ASAP7_75t_L g851 ( .A(n_14), .Y(n_851) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_15), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_16), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_17), .Y(n_830) );
OAI22xp5_ASAP7_75t_SL g110 ( .A1(n_19), .A2(n_76), .B1(n_111), .B2(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_22), .B(n_470), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_23), .A2(n_102), .B1(n_129), .B2(n_132), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_24), .A2(n_43), .B1(n_173), .B2(n_175), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_25), .B(n_130), .Y(n_223) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_26), .A2(n_60), .B(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_27), .A2(n_820), .B1(n_824), .B2(n_825), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_27), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_29), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_30), .Y(n_649) );
INVx4_ASAP7_75t_R g567 ( .A(n_31), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_32), .B(n_136), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_33), .A2(n_51), .B1(n_189), .B2(n_191), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_34), .A2(n_71), .B1(n_822), .B2(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_34), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_35), .A2(n_57), .B1(n_129), .B2(n_191), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_36), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_37), .B(n_173), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_38), .Y(n_236) );
INVx1_ASAP7_75t_L g477 ( .A(n_39), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_40), .B(n_245), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_SL g516 ( .A1(n_41), .A2(n_135), .B(n_139), .C(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_42), .A2(n_58), .B1(n_139), .B2(n_191), .Y(n_647) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_44), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_45), .A2(n_90), .B1(n_139), .B2(n_209), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_46), .A2(n_50), .B1(n_139), .B2(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_48), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_49), .A2(n_62), .B1(n_129), .B2(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g601 ( .A(n_52), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_53), .B(n_139), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_54), .Y(n_542) );
INVx2_ASAP7_75t_L g486 ( .A(n_55), .Y(n_486) );
INVx1_ASAP7_75t_L g473 ( .A(n_56), .Y(n_473) );
BUFx3_ASAP7_75t_L g494 ( .A(n_56), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_59), .A2(n_91), .B1(n_139), .B2(n_191), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_61), .Y(n_568) );
XNOR2xp5_ASAP7_75t_SL g820 ( .A(n_63), .B(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_65), .A2(n_79), .B1(n_138), .B2(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_66), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_67), .A2(n_81), .B1(n_139), .B2(n_161), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_68), .A2(n_101), .B1(n_129), .B2(n_159), .Y(n_233) );
AND2x4_ASAP7_75t_L g125 ( .A(n_69), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g148 ( .A(n_70), .Y(n_148) );
INVx1_ASAP7_75t_L g822 ( .A(n_71), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_72), .A2(n_93), .B1(n_189), .B2(n_191), .Y(n_576) );
AO22x1_ASAP7_75t_L g533 ( .A1(n_73), .A2(n_80), .B1(n_175), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g126 ( .A(n_74), .Y(n_126) );
AND2x2_ASAP7_75t_L g520 ( .A(n_75), .B(n_229), .Y(n_520) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_77), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_78), .B(n_212), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_82), .B(n_245), .Y(n_543) );
INVx2_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_84), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_85), .B(n_229), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_86), .A2(n_100), .B1(n_191), .B2(n_212), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_87), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_88), .B(n_146), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_89), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_92), .B(n_229), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_94), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_95), .B(n_229), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_96), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g500 ( .A(n_96), .Y(n_500) );
NAND2xp33_ASAP7_75t_L g226 ( .A(n_97), .B(n_130), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_98), .A2(n_163), .B(n_212), .C(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g569 ( .A(n_99), .B(n_570), .Y(n_569) );
NAND2xp33_ASAP7_75t_L g547 ( .A(n_103), .B(n_174), .Y(n_547) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_483), .B(n_487), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2x1_ASAP7_75t_L g107 ( .A(n_108), .B(n_480), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_468), .B(n_479), .Y(n_108) );
AOI21x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_113), .B(n_466), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_110), .Y(n_467) );
AOI211xp5_ASAP7_75t_SL g480 ( .A1(n_110), .A2(n_113), .B(n_466), .C(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g466 ( .A(n_114), .B(n_467), .Y(n_466) );
OAI22x1_ASAP7_75t_L g496 ( .A1(n_114), .A2(n_497), .B1(n_501), .B2(n_817), .Y(n_496) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_375), .Y(n_114) );
NOR2x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_314), .Y(n_115) );
NAND4xp25_ASAP7_75t_L g116 ( .A(n_117), .B(n_265), .C(n_284), .D(n_295), .Y(n_116) );
O2A1O1Ixp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_196), .B(n_203), .C(n_237), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_168), .Y(n_118) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_119), .B(n_330), .C(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g411 ( .A(n_119), .B(n_293), .Y(n_411) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_152), .Y(n_119) );
AND2x2_ASAP7_75t_L g255 ( .A(n_120), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g273 ( .A(n_120), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g290 ( .A(n_120), .Y(n_290) );
AND2x2_ASAP7_75t_L g335 ( .A(n_120), .B(n_170), .Y(n_335) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g200 ( .A(n_121), .Y(n_200) );
AND2x4_ASAP7_75t_L g283 ( .A(n_121), .B(n_274), .Y(n_283) );
AO31x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .A3(n_143), .B(n_149), .Y(n_121) );
AO31x2_ASAP7_75t_L g231 ( .A1(n_122), .A2(n_164), .A3(n_232), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_123), .A2(n_562), .B(n_565), .Y(n_561) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AO31x2_ASAP7_75t_L g153 ( .A1(n_124), .A2(n_154), .A3(n_164), .B(n_166), .Y(n_153) );
AO31x2_ASAP7_75t_L g170 ( .A1(n_124), .A2(n_171), .A3(n_180), .B(n_182), .Y(n_170) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_124), .A2(n_243), .A3(n_247), .B(n_248), .Y(n_242) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_124), .A2(n_151), .A3(n_554), .B(n_557), .Y(n_553) );
BUFx10_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g193 ( .A(n_125), .Y(n_193) );
INVx1_ASAP7_75t_L g519 ( .A(n_125), .Y(n_519) );
BUFx10_ASAP7_75t_L g551 ( .A(n_125), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B1(n_137), .B2(n_140), .Y(n_127) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_130), .Y(n_534) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g133 ( .A(n_131), .Y(n_133) );
INVx3_ASAP7_75t_L g139 ( .A(n_131), .Y(n_139) );
INVx1_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
INVx2_ASAP7_75t_L g210 ( .A(n_131), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_131), .Y(n_212) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_131), .Y(n_245) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_133), .B(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_134), .A2(n_155), .B1(n_160), .B2(n_162), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_134), .A2(n_140), .B1(n_172), .B2(n_177), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_134), .A2(n_140), .B1(n_188), .B2(n_190), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_134), .A2(n_208), .B1(n_211), .B2(n_213), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_134), .A2(n_225), .B(n_226), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_134), .A2(n_162), .B1(n_233), .B2(n_234), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_134), .A2(n_140), .B1(n_244), .B2(n_246), .Y(n_243) );
OAI22x1_ASAP7_75t_L g554 ( .A1(n_134), .A2(n_213), .B1(n_555), .B2(n_556), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_134), .A2(n_213), .B1(n_576), .B2(n_577), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_134), .A2(n_529), .B1(n_646), .B2(n_647), .Y(n_645) );
INVx6_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
O2A1O1Ixp5_ASAP7_75t_L g221 ( .A1(n_135), .A2(n_161), .B(n_222), .C(n_223), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_135), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_135), .A2(n_547), .B(n_548), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_135), .A2(n_528), .B(n_533), .C(n_536), .Y(n_587) );
BUFx8_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
INVx1_ASAP7_75t_L g515 ( .A(n_136), .Y(n_515) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
INVx4_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g529 ( .A(n_141), .Y(n_529) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g545 ( .A(n_142), .Y(n_545) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_143), .A2(n_187), .A3(n_192), .B(n_194), .Y(n_186) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_143), .A2(n_561), .B(n_569), .Y(n_560) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_SL g166 ( .A(n_145), .B(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_145), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g151 ( .A(n_146), .Y(n_151) );
INVx2_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_146), .A2(n_519), .B(n_531), .Y(n_536) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_151), .B(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g201 ( .A(n_152), .B(n_202), .Y(n_201) );
AND2x4_ASAP7_75t_L g258 ( .A(n_152), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_152), .Y(n_281) );
INVx1_ASAP7_75t_L g292 ( .A(n_152), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_152), .B(n_184), .Y(n_301) );
INVx2_ASAP7_75t_L g308 ( .A(n_152), .Y(n_308) );
INVx4_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g253 ( .A(n_153), .B(n_170), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_153), .B(n_260), .Y(n_326) );
AND2x2_ASAP7_75t_L g334 ( .A(n_153), .B(n_186), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_153), .B(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g387 ( .A(n_153), .Y(n_387) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_158), .B(n_564), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_161), .A2(n_542), .B(n_543), .C(n_544), .Y(n_541) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
AOI21x1_ASAP7_75t_L g507 ( .A1(n_164), .A2(n_508), .B(n_520), .Y(n_507) );
AO31x2_ASAP7_75t_L g574 ( .A1(n_164), .A2(n_192), .A3(n_575), .B(n_579), .Y(n_574) );
BUFx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_165), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g570 ( .A(n_165), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_165), .B(n_477), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_165), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g403 ( .A(n_169), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_184), .Y(n_169) );
INVx1_ASAP7_75t_L g202 ( .A(n_170), .Y(n_202) );
INVx1_ASAP7_75t_L g260 ( .A(n_170), .Y(n_260) );
INVx2_ASAP7_75t_L g294 ( .A(n_170), .Y(n_294) );
OR2x2_ASAP7_75t_L g298 ( .A(n_170), .B(n_186), .Y(n_298) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_170), .Y(n_347) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_174), .A2(n_179), .B1(n_567), .B2(n_568), .Y(n_566) );
OAI21xp33_ASAP7_75t_SL g597 ( .A1(n_175), .A2(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AO31x2_ASAP7_75t_L g206 ( .A1(n_180), .A2(n_192), .A3(n_207), .B(n_214), .Y(n_206) );
BUFx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_181), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_SL g219 ( .A(n_181), .Y(n_219) );
INVx4_ASAP7_75t_L g229 ( .A(n_181), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_181), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_181), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g605 ( .A(n_181), .B(n_551), .Y(n_605) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g320 ( .A(n_185), .B(n_200), .Y(n_320) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
INVx2_ASAP7_75t_L g274 ( .A(n_186), .Y(n_274) );
AND2x4_ASAP7_75t_L g293 ( .A(n_186), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g381 ( .A(n_186), .Y(n_381) );
INVx2_ASAP7_75t_L g578 ( .A(n_191), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_191), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_SL g227 ( .A(n_193), .Y(n_227) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_201), .Y(n_197) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g299 ( .A(n_199), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_199), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g362 ( .A(n_200), .Y(n_362) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2x1_ASAP7_75t_L g204 ( .A(n_205), .B(n_216), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_205), .B(n_217), .Y(n_312) );
INVx1_ASAP7_75t_L g410 ( .A(n_205), .Y(n_410) );
BUFx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g250 ( .A(n_206), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g264 ( .A(n_206), .B(n_242), .Y(n_264) );
AND2x4_ASAP7_75t_L g287 ( .A(n_206), .B(n_230), .Y(n_287) );
INVx2_ASAP7_75t_L g304 ( .A(n_206), .Y(n_304) );
AND2x2_ASAP7_75t_L g330 ( .A(n_206), .B(n_231), .Y(n_330) );
INVx1_ASAP7_75t_L g395 ( .A(n_206), .Y(n_395) );
INVx2_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_210), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_213), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g355 ( .A(n_216), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_230), .Y(n_216) );
AND2x2_ASAP7_75t_L g321 ( .A(n_217), .B(n_278), .Y(n_321) );
AND2x4_ASAP7_75t_L g337 ( .A(n_217), .B(n_304), .Y(n_337) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g331 ( .A(n_218), .Y(n_331) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_218) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_252) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_224), .B(n_227), .Y(n_220) );
INVx2_ASAP7_75t_L g247 ( .A(n_229), .Y(n_247) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_229), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
INVx3_ASAP7_75t_L g269 ( .A(n_230), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_230), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_230), .B(n_398), .Y(n_397) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g303 ( .A(n_231), .B(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g427 ( .A(n_231), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_253), .A3(n_254), .B1(n_255), .B2(n_257), .B3(n_261), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_250), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g361 ( .A(n_241), .B(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g270 ( .A(n_242), .B(n_252), .Y(n_270) );
INVx2_ASAP7_75t_L g278 ( .A(n_242), .Y(n_278) );
INVx1_ASAP7_75t_L g286 ( .A(n_242), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_245), .B(n_511), .Y(n_510) );
AO31x2_ASAP7_75t_L g644 ( .A1(n_247), .A2(n_551), .A3(n_645), .B(n_648), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_250), .A2(n_306), .B1(n_309), .B2(n_313), .Y(n_305) );
OR2x2_ASAP7_75t_L g445 ( .A(n_250), .B(n_263), .Y(n_445) );
AND2x4_ASAP7_75t_L g349 ( .A(n_251), .B(n_311), .Y(n_349) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_252), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_253), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_253), .B(n_289), .Y(n_391) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g364 ( .A(n_255), .Y(n_364) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g422 ( .A(n_258), .B(n_290), .Y(n_422) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_258), .B(n_289), .Y(n_440) );
AND2x2_ASAP7_75t_L g464 ( .A(n_258), .B(n_283), .Y(n_464) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g454 ( .A(n_262), .B(n_331), .Y(n_454) );
NOR2x1p5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g388 ( .A(n_263), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g356 ( .A(n_264), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_271), .B1(n_275), .B2(n_279), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g363 ( .A(n_268), .B(n_331), .Y(n_363) );
AND2x2_ASAP7_75t_L g400 ( .A(n_268), .B(n_349), .Y(n_400) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_269), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g441 ( .A(n_269), .B(n_270), .Y(n_441) );
AND2x2_ASAP7_75t_L g302 ( .A(n_270), .B(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g421 ( .A(n_270), .B(n_287), .Y(n_421) );
AND2x2_ASAP7_75t_L g465 ( .A(n_270), .B(n_330), .Y(n_465) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_275), .A2(n_400), .B1(n_401), .B2(n_404), .C1(n_406), .C2(n_407), .Y(n_399) );
AND2x2_ASAP7_75t_L g322 ( .A(n_276), .B(n_290), .Y(n_322) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g353 ( .A(n_277), .Y(n_353) );
INVxp67_ASAP7_75t_SL g398 ( .A(n_277), .Y(n_398) );
INVx2_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g368 ( .A(n_281), .Y(n_368) );
INVx2_ASAP7_75t_L g374 ( .A(n_282), .Y(n_374) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g358 ( .A(n_283), .B(n_347), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x4_ASAP7_75t_L g389 ( .A(n_286), .B(n_337), .Y(n_389) );
INVx2_ASAP7_75t_L g436 ( .A(n_286), .Y(n_436) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g379 ( .A(n_290), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g413 ( .A(n_290), .B(n_298), .Y(n_413) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_293), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g425 ( .A(n_293), .B(n_341), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B(n_302), .C(n_305), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OR2x2_ASAP7_75t_L g306 ( .A(n_298), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g342 ( .A(n_298), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_299), .B(n_334), .Y(n_438) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g414 ( .A(n_301), .B(n_383), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_303), .B(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_303), .A2(n_319), .B1(n_361), .B2(n_363), .Y(n_360) );
AND2x2_ASAP7_75t_L g366 ( .A(n_303), .B(n_331), .Y(n_366) );
AND2x2_ASAP7_75t_L g435 ( .A(n_303), .B(n_436), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_L g428 ( .A1(n_306), .A2(n_408), .B(n_429), .C(n_432), .Y(n_428) );
INVx2_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g419 ( .A(n_311), .Y(n_419) );
INVx1_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_313), .A2(n_360), .B1(n_364), .B2(n_365), .Y(n_359) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_327), .C(n_350), .Y(n_314) );
AO22x1_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B1(n_322), .B2(n_323), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_320), .Y(n_453) );
OR2x2_ASAP7_75t_L g460 ( .A(n_320), .B(n_341), .Y(n_460) );
AND2x2_ASAP7_75t_L g372 ( .A(n_321), .B(n_330), .Y(n_372) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g448 ( .A(n_326), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .C(n_338), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
AND2x4_ASAP7_75t_SL g406 ( .A(n_330), .B(n_349), .Y(n_406) );
INVx1_ASAP7_75t_SL g417 ( .A(n_330), .Y(n_417) );
OR2x2_ASAP7_75t_L g369 ( .A(n_331), .B(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_336), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x4_ASAP7_75t_L g346 ( .A(n_334), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g404 ( .A(n_335), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g426 ( .A(n_337), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g451 ( .A(n_337), .B(n_431), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_345), .B2(n_348), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x4_ASAP7_75t_L g386 ( .A(n_342), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g408 ( .A(n_342), .Y(n_408) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g463 ( .A(n_346), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_359), .C(n_367), .Y(n_350) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g432 ( .A(n_353), .Y(n_432) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_358), .A2(n_456), .B1(n_459), .B2(n_461), .C1(n_463), .C2(n_465), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_361), .B(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_371), .C(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_433), .Y(n_375) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_399), .C(n_409), .D(n_420), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_388), .B1(n_390), .B2(n_392), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .C(n_385), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_379), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_383), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g430 ( .A(n_395), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_397), .Y(n_462) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_412), .C(n_418), .Y(n_409) );
AOI21xp33_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_413), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_423), .B2(n_426), .C(n_428), .Y(n_420) );
INVx1_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
AOI31xp33_ASAP7_75t_L g442 ( .A1(n_424), .A2(n_443), .A3(n_444), .B(n_445), .Y(n_442) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_427), .Y(n_431) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_446), .C(n_455), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_439), .B2(n_441), .C(n_442), .Y(n_434) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g443 ( .A(n_441), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_449), .B1(n_452), .B2(n_454), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_476), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_470), .B(n_476), .Y(n_482) );
AND2x6_ASAP7_75t_SL g470 ( .A(n_471), .B(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_473), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_474), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_475), .B(n_494), .Y(n_838) );
OAI21xp33_ASAP7_75t_L g829 ( .A1(n_479), .A2(n_830), .B(n_831), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g491 ( .A(n_486), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_486), .B(n_836), .Y(n_835) );
OAI21x1_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_495), .B(n_828), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx6_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x6_ASAP7_75t_SL g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_819), .B1(n_826), .B2(n_827), .Y(n_495) );
INVx1_ASAP7_75t_L g826 ( .A(n_496), .Y(n_826) );
INVx4_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR3xp33_ASAP7_75t_L g843 ( .A(n_499), .B(n_844), .C(n_847), .Y(n_843) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g818 ( .A(n_500), .Y(n_818) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_717), .Y(n_502) );
NAND3xp33_ASAP7_75t_SL g503 ( .A(n_504), .B(n_620), .C(n_679), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_521), .B1(n_607), .B2(n_613), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g676 ( .A(n_506), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_506), .B(n_594), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_506), .B(n_640), .Y(n_787) );
AND2x2_ASAP7_75t_L g793 ( .A(n_506), .B(n_619), .Y(n_793) );
INVxp67_ASAP7_75t_L g798 ( .A(n_506), .Y(n_798) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g611 ( .A(n_507), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_516), .B(n_519), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B(n_514), .Y(n_509) );
BUFx4f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_515), .B(n_601), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_571), .B(n_580), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_552), .Y(n_523) );
INVx1_ASAP7_75t_L g714 ( .A(n_524), .Y(n_714) );
AND2x2_ASAP7_75t_L g743 ( .A(n_524), .B(n_705), .Y(n_743) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_537), .Y(n_524) );
AND2x2_ASAP7_75t_L g637 ( .A(n_525), .B(n_560), .Y(n_637) );
INVx1_ASAP7_75t_L g692 ( .A(n_525), .Y(n_692) );
AND2x2_ASAP7_75t_L g742 ( .A(n_525), .B(n_559), .Y(n_742) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g617 ( .A(n_526), .B(n_559), .Y(n_617) );
AND2x4_ASAP7_75t_L g761 ( .A(n_526), .B(n_560), .Y(n_761) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_532), .B(n_535), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI21x1_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_529), .A2(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g686 ( .A(n_537), .Y(n_686) );
AND2x2_ASAP7_75t_L g755 ( .A(n_537), .B(n_560), .Y(n_755) );
AND2x2_ASAP7_75t_L g762 ( .A(n_537), .B(n_588), .Y(n_762) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g584 ( .A(n_538), .Y(n_584) );
BUFx3_ASAP7_75t_L g619 ( .A(n_538), .Y(n_619) );
AND2x2_ASAP7_75t_L g630 ( .A(n_538), .B(n_616), .Y(n_630) );
AND2x2_ASAP7_75t_L g693 ( .A(n_538), .B(n_553), .Y(n_693) );
AND2x2_ASAP7_75t_L g698 ( .A(n_538), .B(n_560), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OAI21x1_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B(n_549), .Y(n_540) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_552), .B(n_704), .Y(n_806) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_559), .Y(n_552) );
INVx2_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
OR2x2_ASAP7_75t_L g591 ( .A(n_553), .B(n_560), .Y(n_591) );
INVx2_ASAP7_75t_L g616 ( .A(n_553), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_553), .B(n_586), .Y(n_632) );
AND2x2_ASAP7_75t_L g705 ( .A(n_553), .B(n_560), .Y(n_705) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g633 ( .A(n_560), .Y(n_633) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_572), .B(n_668), .Y(n_814) );
BUFx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g626 ( .A(n_573), .Y(n_626) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g606 ( .A(n_574), .Y(n_606) );
AND2x2_ASAP7_75t_L g612 ( .A(n_574), .B(n_594), .Y(n_612) );
INVx1_ASAP7_75t_L g660 ( .A(n_574), .Y(n_660) );
OR2x2_ASAP7_75t_L g665 ( .A(n_574), .B(n_644), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_574), .B(n_644), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_574), .B(n_643), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_574), .B(n_611), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_589), .B(n_592), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
OR2x2_ASAP7_75t_L g590 ( .A(n_583), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g741 ( .A(n_583), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g771 ( .A(n_583), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_584), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g739 ( .A(n_584), .Y(n_739) );
OR2x2_ASAP7_75t_L g652 ( .A(n_585), .B(n_653), .Y(n_652) );
INVxp33_ASAP7_75t_L g770 ( .A(n_585), .Y(n_770) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx2_ASAP7_75t_L g674 ( .A(n_586), .Y(n_674) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g628 ( .A(n_588), .Y(n_628) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g736 ( .A1(n_590), .A2(n_661), .B1(n_666), .B2(n_737), .C(n_740), .Y(n_736) );
OR2x2_ASAP7_75t_L g723 ( .A(n_591), .B(n_674), .Y(n_723) );
INVx2_ASAP7_75t_L g772 ( .A(n_591), .Y(n_772) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g672 ( .A(n_593), .Y(n_672) );
OR2x2_ASAP7_75t_L g675 ( .A(n_593), .B(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_593), .Y(n_716) );
OR2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_606), .Y(n_593) );
NAND2x1p5_ASAP7_75t_SL g625 ( .A(n_594), .B(n_610), .Y(n_625) );
INVx3_ASAP7_75t_L g640 ( .A(n_594), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_594), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_594), .Y(n_663) );
AND2x2_ASAP7_75t_L g744 ( .A(n_594), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g751 ( .A(n_594), .B(n_658), .Y(n_751) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_602), .B(n_605), .Y(n_596) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .Y(n_607) );
AND2x2_ASAP7_75t_L g803 ( .A(n_608), .B(n_662), .Y(n_803) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g707 ( .A(n_610), .B(n_677), .Y(n_707) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g642 ( .A(n_611), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g668 ( .A(n_611), .B(n_644), .Y(n_668) );
AND2x4_ASAP7_75t_L g765 ( .A(n_612), .B(n_735), .Y(n_765) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g684 ( .A(n_617), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_618), .B(n_705), .Y(n_789) );
AND2x2_ASAP7_75t_L g796 ( .A(n_618), .B(n_756), .Y(n_796) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g721 ( .A(n_619), .Y(n_721) );
AOI321xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_634), .A3(n_650), .B1(n_651), .B2(n_654), .C(n_669), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_622), .B(n_631), .Y(n_621) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_627), .B(n_629), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_624), .A2(n_635), .B(n_638), .Y(n_634) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
OR2x2_ASAP7_75t_L g733 ( .A(n_625), .B(n_665), .Y(n_733) );
INVx1_ASAP7_75t_L g725 ( .A(n_626), .Y(n_725) );
INVx2_ASAP7_75t_L g710 ( .A(n_627), .Y(n_710) );
OAI32xp33_ASAP7_75t_L g813 ( .A1(n_627), .A2(n_775), .A3(n_786), .B1(n_814), .B2(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g728 ( .A(n_628), .Y(n_728) );
INVx1_ASAP7_75t_L g678 ( .A(n_629), .Y(n_678) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_SL g766 ( .A(n_630), .B(n_673), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_631), .B(n_635), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_631), .A2(n_707), .B1(n_768), .B2(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g756 ( .A(n_632), .Y(n_756) );
INVx1_ASAP7_75t_L g653 ( .A(n_633), .Y(n_653) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g738 ( .A(n_637), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_638), .B(n_655), .C(n_661), .D(n_666), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVxp67_ASAP7_75t_L g680 ( .A(n_639), .Y(n_680) );
AND2x2_ASAP7_75t_L g759 ( .A(n_639), .B(n_668), .Y(n_759) );
OR2x2_ASAP7_75t_L g768 ( .A(n_639), .B(n_642), .Y(n_768) );
AND2x2_ASAP7_75t_L g792 ( .A(n_639), .B(n_664), .Y(n_792) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g706 ( .A(n_640), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g713 ( .A(n_640), .B(n_660), .Y(n_713) );
INVx1_ASAP7_75t_L g777 ( .A(n_641), .Y(n_777) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g685 ( .A(n_642), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g735 ( .A(n_642), .Y(n_735) );
INVx1_ASAP7_75t_L g677 ( .A(n_643), .Y(n_677) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g658 ( .A(n_644), .Y(n_658) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
AND2x4_ASAP7_75t_L g671 ( .A(n_657), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g712 ( .A(n_657), .Y(n_712) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_659), .Y(n_776) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x2_ASAP7_75t_L g667 ( .A(n_663), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g753 ( .A(n_665), .Y(n_753) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g730 ( .A(n_668), .Y(n_730) );
AND2x2_ASAP7_75t_L g773 ( .A(n_668), .B(n_713), .Y(n_773) );
O2A1O1Ixp33_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_673), .B(n_675), .C(n_678), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g784 ( .A(n_673), .B(n_762), .Y(n_784) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g688 ( .A(n_676), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B(n_694), .C(n_708), .Y(n_679) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B(n_687), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_683), .A2(n_791), .B(n_794), .Y(n_790) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g704 ( .A(n_686), .Y(n_704) );
AND2x2_ASAP7_75t_L g764 ( .A(n_686), .B(n_761), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g783 ( .A(n_691), .Y(n_783) );
AND2x2_ASAP7_75t_L g809 ( .A(n_691), .B(n_772), .Y(n_809) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g697 ( .A(n_692), .Y(n_697) );
INVx2_ASAP7_75t_L g748 ( .A(n_693), .Y(n_748) );
NAND2x1_ASAP7_75t_L g782 ( .A(n_693), .B(n_783), .Y(n_782) );
AOI33xp33_ASAP7_75t_L g800 ( .A1(n_693), .A2(n_713), .A3(n_751), .B1(n_761), .B2(n_793), .B3(n_855), .Y(n_800) );
OAI22xp33_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_699), .B1(n_702), .B2(n_706), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
AND2x2_ASAP7_75t_L g727 ( .A(n_698), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_699), .B(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
OR2x2_ASAP7_75t_L g812 ( .A(n_701), .B(n_746), .Y(n_812) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
OAI22xp33_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_711), .B1(n_714), .B2(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_712), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_712), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g734 ( .A(n_713), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g799 ( .A(n_713), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_778), .Y(n_717) );
NOR4xp25_ASAP7_75t_L g718 ( .A(n_719), .B(n_736), .C(n_757), .D(n_774), .Y(n_718) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_724), .B1(n_726), .B2(n_729), .C(n_731), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_SL g774 ( .A1(n_720), .A2(n_775), .B(n_776), .C(n_777), .Y(n_774) );
NAND2x1_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g807 ( .A(n_723), .Y(n_807) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_727), .A2(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OR2x6_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_743), .B(n_744), .C(n_747), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g786 ( .A(n_746), .B(n_787), .Y(n_786) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_746), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_752), .B2(n_754), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_763), .C(n_769), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_761), .A2(n_809), .B1(n_810), .B2(n_811), .C(n_813), .Y(n_808) );
INVx3_ASAP7_75t_L g816 ( .A(n_761), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_763) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g775 ( .A(n_772), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_801), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_790), .Y(n_779) );
O2A1O1Ixp33_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_784), .B(n_785), .C(n_788), .Y(n_780) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_784), .B(n_805), .C(n_807), .Y(n_804) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
OAI21xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_797), .B(n_800), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_804), .B(n_808), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g837 ( .A(n_818), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g827 ( .A(n_819), .Y(n_827) );
INVx1_ASAP7_75t_L g825 ( .A(n_820), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx10_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx3_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
BUFx12f_ASAP7_75t_L g853 ( .A(n_841), .Y(n_853) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g842 ( .A(n_843), .B(n_848), .Y(n_842) );
INVx2_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
NOR2x1p5_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx4f_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
endmodule