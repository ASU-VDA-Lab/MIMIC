module real_aes_7592_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_887;
wire n_599;
wire n_436;
wire n_1066;
wire n_684;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1205;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1170;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_635;
wire n_673;
wire n_518;
wire n_1192;
wire n_905;
wire n_878;
wire n_1067;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1110;
wire n_458;
wire n_1200;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_1123;
wire n_1034;
wire n_491;
wire n_923;
wire n_571;
wire n_694;
wire n_894;
wire n_952;
wire n_429;
wire n_1166;
wire n_1137;
wire n_448;
wire n_545;
wire n_556;
wire n_752;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_1021;
wire n_700;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1160;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_994;
wire n_578;
wire n_528;
wire n_495;
wire n_892;
wire n_1072;
wire n_1078;
wire n_938;
wire n_744;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_1199;
wire n_467;
wire n_875;
wire n_951;
wire n_992;
wire n_774;
wire n_813;
wire n_981;
wire n_791;
wire n_976;
wire n_466;
wire n_559;
wire n_872;
wire n_636;
wire n_1053;
wire n_1049;
wire n_477;
wire n_906;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1070;
wire n_726;
wire n_1189;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_1168;
wire n_746;
wire n_1025;
wire n_1148;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_725;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_1198;
wire n_782;
wire n_443;
wire n_565;
wire n_812;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_817;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_1196;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_1100;
wire n_1193;
wire n_1167;
wire n_1174;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_1149;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_1031;
wire n_432;
wire n_1037;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_1202;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_1179;
wire n_1201;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_1171;
wire n_1203;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1157;
wire n_1132;
wire n_853;
wire n_810;
wire n_1079;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1014;
wire n_1028;
wire n_1187;
wire n_1083;
wire n_727;
wire n_1056;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_1165;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1182;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_1204;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_831;
wire n_487;
wire n_899;
wire n_526;
wire n_928;
wire n_637;
wire n_653;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_1052;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_982;
wire n_717;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_1162;
wire n_861;
wire n_705;
wire n_1191;
wire n_1195;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_1175;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_1150;
wire n_1184;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_1045;
wire n_473;
wire n_566;
wire n_967;
wire n_719;
wire n_837;
wire n_871;
wire n_1159;
wire n_474;
wire n_1156;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_968;
wire n_743;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_1097;
wire n_661;
wire n_463;
wire n_1185;
wire n_804;
wire n_1076;
wire n_447;
wire n_1101;
wire n_1102;
wire n_1173;
wire n_603;
wire n_854;
wire n_403;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_1061;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_0), .A2(n_172), .B1(n_708), .B2(n_847), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_1), .B(n_671), .Y(n_793) );
XOR2x2_ASAP7_75t_L g809 ( .A(n_2), .B(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_3), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_4), .A2(n_299), .B1(n_771), .B2(n_911), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_5), .A2(n_165), .B1(n_530), .B2(n_821), .C(n_1056), .Y(n_1055) );
OA22x2_ASAP7_75t_L g894 ( .A1(n_6), .A2(n_895), .B1(n_896), .B2(n_916), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_6), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_7), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_8), .A2(n_89), .B1(n_593), .B2(n_914), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_9), .A2(n_358), .B1(n_583), .B2(n_595), .Y(n_1037) );
AOI22x1_ASAP7_75t_L g1172 ( .A1(n_10), .A2(n_1173), .B1(n_1198), .B2(n_1199), .Y(n_1172) );
INVx1_ASAP7_75t_L g1198 ( .A(n_10), .Y(n_1198) );
AOI22xp5_ASAP7_75t_SL g706 ( .A1(n_11), .A2(n_394), .B1(n_707), .B2(n_708), .Y(n_706) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_12), .A2(n_221), .B1(n_425), .B2(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g1145 ( .A(n_12), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_13), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g1106 ( .A1(n_14), .A2(n_204), .B1(n_814), .B2(n_885), .Y(n_1106) );
CKINVDCx20_ASAP7_75t_R g1196 ( .A(n_15), .Y(n_1196) );
AOI222xp33_ASAP7_75t_L g1169 ( .A1(n_16), .A2(n_58), .B1(n_330), .B2(n_567), .C1(n_680), .C2(n_1060), .Y(n_1169) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_17), .A2(n_301), .B1(n_551), .B2(n_789), .Y(n_788) );
AOI22xp5_ASAP7_75t_SL g701 ( .A1(n_18), .A2(n_248), .B1(n_541), .B2(n_702), .Y(n_701) );
AO22x1_ASAP7_75t_L g859 ( .A1(n_19), .A2(n_860), .B1(n_887), .B2(n_888), .Y(n_859) );
INVx1_ASAP7_75t_L g887 ( .A(n_19), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g997 ( .A(n_20), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_21), .A2(n_26), .B1(n_537), .B2(n_725), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_22), .A2(n_397), .B1(n_456), .B2(n_599), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_23), .A2(n_388), .B1(n_440), .B2(n_880), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g1094 ( .A(n_24), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_25), .A2(n_383), .B1(n_623), .B2(n_734), .Y(n_816) );
INVx1_ASAP7_75t_L g826 ( .A(n_27), .Y(n_826) );
AOI221xp5_ASAP7_75t_L g1164 ( .A1(n_28), .A2(n_251), .B1(n_821), .B2(n_1165), .C(n_1166), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_29), .A2(n_375), .B1(n_452), .B2(n_623), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_30), .A2(n_174), .B1(n_698), .B2(n_699), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_31), .A2(n_349), .B1(n_624), .B2(n_802), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_32), .A2(n_97), .B1(n_495), .B2(n_568), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_33), .A2(n_638), .B1(n_681), .B2(n_682), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_33), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g907 ( .A(n_34), .Y(n_907) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_35), .A2(n_106), .B1(n_425), .B2(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_36), .A2(n_259), .B1(n_732), .B2(n_738), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g1168 ( .A(n_37), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_38), .A2(n_278), .B1(n_446), .B2(n_1039), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_39), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_40), .A2(n_255), .B1(n_531), .B2(n_839), .Y(n_1075) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_41), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g1073 ( .A1(n_42), .A2(n_341), .B1(n_789), .B2(n_1074), .Y(n_1073) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_43), .A2(n_332), .B1(n_589), .B2(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_44), .A2(n_227), .B1(n_519), .B2(n_521), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g1070 ( .A(n_45), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_46), .A2(n_231), .B1(n_521), .B2(n_595), .Y(n_886) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_47), .A2(n_145), .B1(n_294), .B2(n_678), .C1(n_679), .C2(n_680), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_48), .B(n_573), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g1058 ( .A(n_49), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_50), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_51), .Y(n_1193) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_52), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_53), .A2(n_196), .B1(n_573), .B2(n_691), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_54), .B(n_825), .Y(n_932) );
AOI222xp33_ASAP7_75t_L g1059 ( .A1(n_55), .A2(n_212), .B1(n_323), .B2(n_691), .C1(n_722), .C2(n_1060), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_56), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_57), .A2(n_337), .B1(n_593), .B2(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_59), .A2(n_215), .B1(n_452), .B2(n_456), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g1160 ( .A(n_60), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_61), .A2(n_188), .B1(n_440), .B2(n_445), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_62), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_63), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_64), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_65), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_66), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_67), .A2(n_376), .B1(n_441), .B2(n_592), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_68), .A2(n_296), .B1(n_525), .B2(n_769), .Y(n_797) );
AOI22xp5_ASAP7_75t_SL g602 ( .A1(n_69), .A2(n_603), .B1(n_627), .B2(n_628), .Y(n_602) );
CKINVDCx16_ASAP7_75t_R g628 ( .A(n_69), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_70), .A2(n_205), .B1(n_418), .B2(n_598), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_71), .A2(n_126), .B1(n_465), .B2(n_911), .Y(n_1186) );
INVx1_ASAP7_75t_L g711 ( .A(n_72), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_73), .A2(n_102), .B1(n_465), .B2(n_882), .Y(n_881) );
AOI222xp33_ASAP7_75t_L g545 ( .A1(n_74), .A2(n_203), .B1(n_241), .B2(n_546), .C1(n_547), .C2(n_549), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_75), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_76), .Y(n_613) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_77), .A2(n_206), .B1(n_538), .B2(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g855 ( .A1(n_78), .A2(n_268), .B1(n_710), .B2(n_734), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_79), .A2(n_280), .B1(n_418), .B2(n_435), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g1078 ( .A1(n_80), .A2(n_81), .B1(n_654), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_82), .A2(n_144), .B1(n_525), .B2(n_620), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_83), .A2(n_235), .B1(n_519), .B2(n_938), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g1077 ( .A1(n_84), .A2(n_243), .B1(n_445), .B2(n_943), .Y(n_1077) );
AOI22xp5_ASAP7_75t_SL g703 ( .A1(n_85), .A2(n_253), .B1(n_626), .B2(n_704), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_86), .Y(n_1012) );
OA22x2_ASAP7_75t_L g1064 ( .A1(n_87), .A2(n_1065), .B1(n_1066), .B2(n_1085), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g1065 ( .A(n_87), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_88), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_90), .A2(n_128), .B1(n_543), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_91), .A2(n_308), .B1(n_456), .B2(n_523), .Y(n_1104) );
CKINVDCx20_ASAP7_75t_R g1189 ( .A(n_92), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_93), .A2(n_113), .B1(n_435), .B2(n_541), .Y(n_540) );
AO22x2_ASAP7_75t_L g434 ( .A1(n_94), .A2(n_258), .B1(n_425), .B2(n_426), .Y(n_434) );
INVx1_ASAP7_75t_L g1142 ( .A(n_94), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_95), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_96), .A2(n_183), .B1(n_537), .B2(n_994), .Y(n_993) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_98), .Y(n_657) );
AOI22xp5_ASAP7_75t_SL g709 ( .A1(n_99), .A2(n_210), .B1(n_418), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_100), .A2(n_297), .B1(n_543), .B2(n_544), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_101), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_103), .A2(n_414), .B1(n_510), .B2(n_511), .Y(n_413) );
INVx1_ASAP7_75t_L g510 ( .A(n_103), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_104), .A2(n_112), .B1(n_547), .B2(n_549), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_105), .A2(n_177), .B1(n_535), .B2(n_679), .Y(n_1120) );
INVx1_ASAP7_75t_L g1146 ( .A(n_106), .Y(n_1146) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_107), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_108), .B(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_109), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_110), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g1167 ( .A(n_111), .Y(n_1167) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_114), .A2(n_342), .B1(n_535), .B2(n_537), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_115), .A2(n_199), .B1(n_617), .B2(n_854), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_116), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_117), .A2(n_365), .B1(n_583), .B2(n_943), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g1184 ( .A(n_118), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_119), .A2(n_338), .B1(n_525), .B2(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_120), .Y(n_1190) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_121), .A2(n_209), .B1(n_842), .B2(n_843), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_122), .A2(n_372), .B1(n_598), .B2(n_738), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_123), .A2(n_244), .B1(n_418), .B2(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_124), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_125), .A2(n_271), .B1(n_769), .B2(n_1083), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_127), .A2(n_140), .B1(n_548), .B2(n_551), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g1053 ( .A(n_129), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_130), .A2(n_344), .B1(n_543), .B2(n_771), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_131), .A2(n_245), .B1(n_535), .B2(n_568), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_132), .A2(n_380), .B1(n_775), .B2(n_777), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_133), .A2(n_355), .B1(n_551), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_134), .A2(n_315), .B1(n_1039), .B2(n_1181), .Y(n_1180) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_135), .A2(n_153), .B1(n_643), .B2(n_938), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_136), .A2(n_190), .B1(n_531), .B2(n_669), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_137), .A2(n_373), .B1(n_595), .B2(n_598), .Y(n_594) );
XNOR2x2_ASAP7_75t_L g1030 ( .A(n_138), .B(n_1031), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_139), .A2(n_151), .B1(n_519), .B2(n_643), .Y(n_985) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_141), .A2(n_214), .B1(n_738), .B2(n_1151), .C(n_1153), .Y(n_1150) );
INVx1_ASAP7_75t_L g803 ( .A(n_142), .Y(n_803) );
AND2x6_ASAP7_75t_L g403 ( .A(n_143), .B(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_143), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_146), .A2(n_382), .B1(n_456), .B2(n_707), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_147), .A2(n_187), .B1(n_617), .B2(n_735), .Y(n_1028) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_148), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g840 ( .A(n_149), .B(n_530), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_150), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g942 ( .A1(n_152), .A2(n_360), .B1(n_734), .B2(n_943), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_154), .A2(n_192), .B1(n_446), .B2(n_620), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_155), .B(n_839), .Y(n_838) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_156), .A2(n_267), .B1(n_721), .B2(n_722), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_157), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_158), .Y(n_641) );
AO22x1_ASAP7_75t_L g1044 ( .A1(n_159), .A2(n_1045), .B1(n_1061), .B2(n_1062), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g1061 ( .A(n_159), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g1122 ( .A1(n_160), .A2(n_178), .B1(n_735), .B2(n_1123), .Y(n_1122) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_161), .A2(n_399), .B(n_408), .C(n_1147), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_162), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_163), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g1043 ( .A1(n_164), .A2(n_207), .B1(n_350), .B2(n_680), .C1(n_721), .C2(n_825), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_166), .A2(n_306), .B1(n_519), .B2(n_885), .Y(n_884) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_167), .A2(n_252), .B1(n_425), .B2(n_429), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g1143 ( .A(n_167), .B(n_1144), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_168), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g1194 ( .A(n_169), .Y(n_1194) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_170), .A2(n_198), .B1(n_620), .B2(n_1034), .C(n_1159), .Y(n_1158) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_171), .A2(n_181), .B1(n_583), .B2(n_584), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g967 ( .A(n_173), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_175), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_176), .A2(n_202), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_179), .A2(n_260), .B1(n_441), .B2(n_543), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_180), .A2(n_189), .B1(n_669), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_182), .A2(n_331), .B1(n_586), .B2(n_589), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_184), .A2(n_322), .B1(n_440), .B2(n_598), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_185), .A2(n_201), .B1(n_623), .B2(n_1034), .C(n_1047), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_186), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_191), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_193), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g902 ( .A(n_194), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_195), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_197), .A2(n_303), .B1(n_544), .B2(n_644), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_200), .A2(n_300), .B1(n_461), .B2(n_771), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g1179 ( .A(n_208), .Y(n_1179) );
AOI22xp33_ASAP7_75t_SL g937 ( .A1(n_211), .A2(n_242), .B1(n_541), .B2(n_938), .Y(n_937) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_213), .A2(n_234), .B1(n_462), .B2(n_626), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_216), .A2(n_239), .B1(n_456), .B2(n_619), .C(n_1051), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_217), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_218), .A2(n_345), .B1(n_589), .B2(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_219), .A2(n_352), .B1(n_461), .B2(n_465), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_220), .A2(n_240), .B1(n_456), .B2(n_644), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_222), .B(n_530), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_223), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_224), .A2(n_364), .B1(n_486), .B2(n_551), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_225), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_226), .A2(n_273), .B1(n_486), .B2(n_904), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g1025 ( .A1(n_228), .A2(n_310), .B1(n_771), .B2(n_882), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_229), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_230), .A2(n_371), .B1(n_619), .B2(n_620), .Y(n_618) );
OA22x2_ASAP7_75t_L g922 ( .A1(n_232), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_232), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g1049 ( .A(n_233), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_236), .A2(n_254), .B1(n_523), .B2(n_525), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_237), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_238), .A2(n_334), .B1(n_521), .B2(n_1034), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_246), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_247), .Y(n_689) );
INVx2_ASAP7_75t_L g407 ( .A(n_249), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_250), .A2(n_295), .B1(n_525), .B2(n_802), .Y(n_1111) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_256), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_257), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_261), .A2(n_976), .B1(n_1000), .B2(n_1001), .Y(n_975) );
INVx1_ASAP7_75t_L g1000 ( .A(n_261), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_262), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_263), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g1093 ( .A(n_264), .Y(n_1093) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_265), .Y(n_1021) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_266), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_269), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_270), .Y(n_992) );
OA22x2_ASAP7_75t_L g713 ( .A1(n_272), .A2(n_714), .B1(n_715), .B2(n_741), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_272), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_274), .A2(n_293), .B1(n_592), .B2(n_593), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_275), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_276), .Y(n_953) );
AOI22x1_ASAP7_75t_L g749 ( .A1(n_277), .A2(n_750), .B1(n_778), .B2(n_779), .Y(n_749) );
INVx1_ASAP7_75t_L g778 ( .A(n_277), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g1115 ( .A(n_279), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_281), .Y(n_1019) );
OA22x2_ASAP7_75t_L g945 ( .A1(n_282), .A2(n_946), .B1(n_947), .B2(n_948), .Y(n_945) );
CKINVDCx16_ASAP7_75t_R g946 ( .A(n_282), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_283), .B(n_530), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_284), .A2(n_362), .B1(n_626), .B2(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g425 ( .A(n_285), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_285), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_286), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_287), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_288), .A2(n_347), .B1(n_544), .B2(n_882), .Y(n_965) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_289), .Y(n_1069) );
CKINVDCx20_ASAP7_75t_R g1197 ( .A(n_290), .Y(n_1197) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_291), .A2(n_395), .B1(n_530), .B2(n_669), .C(n_672), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_292), .A2(n_335), .B1(n_462), .B2(n_735), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_298), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_302), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g1156 ( .A(n_304), .Y(n_1156) );
CKINVDCx20_ASAP7_75t_R g1192 ( .A(n_305), .Y(n_1192) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_307), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_309), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_311), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_312), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_313), .A2(n_830), .B1(n_831), .B2(n_856), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_313), .Y(n_830) );
XNOR2x1_ASAP7_75t_L g1089 ( .A(n_314), .B(n_1090), .Y(n_1089) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_316), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_317), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_318), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_319), .A2(n_369), .B1(n_538), .B2(n_698), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_320), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_321), .Y(n_1125) );
INVx1_ASAP7_75t_L g406 ( .A(n_324), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_325), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_326), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_327), .Y(n_1015) );
INVx1_ASAP7_75t_L g404 ( .A(n_328), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g955 ( .A(n_329), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_333), .A2(n_379), .B1(n_623), .B2(n_624), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_336), .A2(n_390), .B1(n_495), .B2(n_789), .Y(n_1097) );
XOR2xp5_ASAP7_75t_L g1148 ( .A(n_339), .B(n_1149), .Y(n_1148) );
XOR2x2_ASAP7_75t_L g1008 ( .A(n_340), .B(n_1009), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g999 ( .A(n_343), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g1176 ( .A(n_346), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_348), .B(n_820), .Y(n_1118) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_351), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_353), .A2(n_387), .B1(n_537), .B2(n_574), .Y(n_1116) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_354), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_356), .B(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_357), .A2(n_396), .B1(n_820), .B2(n_821), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g1154 ( .A(n_359), .Y(n_1154) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_361), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_363), .A2(n_374), .B1(n_710), .B2(n_1039), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_366), .A2(n_391), .B1(n_543), .B2(n_589), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g1185 ( .A(n_367), .Y(n_1185) );
CKINVDCx20_ASAP7_75t_R g935 ( .A(n_368), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_370), .B(n_671), .Y(n_1119) );
CKINVDCx20_ASAP7_75t_R g1052 ( .A(n_377), .Y(n_1052) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_378), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_381), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_384), .B(n_548), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_385), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_386), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_389), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_392), .B(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_393), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_400), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_405), .Y(n_402) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_404), .Y(n_1138) );
OAI21xp5_ASAP7_75t_L g1204 ( .A1(n_405), .A2(n_1137), .B(n_1205), .Y(n_1204) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_891), .B1(n_1132), .B2(n_1133), .C(n_1134), .Y(n_408) );
INVx1_ASAP7_75t_L g1133 ( .A(n_409), .Y(n_1133) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_633), .B1(n_889), .B2(n_890), .Y(n_409) );
INVx1_ASAP7_75t_L g890 ( .A(n_410), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_554), .B1(n_631), .B2(n_632), .Y(n_410) );
INVx1_ASAP7_75t_L g631 ( .A(n_411), .Y(n_631) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_512), .B1(n_513), .B2(n_553), .Y(n_412) );
INVx1_ASAP7_75t_L g553 ( .A(n_413), .Y(n_553) );
INVx1_ASAP7_75t_SL g511 ( .A(n_414), .Y(n_511) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_415), .B(n_469), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_450), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_439), .Y(n_416) );
INVx1_ASAP7_75t_L g658 ( .A(n_418), .Y(n_658) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g619 ( .A(n_419), .Y(n_619) );
INVx4_ASAP7_75t_L g734 ( .A(n_419), .Y(n_734) );
INVx4_ASAP7_75t_L g914 ( .A(n_419), .Y(n_914) );
INVx11_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx11_ASAP7_75t_L g520 ( .A(n_420), .Y(n_520) );
AND2x6_ASAP7_75t_L g420 ( .A(n_421), .B(n_430), .Y(n_420) );
AND2x4_ASAP7_75t_L g533 ( .A(n_421), .B(n_455), .Y(n_533) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g473 ( .A(n_422), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g438 ( .A(n_423), .B(n_428), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_423), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g483 ( .A(n_424), .B(n_428), .Y(n_483) );
AND2x2_ASAP7_75t_L g490 ( .A(n_424), .B(n_432), .Y(n_490) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_427), .Y(n_429) );
INVx2_ASAP7_75t_L g444 ( .A(n_428), .Y(n_444) );
INVx1_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
AND2x4_ASAP7_75t_L g437 ( .A(n_430), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g442 ( .A(n_430), .B(n_443), .Y(n_442) );
AND2x6_ASAP7_75t_L g482 ( .A(n_430), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
AND2x2_ASAP7_75t_L g455 ( .A(n_431), .B(n_434), .Y(n_455) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g448 ( .A(n_432), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_432), .B(n_434), .Y(n_459) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g449 ( .A(n_434), .Y(n_449) );
INVx1_ASAP7_75t_L g489 ( .A(n_434), .Y(n_489) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g620 ( .A(n_436), .Y(n_620) );
INVx2_ASAP7_75t_L g710 ( .A(n_436), .Y(n_710) );
INVx2_ASAP7_75t_L g885 ( .A(n_436), .Y(n_885) );
INVx6_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g584 ( .A(n_437), .Y(n_584) );
BUFx3_ASAP7_75t_L g735 ( .A(n_437), .Y(n_735) );
BUFx3_ASAP7_75t_L g943 ( .A(n_437), .Y(n_943) );
AND2x2_ASAP7_75t_L g464 ( .A(n_438), .B(n_448), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_438), .B(n_455), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_438), .B(n_448), .Y(n_651) );
AND2x6_ASAP7_75t_L g671 ( .A(n_438), .B(n_455), .Y(n_671) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx3_ASAP7_75t_L g583 ( .A(n_441), .Y(n_583) );
INVx3_ASAP7_75t_L g739 ( .A(n_441), .Y(n_739) );
BUFx6f_ASAP7_75t_L g854 ( .A(n_441), .Y(n_854) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g524 ( .A(n_442), .Y(n_524) );
BUFx2_ASAP7_75t_SL g623 ( .A(n_442), .Y(n_623) );
BUFx2_ASAP7_75t_SL g702 ( .A(n_442), .Y(n_702) );
AND2x2_ASAP7_75t_L g447 ( .A(n_443), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g454 ( .A(n_443), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g457 ( .A(n_443), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_443), .B(n_448), .Y(n_667) );
AND2x2_ASAP7_75t_L g488 ( .A(n_444), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g525 ( .A(n_447), .Y(n_525) );
BUFx3_ASAP7_75t_L g597 ( .A(n_447), .Y(n_597) );
BUFx3_ASAP7_75t_L g707 ( .A(n_447), .Y(n_707) );
INVx1_ASAP7_75t_L g509 ( .A(n_449), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g880 ( .A(n_453), .Y(n_880) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g541 ( .A(n_454), .Y(n_541) );
BUFx3_ASAP7_75t_L g599 ( .A(n_454), .Y(n_599) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_454), .Y(n_624) );
BUFx3_ASAP7_75t_L g644 ( .A(n_454), .Y(n_644) );
INVx1_ASAP7_75t_L g474 ( .A(n_455), .Y(n_474) );
INVx1_ASAP7_75t_L g1157 ( .A(n_456), .Y(n_1157) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g521 ( .A(n_457), .Y(n_521) );
BUFx2_ASAP7_75t_SL g593 ( .A(n_457), .Y(n_593) );
BUFx3_ASAP7_75t_L g647 ( .A(n_457), .Y(n_647) );
BUFx2_ASAP7_75t_L g708 ( .A(n_457), .Y(n_708) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_457), .Y(n_732) );
BUFx3_ASAP7_75t_L g769 ( .A(n_457), .Y(n_769) );
INVx1_ASAP7_75t_L g974 ( .A(n_457), .Y(n_974) );
AND2x2_ASAP7_75t_L g802 ( .A(n_458), .B(n_502), .Y(n_802) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x6_ASAP7_75t_L g467 ( .A(n_459), .B(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g911 ( .A(n_462), .Y(n_911) );
INVx5_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
INVx4_ASAP7_75t_L g588 ( .A(n_463), .Y(n_588) );
INVx2_ASAP7_75t_L g814 ( .A(n_463), .Y(n_814) );
BUFx3_ASAP7_75t_L g851 ( .A(n_463), .Y(n_851) );
INVx1_ASAP7_75t_L g1080 ( .A(n_463), .Y(n_1080) );
INVx8_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_465), .Y(n_1054) );
BUFx4f_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g544 ( .A(n_466), .Y(n_544) );
BUFx2_ASAP7_75t_L g626 ( .A(n_466), .Y(n_626) );
BUFx2_ASAP7_75t_L g654 ( .A(n_466), .Y(n_654) );
BUFx2_ASAP7_75t_L g1163 ( .A(n_466), .Y(n_1163) );
INVx6_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g589 ( .A(n_467), .Y(n_589) );
INVx1_ASAP7_75t_L g771 ( .A(n_467), .Y(n_771) );
INVx1_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .C(n_497), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_475), .B2(n_476), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_472), .A2(n_476), .B1(n_758), .B2(n_759), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_472), .A2(n_563), .B1(n_928), .B2(n_929), .Y(n_927) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_473), .Y(n_561) );
INVx2_ASAP7_75t_L g865 ( .A(n_473), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_473), .A2(n_476), .B1(n_1093), .B2(n_1094), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_476), .A2(n_863), .B1(n_864), .B2(n_866), .Y(n_862) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g528 ( .A(n_477), .Y(n_528) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g563 ( .A(n_478), .Y(n_563) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_484), .B1(n_485), .B2(n_491), .C(n_492), .Y(n_479) );
INVx1_ASAP7_75t_L g678 ( .A(n_480), .Y(n_678) );
OAI222xp33_ASAP7_75t_L g1068 ( .A1(n_480), .A2(n_485), .B1(n_572), .B2(n_1069), .C1(n_1070), .C2(n_1071), .Y(n_1068) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_481), .A2(n_689), .B(n_690), .Y(n_688) );
INVx4_ASAP7_75t_L g1060 ( .A(n_481), .Y(n_1060) );
OAI21xp5_ASAP7_75t_L g1114 ( .A1(n_481), .A2(n_1115), .B(n_1116), .Y(n_1114) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
INVx2_ASAP7_75t_SL g570 ( .A(n_482), .Y(n_570) );
INVx2_ASAP7_75t_L g718 ( .A(n_482), .Y(n_718) );
INVx2_ASAP7_75t_L g753 ( .A(n_482), .Y(n_753) );
BUFx3_ASAP7_75t_L g825 ( .A(n_482), .Y(n_825) );
INVx1_ASAP7_75t_L g507 ( .A(n_483), .Y(n_507) );
AND2x4_ASAP7_75t_L g538 ( .A(n_483), .B(n_509), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_485), .A2(n_753), .B1(n_754), .B2(n_755), .C(n_756), .Y(n_752) );
OAI222xp33_ASAP7_75t_L g995 ( .A1(n_485), .A2(n_870), .B1(n_996), .B2(n_997), .C1(n_998), .C2(n_999), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_487), .Y(n_568) );
BUFx4f_ASAP7_75t_SL g679 ( .A(n_487), .Y(n_679) );
BUFx2_ASAP7_75t_L g721 ( .A(n_487), .Y(n_721) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_489), .Y(n_496) );
AND2x4_ASAP7_75t_L g495 ( .A(n_490), .B(n_496), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_490), .B(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g535 ( .A(n_490), .B(n_536), .Y(n_535) );
INVxp67_ASAP7_75t_L g998 ( .A(n_493), .Y(n_998) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx3_ASAP7_75t_L g722 ( .A(n_494), .Y(n_722) );
INVx2_ASAP7_75t_L g905 ( .A(n_494), .Y(n_905) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx12f_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_495), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B1(n_503), .B2(n_504), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_499), .A2(n_506), .B1(n_612), .B2(n_613), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_499), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
INVx3_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g674 ( .A(n_500), .Y(n_674) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g577 ( .A(n_501), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_501), .A2(n_763), .B1(n_899), .B2(n_900), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_501), .A2(n_506), .B1(n_934), .B2(n_935), .Y(n_933) );
OAI22xp33_ASAP7_75t_SL g959 ( .A1(n_501), .A2(n_504), .B1(n_960), .B2(n_961), .Y(n_959) );
HB1xp67_ASAP7_75t_L g1020 ( .A(n_501), .Y(n_1020) );
OAI22xp5_ASAP7_75t_SL g576 ( .A1(n_504), .A2(n_577), .B1(n_578), .B2(n_579), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_504), .A2(n_577), .B1(n_875), .B2(n_876), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_504), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1018) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g763 ( .A(n_505), .Y(n_763) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g676 ( .A(n_506), .Y(n_676) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AO22x1_ASAP7_75t_L g601 ( .A1(n_514), .A2(n_515), .B1(n_602), .B2(n_629), .Y(n_601) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
XOR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_552), .Y(n_515) );
NAND4xp75_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .C(n_539), .D(n_545), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx5_ASAP7_75t_SL g592 ( .A(n_520), .Y(n_592) );
INVx4_ASAP7_75t_L g1039 ( .A(n_520), .Y(n_1039) );
INVx1_ASAP7_75t_L g1083 ( .A(n_520), .Y(n_1083) );
INVx2_ASAP7_75t_SL g1123 ( .A(n_520), .Y(n_1123) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g938 ( .A(n_524), .Y(n_938) );
OA211x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .C(n_534), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_528), .A2(n_561), .B1(n_606), .B2(n_607), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_528), .A2(n_561), .B1(n_907), .B2(n_908), .Y(n_906) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx5_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g728 ( .A(n_532), .Y(n_728) );
INVx2_ASAP7_75t_L g792 ( .A(n_532), .Y(n_792) );
INVx2_ASAP7_75t_L g820 ( .A(n_532), .Y(n_820) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g698 ( .A(n_535), .Y(n_698) );
INVx1_ASAP7_75t_L g726 ( .A(n_535), .Y(n_726) );
BUFx2_ASAP7_75t_L g994 ( .A(n_535), .Y(n_994) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_535), .Y(n_1074) );
INVx1_ASAP7_75t_SL g844 ( .A(n_537), .Y(n_844) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_SL g699 ( .A(n_538), .Y(n_699) );
BUFx3_ASAP7_75t_L g789 ( .A(n_538), .Y(n_789) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g972 ( .A(n_541), .Y(n_972) );
HB1xp67_ASAP7_75t_L g1178 ( .A(n_541), .Y(n_1178) );
INVx2_ASAP7_75t_L g834 ( .A(n_546), .Y(n_834) );
INVx2_ASAP7_75t_SL g870 ( .A(n_546), .Y(n_870) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g692 ( .A(n_548), .Y(n_692) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx4f_ASAP7_75t_SL g680 ( .A(n_551), .Y(n_680) );
INVx2_ASAP7_75t_L g632 ( .A(n_554), .Y(n_632) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_600), .B1(n_601), .B2(n_630), .Y(n_555) );
INVx2_ASAP7_75t_L g630 ( .A(n_556), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_556), .A2(n_630), .B1(n_713), .B2(n_742), .Y(n_712) );
XNOR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_580), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_565), .C(n_576), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g952 ( .A(n_561), .Y(n_952) );
OAI221xp5_ASAP7_75t_SL g988 ( .A1(n_561), .A2(n_989), .B1(n_990), .B2(n_992), .C(n_993), .Y(n_988) );
BUFx3_ASAP7_75t_L g954 ( .A(n_563), .Y(n_954) );
INVx2_ASAP7_75t_L g991 ( .A(n_563), .Y(n_991) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_570), .B2(n_571), .C1(n_572), .C2(n_575), .Y(n_565) );
OAI222xp33_ASAP7_75t_L g1191 ( .A1(n_566), .A2(n_870), .B1(n_872), .B2(n_1192), .C1(n_1193), .C2(n_1194), .Y(n_1191) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_570), .A2(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_577), .A2(n_763), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_590), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
INVx1_ASAP7_75t_L g776 ( .A(n_584), .Y(n_776) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g704 ( .A(n_588), .Y(n_704) );
BUFx6f_ASAP7_75t_L g882 ( .A(n_588), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
INVx1_ASAP7_75t_L g980 ( .A(n_593), .Y(n_980) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx4f_ASAP7_75t_SL g617 ( .A(n_597), .Y(n_617) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g629 ( .A(n_602), .Y(n_629) );
INVx2_ASAP7_75t_L g627 ( .A(n_603), .Y(n_627) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_614), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .C(n_611), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_621), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx2_ASAP7_75t_L g660 ( .A(n_620), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g663 ( .A(n_623), .Y(n_663) );
INVx4_ASAP7_75t_L g848 ( .A(n_624), .Y(n_848) );
INVx1_ASAP7_75t_L g889 ( .A(n_633), .Y(n_889) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_745), .Y(n_633) );
XOR2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_683), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g682 ( .A(n_638), .Y(n_682) );
AND4x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_655), .C(n_668), .D(n_677), .Y(n_638) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_640), .B(n_648), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_645), .B2(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_650), .A2(n_1052), .B1(n_1053), .B2(n_1054), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_650), .A2(n_1160), .B1(n_1161), .B2(n_1162), .Y(n_1159) );
BUFx2_ASAP7_75t_R g650 ( .A(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_661), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_660), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_660), .A2(n_665), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_661) );
OAI221xp5_ASAP7_75t_SL g978 ( .A1(n_665), .A2(n_979), .B1(n_980), .B2(n_981), .C(n_982), .Y(n_978) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g969 ( .A(n_666), .Y(n_969) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g695 ( .A(n_670), .Y(n_695) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
BUFx4f_ASAP7_75t_L g821 ( .A(n_671), .Y(n_821) );
BUFx2_ASAP7_75t_L g839 ( .A(n_671), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_674), .A2(n_868), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_674), .A2(n_676), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_674), .A2(n_763), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_712), .B1(n_743), .B2(n_744), .Y(n_683) );
INVx2_ASAP7_75t_L g744 ( .A(n_684), .Y(n_744) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
XOR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_711), .Y(n_685) );
NAND3x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_700), .C(n_705), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_688), .B(n_693), .Y(n_687) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .C(n_697), .Y(n_693) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
BUFx2_ASAP7_75t_L g777 ( .A(n_707), .Y(n_777) );
INVx1_ASAP7_75t_L g1152 ( .A(n_707), .Y(n_1152) );
INVx1_ASAP7_75t_L g743 ( .A(n_712), .Y(n_743) );
INVx1_ASAP7_75t_L g742 ( .A(n_713), .Y(n_742) );
INVx2_ASAP7_75t_L g741 ( .A(n_715), .Y(n_741) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_729), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_723), .Y(n_716) );
OAI21xp5_ASAP7_75t_SL g717 ( .A1(n_718), .A2(n_719), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g868 ( .A(n_721), .Y(n_868) );
INVx2_ASAP7_75t_L g872 ( .A(n_722), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g842 ( .A(n_726), .Y(n_842) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_736), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx3_ASAP7_75t_L g1183 ( .A(n_735), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI221xp5_ASAP7_75t_SL g1175 ( .A1(n_739), .A2(n_1176), .B1(n_1177), .B2(n_1179), .C(n_1180), .Y(n_1175) );
XNOR2x1_ASAP7_75t_L g745 ( .A(n_746), .B(n_805), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_780), .B1(n_781), .B2(n_804), .Y(n_748) );
INVx1_ASAP7_75t_L g804 ( .A(n_749), .Y(n_804) );
INVx2_ASAP7_75t_SL g779 ( .A(n_750), .Y(n_779) );
AND2x4_ASAP7_75t_L g750 ( .A(n_751), .B(n_764), .Y(n_750) );
NOR3xp33_ASAP7_75t_SL g751 ( .A(n_752), .B(n_757), .C(n_760), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_753), .A2(n_787), .B(n_788), .Y(n_786) );
OAI21xp33_ASAP7_75t_L g901 ( .A1(n_753), .A2(n_902), .B(n_903), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g1014 ( .A1(n_753), .A2(n_872), .B1(n_1015), .B2(n_1016), .C(n_1017), .Y(n_1014) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_772), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_770), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
HB1xp67_ASAP7_75t_L g1181 ( .A(n_769), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
XOR2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_803), .Y(n_783) );
NAND2x1p5_ASAP7_75t_L g784 ( .A(n_785), .B(n_795), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_790), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .C(n_794), .Y(n_790) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_799), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
BUFx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_858), .B2(n_859), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AO22x1_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_828), .B1(n_829), .B2(n_857), .Y(n_808) );
INVx1_ASAP7_75t_SL g857 ( .A(n_809), .Y(n_857) );
NOR4xp75_ASAP7_75t_L g810 ( .A(n_811), .B(n_815), .C(n_818), .D(n_823), .Y(n_810) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_812), .B(n_813), .Y(n_811) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_814), .Y(n_983) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_816), .B(n_817), .Y(n_815) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_819), .B(n_822), .Y(n_818) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_820), .Y(n_1165) );
OAI21xp5_ASAP7_75t_SL g823 ( .A1(n_824), .A2(n_826), .B(n_827), .Y(n_823) );
OAI21xp33_ASAP7_75t_SL g956 ( .A1(n_824), .A2(n_957), .B(n_958), .Y(n_956) );
OAI21xp33_ASAP7_75t_L g1095 ( .A1(n_824), .A2(n_1096), .B(n_1097), .Y(n_1095) );
INVx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g856 ( .A(n_831), .Y(n_856) );
NAND3x1_ASAP7_75t_L g831 ( .A(n_832), .B(n_845), .C(n_852), .Y(n_831) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_837), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g833 ( .A1(n_834), .A2(n_835), .B(n_836), .Y(n_833) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_840), .C(n_841), .Y(n_837) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
INVx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx4_ASAP7_75t_L g1034 ( .A(n_848), .Y(n_1034) );
INVx3_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_SL g888 ( .A(n_860), .Y(n_888) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_877), .Y(n_860) );
NOR3xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_867), .C(n_874), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g1011 ( .A1(n_864), .A2(n_990), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OAI222xp33_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_870), .B2(n_871), .C1(n_872), .C2(n_873), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g877 ( .A(n_878), .B(n_883), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_881), .Y(n_878) );
NAND2xp5_ASAP7_75t_SL g883 ( .A(n_884), .B(n_886), .Y(n_883) );
INVx1_ASAP7_75t_L g1132 ( .A(n_891), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_1004), .B2(n_1131), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
AOI22x1_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_917), .B1(n_918), .B2(n_1003), .Y(n_893) );
INVx1_ASAP7_75t_L g1003 ( .A(n_894), .Y(n_1003) );
INVx2_ASAP7_75t_L g916 ( .A(n_896), .Y(n_916) );
NAND2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_909), .Y(n_896) );
NOR3xp33_ASAP7_75t_SL g897 ( .A(n_898), .B(n_901), .C(n_906), .Y(n_897) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
AND4x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_912), .C(n_913), .D(n_915), .Y(n_909) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
AO22x2_ASAP7_75t_SL g918 ( .A1(n_919), .A2(n_920), .B1(n_975), .B2(n_1002), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_922), .B1(n_944), .B2(n_945), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AND3x1_ASAP7_75t_L g925 ( .A(n_926), .B(n_936), .C(n_940), .Y(n_925) );
NOR3xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .C(n_933), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
AND2x2_ASAP7_75t_L g936 ( .A(n_937), .B(n_939), .Y(n_936) );
AND2x2_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx2_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_962), .Y(n_948) );
NOR3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_956), .C(n_959), .Y(n_949) );
OAI22xp5_ASAP7_75t_SL g950 ( .A1(n_951), .A2(n_953), .B1(n_954), .B2(n_955), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_951), .A2(n_990), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
NOR3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_966), .C(n_970), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_965), .Y(n_963) );
OAI221xp5_ASAP7_75t_SL g1182 ( .A1(n_969), .A2(n_1183), .B1(n_1184), .B2(n_1185), .C(n_1186), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_971), .A2(n_972), .B1(n_973), .B2(n_974), .Y(n_970) );
INVx2_ASAP7_75t_L g1002 ( .A(n_975), .Y(n_1002) );
INVx1_ASAP7_75t_L g1001 ( .A(n_976), .Y(n_1001) );
AND2x2_ASAP7_75t_SL g976 ( .A(n_977), .B(n_987), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_984), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_986), .Y(n_984) );
NOR2xp33_ASAP7_75t_SL g987 ( .A(n_988), .B(n_995), .Y(n_987) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1004), .Y(n_1131) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1063), .B1(n_1129), .B2(n_1130), .Y(n_1004) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1005), .Y(n_1129) );
XOR2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1044), .Y(n_1005) );
OAI22xp5_ASAP7_75t_SL g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1029), .B2(n_1030), .Y(n_1006) );
OA22x2_ASAP7_75t_L g1087 ( .A1(n_1007), .A2(n_1008), .B1(n_1088), .B2(n_1126), .Y(n_1087) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1022), .Y(n_1009) );
NOR3xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1014), .C(n_1018), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1026), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
NAND4xp75_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1036), .C(n_1040), .D(n_1043), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1035), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_1039), .Y(n_1155) );
AND2x2_ASAP7_75t_SL g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1045), .Y(n_1062) );
AND4x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1050), .C(n_1055), .D(n_1059), .Y(n_1045) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1063), .Y(n_1130) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1086), .B1(n_1127), .B2(n_1128), .Y(n_1063) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1064), .Y(n_1127) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1066), .Y(n_1085) );
NAND3xp33_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1076), .C(n_1081), .Y(n_1066) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1072), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1075), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1084), .Y(n_1081) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1087), .Y(n_1128) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1088), .Y(n_1126) );
XOR2x2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1108), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1101), .Y(n_1090) );
NOR3xp33_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1095), .C(n_1098), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
XOR2x2_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1125), .Y(n_1108) );
NAND3x1_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1113), .C(n_1121), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
NOR2x1_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1117), .Y(n_1113) );
NAND3xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1119), .C(n_1120), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1124), .Y(n_1121) );
INVx1_ASAP7_75t_SL g1134 ( .A(n_1135), .Y(n_1134) );
NOR2x1_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1140), .Y(n_1135) );
OR2x2_ASAP7_75t_SL g1202 ( .A(n_1136), .B(n_1141), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1139), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1137), .B(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1138), .B(n_1171), .Y(n_1205) );
CKINVDCx16_ASAP7_75t_R g1171 ( .A(n_1139), .Y(n_1171) );
CKINVDCx20_ASAP7_75t_R g1140 ( .A(n_1141), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1146), .Y(n_1144) );
OAI222xp33_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1170), .B1(n_1172), .B2(n_1198), .C1(n_1200), .C2(n_1203), .Y(n_1147) );
AND4x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1158), .C(n_1164), .D(n_1169), .Y(n_1149) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1155), .B1(n_1156), .B2(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_SL g1199 ( .A(n_1173), .Y(n_1199) );
AND2x2_ASAP7_75t_SL g1173 ( .A(n_1174), .B(n_1187), .Y(n_1173) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1182), .Y(n_1174) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
NOR3xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1191), .C(n_1195), .Y(n_1187) );
CKINVDCx20_ASAP7_75t_R g1200 ( .A(n_1201), .Y(n_1200) );
CKINVDCx20_ASAP7_75t_R g1201 ( .A(n_1202), .Y(n_1201) );
CKINVDCx16_ASAP7_75t_R g1203 ( .A(n_1204), .Y(n_1203) );
endmodule