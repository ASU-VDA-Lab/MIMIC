module real_aes_16048_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AND2x4_ASAP7_75t_L g116 ( .A(n_0), .B(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_1), .A2(n_525), .B1(n_526), .B2(n_528), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_1), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_2), .A2(n_35), .B1(n_152), .B2(n_244), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_3), .A2(n_12), .B1(n_557), .B2(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g117 ( .A(n_4), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_5), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_6), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_7), .A2(n_13), .B1(n_558), .B2(n_594), .Y(n_593) );
XNOR2xp5_ASAP7_75t_L g526 ( .A(n_8), .B(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g112 ( .A(n_9), .B(n_31), .Y(n_112) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_10), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_11), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_14), .B(n_167), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_15), .A2(n_102), .B1(n_197), .B2(n_557), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_16), .A2(n_32), .B1(n_575), .B2(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_17), .B(n_167), .Y(n_572) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_18), .A2(n_48), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_19), .B(n_248), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_20), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_20), .A2(n_95), .B1(n_630), .B2(n_864), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_21), .A2(n_39), .B1(n_204), .B2(n_219), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_22), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_23), .A2(n_45), .B1(n_219), .B2(n_557), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_24), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_25), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_26), .B(n_227), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_27), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g527 ( .A(n_28), .B(n_40), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_29), .B(n_145), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_30), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_33), .A2(n_86), .B1(n_152), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_34), .A2(n_38), .B1(n_152), .B2(n_560), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_36), .A2(n_51), .B1(n_557), .B2(n_612), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_37), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_41), .B(n_167), .Y(n_215) );
INVx2_ASAP7_75t_L g128 ( .A(n_42), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_43), .B(n_200), .Y(n_242) );
BUFx3_ASAP7_75t_L g111 ( .A(n_44), .Y(n_111) );
INVx1_ASAP7_75t_L g878 ( .A(n_44), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_46), .B(n_186), .Y(n_250) );
XOR2x2_ASAP7_75t_L g134 ( .A(n_47), .B(n_135), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_47), .A2(n_866), .B1(n_867), .B2(n_870), .Y(n_865) );
INVx1_ASAP7_75t_L g870 ( .A(n_47), .Y(n_870) );
AND2x2_ASAP7_75t_L g278 ( .A(n_49), .B(n_186), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_50), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_52), .B(n_227), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_53), .B(n_204), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_54), .A2(n_73), .B1(n_204), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_55), .A2(n_76), .B1(n_152), .B2(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_56), .B(n_308), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_57), .A2(n_156), .B(n_165), .C(n_271), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_58), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_59), .A2(n_99), .B1(n_557), .B2(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g148 ( .A(n_60), .Y(n_148) );
AND2x4_ASAP7_75t_L g170 ( .A(n_61), .B(n_171), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_62), .A2(n_63), .B1(n_219), .B2(n_231), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_64), .A2(n_83), .B1(n_868), .B2(n_869), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_64), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_65), .B(n_145), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_66), .B(n_186), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_67), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_68), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g171 ( .A(n_69), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_70), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_71), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_72), .B(n_145), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_74), .B(n_152), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_75), .B(n_200), .C(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_77), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g158 ( .A(n_78), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_79), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_80), .B(n_167), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_81), .B(n_161), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_82), .A2(n_98), .B1(n_165), .B2(n_219), .Y(n_544) );
INVx1_ASAP7_75t_L g869 ( .A(n_83), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_84), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_85), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_87), .A2(n_92), .B1(n_226), .B2(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_88), .B(n_167), .Y(n_199) );
NAND2xp33_ASAP7_75t_SL g184 ( .A(n_89), .B(n_155), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_90), .B(n_198), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_91), .B(n_145), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_93), .Y(n_597) );
INVx1_ASAP7_75t_L g115 ( .A(n_94), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_94), .B(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g864 ( .A(n_95), .Y(n_864) );
NAND2xp33_ASAP7_75t_L g576 ( .A(n_96), .B(n_167), .Y(n_576) );
NAND2xp33_ASAP7_75t_L g154 ( .A(n_97), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_100), .B(n_186), .Y(n_310) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_101), .B(n_155), .C(n_179), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_103), .B(n_152), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_104), .B(n_227), .Y(n_306) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_118), .B(n_889), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx12f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx12f_ASAP7_75t_L g892 ( .A(n_108), .Y(n_892) );
OR2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_113), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g851 ( .A(n_110), .B(n_124), .Y(n_851) );
NOR2x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_112), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_114), .Y(n_855) );
AND3x2_ASAP7_75t_L g876 ( .A(n_114), .B(n_131), .C(n_877), .Y(n_876) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g124 ( .A(n_115), .Y(n_124) );
OR2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_879), .Y(n_118) );
OAI211xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_132), .B(n_529), .C(n_856), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
NOR2xp67_ASAP7_75t_SL g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx4_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
NOR2x1_ASAP7_75t_R g854 ( .A(n_125), .B(n_855), .Y(n_854) );
INVx5_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_128), .B(n_850), .Y(n_849) );
INVx3_ASAP7_75t_L g859 ( .A(n_128), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x6_ASAP7_75t_SL g881 ( .A(n_131), .B(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B1(n_523), .B2(n_524), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_135), .Y(n_873) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_455), .Y(n_135) );
NAND4xp25_ASAP7_75t_L g136 ( .A(n_137), .B(n_330), .C(n_370), .D(n_419), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_138), .B(n_279), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_189), .B1(n_251), .B2(n_260), .Y(n_138) );
INVx1_ASAP7_75t_L g451 ( .A(n_139), .Y(n_451) );
INVx1_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_140), .B(n_298), .Y(n_367) );
AND2x2_ASAP7_75t_L g398 ( .A(n_140), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_172), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_141), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g322 ( .A(n_141), .Y(n_322) );
AND2x2_ASAP7_75t_L g497 ( .A(n_141), .B(n_365), .Y(n_497) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx2_ASAP7_75t_L g262 ( .A(n_142), .Y(n_262) );
AND2x2_ASAP7_75t_L g350 ( .A(n_142), .B(n_312), .Y(n_350) );
AND2x2_ASAP7_75t_L g394 ( .A(n_142), .B(n_299), .Y(n_394) );
OR2x2_ASAP7_75t_L g412 ( .A(n_142), .B(n_413), .Y(n_412) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g316 ( .A(n_143), .B(n_299), .Y(n_316) );
BUFx2_ASAP7_75t_L g373 ( .A(n_143), .Y(n_373) );
OR2x2_ASAP7_75t_L g381 ( .A(n_143), .B(n_339), .Y(n_381) );
INVx1_ASAP7_75t_L g436 ( .A(n_143), .Y(n_436) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx2_ASAP7_75t_L g584 ( .A(n_145), .Y(n_584) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_SL g168 ( .A(n_146), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_SL g175 ( .A(n_146), .Y(n_175) );
INVx2_ASAP7_75t_L g211 ( .A(n_146), .Y(n_211) );
BUFx3_ASAP7_75t_L g540 ( .A(n_146), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_146), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g568 ( .A(n_146), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_146), .B(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_146), .B(n_607), .Y(n_606) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_159), .B(n_168), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_156), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g275 ( .A1(n_152), .A2(n_219), .B1(n_276), .B2(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g558 ( .A(n_152), .Y(n_558) );
INVx4_ASAP7_75t_L g560 ( .A(n_152), .Y(n_560) );
INVx1_ASAP7_75t_L g612 ( .A(n_152), .Y(n_612) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_153), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_153), .Y(n_165) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_153), .Y(n_167) );
INVx1_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
INVx1_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_153), .Y(n_219) );
INVx1_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_153), .Y(n_231) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_153), .Y(n_244) );
INVx2_ASAP7_75t_L g273 ( .A(n_153), .Y(n_273) );
INVx2_ASAP7_75t_L g204 ( .A(n_155), .Y(n_204) );
INVx1_ASAP7_75t_L g575 ( .A(n_155), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_156), .A2(n_182), .B(n_184), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_156), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_156), .A2(n_303), .B(n_304), .Y(n_302) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g163 ( .A(n_158), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
BUFx8_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B1(n_164), .B2(n_166), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_161), .A2(n_202), .B(n_203), .Y(n_201) );
INVx2_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx3_ASAP7_75t_L g233 ( .A(n_163), .Y(n_233) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_167), .A2(n_178), .B(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g248 ( .A(n_167), .Y(n_248) );
INVx3_ASAP7_75t_L g557 ( .A(n_167), .Y(n_557) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_169), .A2(n_177), .B(n_181), .Y(n_176) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_169), .A2(n_195), .B(n_201), .Y(n_194) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_169), .A2(n_213), .B(n_216), .Y(n_212) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_169), .A2(n_241), .B(n_245), .Y(n_240) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_169), .A2(n_302), .B(n_305), .Y(n_301) );
BUFx10_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx10_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
INVx1_ASAP7_75t_L g547 ( .A(n_170), .Y(n_547) );
AND2x2_ASAP7_75t_L g263 ( .A(n_172), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g375 ( .A(n_172), .B(n_352), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_172), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g413 ( .A(n_173), .Y(n_413) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_173), .Y(n_418) );
AND2x2_ASAP7_75t_L g435 ( .A(n_173), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g325 ( .A(n_174), .B(n_265), .Y(n_325) );
INVx1_ASAP7_75t_L g339 ( .A(n_174), .Y(n_339) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_185), .Y(n_174) );
INVx1_ASAP7_75t_L g249 ( .A(n_179), .Y(n_249) );
INVx1_ASAP7_75t_L g545 ( .A(n_179), .Y(n_545) );
INVx1_ASAP7_75t_SL g561 ( .A(n_179), .Y(n_561) );
INVx1_ASAP7_75t_L g603 ( .A(n_183), .Y(n_603) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g193 ( .A(n_187), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_187), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_187), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
INVx2_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
NAND2x1_ASAP7_75t_L g189 ( .A(n_190), .B(n_206), .Y(n_189) );
AND2x4_ASAP7_75t_L g500 ( .A(n_190), .B(n_428), .Y(n_500) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_191), .Y(n_259) );
BUFx3_ASAP7_75t_L g294 ( .A(n_191), .Y(n_294) );
INVx1_ASAP7_75t_L g360 ( .A(n_191), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_191), .B(n_209), .Y(n_363) );
AND2x2_ASAP7_75t_L g388 ( .A(n_191), .B(n_239), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_191), .Y(n_391) );
AND2x2_ASAP7_75t_L g423 ( .A(n_191), .B(n_288), .Y(n_423) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_205), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_193), .A2(n_194), .B(n_205), .Y(n_289) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_193), .A2(n_301), .B(n_310), .Y(n_300) );
OAI21xp33_ASAP7_75t_SL g328 ( .A1(n_193), .A2(n_301), .B(n_310), .Y(n_328) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .C(n_200), .Y(n_195) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_200), .A2(n_217), .B(n_218), .Y(n_216) );
INVx6_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
O2A1O1Ixp5_ASAP7_75t_L g570 ( .A1(n_200), .A2(n_560), .B(n_571), .C(n_572), .Y(n_570) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_221), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g332 ( .A(n_208), .B(n_318), .Y(n_332) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g358 ( .A(n_210), .B(n_345), .Y(n_358) );
AND2x2_ASAP7_75t_L g387 ( .A(n_210), .B(n_223), .Y(n_387) );
OR2x2_ASAP7_75t_L g483 ( .A(n_210), .B(n_223), .Y(n_483) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_210) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_211), .A2(n_240), .B(n_250), .Y(n_239) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_257) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_211), .A2(n_240), .B(n_250), .Y(n_288) );
INVx2_ASAP7_75t_L g226 ( .A(n_219), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_219), .A2(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g362 ( .A(n_221), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g511 ( .A(n_221), .Y(n_511) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_222), .Y(n_253) );
OR2x2_ASAP7_75t_L g445 ( .A(n_222), .B(n_255), .Y(n_445) );
INVx1_ASAP7_75t_L g467 ( .A(n_222), .Y(n_467) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_239), .Y(n_222) );
AND2x2_ASAP7_75t_L g283 ( .A(n_223), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g318 ( .A(n_223), .B(n_288), .Y(n_318) );
INVx1_ASAP7_75t_L g345 ( .A(n_223), .Y(n_345) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_223), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_223), .B(n_239), .Y(n_432) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_234), .A3(n_235), .B(n_236), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_229), .B1(n_230), .B2(n_232), .Y(n_224) );
INVx1_ASAP7_75t_L g594 ( .A(n_227), .Y(n_594) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_229), .A2(n_542), .B1(n_544), .B2(n_545), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_229), .A2(n_556), .B1(n_559), .B2(n_561), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_229), .A2(n_574), .B(n_576), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_229), .A2(n_232), .B1(n_582), .B2(n_583), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_229), .A2(n_561), .B1(n_593), .B2(n_595), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_229), .A2(n_232), .B1(n_602), .B2(n_604), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_229), .A2(n_232), .B1(n_611), .B2(n_613), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_229), .A2(n_232), .B1(n_627), .B2(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g605 ( .A(n_231), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_232), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g309 ( .A(n_233), .Y(n_309) );
INVx2_ASAP7_75t_L g267 ( .A(n_234), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_234), .B(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g596 ( .A(n_234), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g268 ( .A(n_235), .Y(n_268) );
AO31x2_ASAP7_75t_L g580 ( .A1(n_235), .A2(n_581), .A3(n_584), .B(n_585), .Y(n_580) );
AO31x2_ASAP7_75t_L g591 ( .A1(n_235), .A2(n_554), .A3(n_592), .B(n_596), .Y(n_591) );
AO31x2_ASAP7_75t_L g600 ( .A1(n_235), .A2(n_540), .A3(n_601), .B(n_606), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
BUFx2_ASAP7_75t_L g554 ( .A(n_238), .Y(n_554) );
AND2x2_ASAP7_75t_L g369 ( .A(n_239), .B(n_289), .Y(n_369) );
INVx2_ASAP7_75t_L g308 ( .A(n_244), .Y(n_308) );
AOI21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_249), .Y(n_245) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR3x1_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .C(n_258), .Y(n_252) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_255), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g317 ( .A(n_255), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g368 ( .A(n_255), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g408 ( .A(n_255), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_255), .B(n_431), .Y(n_463) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_256), .B(n_344), .Y(n_404) );
AND2x2_ASAP7_75t_L g428 ( .A(n_256), .B(n_288), .Y(n_428) );
BUFx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
BUFx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g439 ( .A(n_259), .B(n_318), .Y(n_439) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_262), .B(n_325), .Y(n_504) );
AND2x4_ASAP7_75t_L g496 ( .A(n_263), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_263), .B(n_316), .Y(n_510) );
INVx2_ASAP7_75t_L g312 ( .A(n_264), .Y(n_312) );
INVx1_ASAP7_75t_L g315 ( .A(n_264), .Y(n_315) );
INVx2_ASAP7_75t_L g400 ( .A(n_264), .Y(n_400) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g384 ( .A(n_265), .Y(n_384) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B(n_278), .Y(n_265) );
NOR2xp67_ASAP7_75t_SL g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g609 ( .A(n_267), .Y(n_609) );
INVx1_ASAP7_75t_L g562 ( .A(n_268), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_SL g543 ( .A(n_273), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_319), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_295), .B1(n_313), .B2(n_317), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B(n_290), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g347 ( .A(n_283), .B(n_294), .Y(n_347) );
AND2x2_ASAP7_75t_L g507 ( .A(n_283), .B(n_388), .Y(n_507) );
BUFx2_ASAP7_75t_L g378 ( .A(n_284), .Y(n_378) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g377 ( .A(n_287), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g292 ( .A(n_288), .Y(n_292) );
INVx1_ASAP7_75t_L g344 ( .A(n_288), .Y(n_344) );
INVx1_ASAP7_75t_L g469 ( .A(n_289), .Y(n_469) );
AOI31xp33_ASAP7_75t_L g487 ( .A1(n_290), .A2(n_488), .A3(n_489), .B(n_490), .Y(n_487) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_292), .B(n_387), .Y(n_486) );
INVx2_ASAP7_75t_L g514 ( .A(n_292), .Y(n_514) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_293), .Y(n_329) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g342 ( .A(n_294), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_294), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g472 ( .A(n_294), .B(n_432), .Y(n_472) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_311), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g383 ( .A(n_299), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g352 ( .A(n_300), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_309), .Y(n_305) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_315), .Y(n_336) );
INVx1_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
INVx1_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
AND2x2_ASAP7_75t_L g417 ( .A(n_316), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g473 ( .A(n_316), .B(n_400), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_317), .A2(n_390), .B(n_392), .Y(n_389) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_329), .Y(n_319) );
NAND3x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .C(n_326), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g491 ( .A(n_322), .B(n_411), .Y(n_491) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2x1_ASAP7_75t_SL g444 ( .A(n_324), .B(n_356), .Y(n_444) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g364 ( .A(n_325), .B(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_326), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_326), .B(n_435), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_326), .B(n_435), .Y(n_508) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g411 ( .A(n_328), .B(n_384), .Y(n_411) );
AND2x2_ASAP7_75t_L g331 ( .A(n_329), .B(n_332), .Y(n_331) );
AOI221x1_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_333), .B1(n_340), .B2(n_349), .C(n_353), .Y(n_330) );
AOI32xp33_ASAP7_75t_L g512 ( .A1(n_332), .A2(n_513), .A3(n_518), .B1(n_519), .B2(n_521), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_337), .B(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g351 ( .A(n_339), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_339), .Y(n_355) );
OR2x2_ASAP7_75t_L g468 ( .A(n_339), .B(n_469), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_346), .C(n_348), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g390 ( .A(n_343), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g407 ( .A(n_343), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_346), .A2(n_443), .B1(n_445), .B2(n_446), .Y(n_442) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g520 ( .A(n_350), .Y(n_520) );
INVx2_ASAP7_75t_L g365 ( .A(n_352), .Y(n_365) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B(n_361), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g489 ( .A(n_358), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_359), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_366), .B2(n_368), .Y(n_361) );
AND2x4_ASAP7_75t_L g458 ( .A(n_364), .B(n_373), .Y(n_458) );
INVx1_ASAP7_75t_L g517 ( .A(n_365), .Y(n_517) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g396 ( .A(n_369), .B(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_369), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_369), .B(n_397), .Y(n_488) );
AOI211x1_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_377), .B(n_379), .C(n_405), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR3x2_ASAP7_75t_L g480 ( .A(n_373), .B(n_375), .C(n_376), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_374), .A2(n_396), .B1(n_398), .B2(n_401), .Y(n_395) );
NOR2x1p5_ASAP7_75t_SL g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_375), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g397 ( .A(n_378), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_385), .B(n_389), .C(n_395), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_387), .B(n_391), .Y(n_402) );
INVx1_ASAP7_75t_L g429 ( .A(n_387), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_387), .B(n_494), .Y(n_502) );
OAI32xp33_ASAP7_75t_L g477 ( .A1(n_388), .A2(n_433), .A3(n_478), .B1(n_480), .B2(n_481), .Y(n_477) );
INVx1_ASAP7_75t_L g494 ( .A(n_388), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_388), .B(n_408), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_391), .B(n_425), .Y(n_460) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g438 ( .A(n_397), .B(n_423), .Y(n_438) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g415 ( .A(n_403), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B1(n_414), .B2(n_416), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g453 ( .A(n_410), .Y(n_453) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g434 ( .A(n_411), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_411), .B(n_418), .Y(n_522) );
INVx1_ASAP7_75t_SL g448 ( .A(n_412), .Y(n_448) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_442), .C(n_449), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_433), .B(n_437), .Y(n_420) );
NOR2xp33_ASAP7_75t_SL g421 ( .A(n_422), .B(n_426), .Y(n_421) );
INVxp67_ASAP7_75t_L g454 ( .A(n_422), .Y(n_454) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g479 ( .A(n_424), .Y(n_479) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .C(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g441 ( .A(n_435), .Y(n_441) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g450 ( .A(n_438), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_443), .A2(n_494), .B1(n_495), .B2(n_498), .C(n_499), .Y(n_493) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI32xp33_ASAP7_75t_L g449 ( .A1(n_446), .A2(n_450), .A3(n_451), .B1(n_452), .B2(n_454), .Y(n_449) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_452), .A2(n_462), .B1(n_463), .B2(n_464), .C(n_470), .Y(n_461) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_474), .C(n_492), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B(n_461), .Y(n_456) );
AOI211x1_ASAP7_75t_L g474 ( .A1(n_457), .A2(n_475), .B(n_477), .C(n_484), .Y(n_474) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2x1_ASAP7_75t_SL g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g476 ( .A(n_467), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AO21x1_ASAP7_75t_L g484 ( .A1(n_473), .A2(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g518 ( .A(n_489), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_505), .Y(n_492) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI21xp33_ASAP7_75t_SL g499 ( .A1(n_500), .A2(n_501), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_509), .Y(n_506) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g515 ( .A(n_514), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_523), .A2(n_530), .B(n_842), .C(n_852), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_523), .A2(n_843), .B(n_844), .Y(n_842) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g843 ( .A(n_532), .Y(n_843) );
NAND4xp75_ASAP7_75t_L g532 ( .A(n_533), .B(n_682), .C(n_758), .D(n_810), .Y(n_532) );
AND3x1_ASAP7_75t_L g533 ( .A(n_534), .B(n_655), .C(n_668), .Y(n_533) );
AOI221x1_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_587), .B1(n_616), .B2(n_620), .C(n_632), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_535), .A2(n_656), .B(n_658), .C(n_659), .Y(n_655) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_550), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g619 ( .A(n_539), .Y(n_619) );
BUFx2_ASAP7_75t_L g637 ( .A(n_539), .Y(n_637) );
OR2x2_ASAP7_75t_L g679 ( .A(n_539), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g686 ( .A(n_539), .B(n_553), .Y(n_686) );
AND2x4_ASAP7_75t_L g721 ( .A(n_539), .B(n_552), .Y(n_721) );
OR2x2_ASAP7_75t_L g764 ( .A(n_539), .B(n_580), .Y(n_764) );
AO31x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .A3(n_546), .B(n_548), .Y(n_539) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_546), .A2(n_609), .A3(n_610), .B(n_614), .Y(n_608) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_SL g577 ( .A(n_547), .Y(n_577) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_565), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_552), .B(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_552), .Y(n_651) );
INVx2_ASAP7_75t_L g678 ( .A(n_552), .Y(n_678) );
INVx3_ASAP7_75t_L g691 ( .A(n_552), .Y(n_691) );
AND2x2_ASAP7_75t_L g809 ( .A(n_552), .B(n_638), .Y(n_809) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g618 ( .A(n_553), .B(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g674 ( .A(n_553), .Y(n_674) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .A3(n_562), .B(n_563), .Y(n_553) );
AO31x2_ASAP7_75t_L g625 ( .A1(n_562), .A2(n_609), .A3(n_626), .B(n_629), .Y(n_625) );
INVxp67_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g694 ( .A(n_566), .Y(n_694) );
INVx1_ASAP7_75t_L g821 ( .A(n_566), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_579), .Y(n_566) );
AND2x2_ASAP7_75t_L g617 ( .A(n_567), .B(n_580), .Y(n_617) );
INVx1_ASAP7_75t_L g680 ( .A(n_567), .Y(n_680) );
OAI21x1_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_578), .Y(n_567) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_568), .A2(n_569), .B(n_578), .Y(n_639) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .B(n_577), .Y(n_569) );
INVx2_ASAP7_75t_L g635 ( .A(n_579), .Y(n_635) );
AND2x2_ASAP7_75t_L g687 ( .A(n_579), .B(n_638), .Y(n_687) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g649 ( .A(n_580), .Y(n_649) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_580), .Y(n_709) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_589), .A2(n_681), .B1(n_685), .B2(n_688), .Y(n_684) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_598), .Y(n_589) );
INVx1_ASAP7_75t_L g702 ( .A(n_590), .Y(n_702) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g622 ( .A(n_591), .B(n_600), .Y(n_622) );
AND2x2_ASAP7_75t_L g653 ( .A(n_591), .B(n_608), .Y(n_653) );
INVx4_ASAP7_75t_SL g664 ( .A(n_591), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_591), .B(n_698), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_591), .B(n_837), .Y(n_836) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g735 ( .A(n_599), .B(n_713), .Y(n_735) );
OR2x2_ASAP7_75t_L g768 ( .A(n_599), .B(n_750), .Y(n_768) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_608), .Y(n_599) );
INVx2_ASAP7_75t_L g642 ( .A(n_600), .Y(n_642) );
INVx1_ASAP7_75t_L g647 ( .A(n_600), .Y(n_647) );
AND2x2_ASAP7_75t_L g654 ( .A(n_600), .B(n_624), .Y(n_654) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_600), .Y(n_670) );
INVx1_ASAP7_75t_L g698 ( .A(n_600), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_600), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g631 ( .A(n_608), .Y(n_631) );
AND2x4_ASAP7_75t_L g641 ( .A(n_608), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g667 ( .A(n_608), .Y(n_667) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_608), .Y(n_744) );
INVx1_ASAP7_75t_L g837 ( .A(n_608), .Y(n_837) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_617), .B(n_690), .Y(n_757) );
AND2x2_ASAP7_75t_L g770 ( .A(n_617), .B(n_686), .Y(n_770) );
AND2x2_ASAP7_75t_L g840 ( .A(n_617), .B(n_691), .Y(n_840) );
AND2x4_ASAP7_75t_L g675 ( .A(n_619), .B(n_638), .Y(n_675) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g742 ( .A(n_622), .B(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g756 ( .A(n_622), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_622), .B(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_623), .B(n_696), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_623), .A2(n_753), .B(n_756), .C(n_757), .Y(n_752) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_631), .Y(n_623) );
AND2x2_ASAP7_75t_L g723 ( .A(n_624), .B(n_664), .Y(n_723) );
INVx3_ASAP7_75t_L g750 ( .A(n_624), .Y(n_750) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g645 ( .A(n_625), .Y(n_645) );
AND2x4_ASAP7_75t_L g671 ( .A(n_625), .B(n_631), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_631), .B(n_664), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_640), .B1(n_648), .B2(n_652), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g789 ( .A(n_634), .Y(n_789) );
AND2x4_ASAP7_75t_L g700 ( .A(n_635), .B(n_680), .Y(n_700) );
INVx1_ASAP7_75t_L g720 ( .A(n_635), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_637), .A2(n_693), .B1(n_703), .B2(n_705), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_637), .B(n_694), .Y(n_751) );
NAND2x1_ASAP7_75t_L g808 ( .A(n_637), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g823 ( .A(n_637), .Y(n_823) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g762 ( .A(n_639), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
AND2x2_ASAP7_75t_L g681 ( .A(n_641), .B(n_663), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_641), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g722 ( .A(n_641), .B(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_641), .Y(n_796) );
NAND2x1p5_ASAP7_75t_L g803 ( .A(n_641), .B(n_704), .Y(n_803) );
AND2x4_ASAP7_75t_L g826 ( .A(n_641), .B(n_754), .Y(n_826) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx3_ASAP7_75t_L g704 ( .A(n_644), .Y(n_704) );
AND2x2_ASAP7_75t_L g716 ( .A(n_644), .B(n_709), .Y(n_716) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g666 ( .A(n_645), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g714 ( .A(n_645), .Y(n_714) );
INVx1_ASAP7_75t_L g657 ( .A(n_646), .Y(n_657) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g814 ( .A(n_647), .B(n_664), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
AND2x2_ASAP7_75t_L g740 ( .A(n_649), .B(n_721), .Y(n_740) );
INVx2_ASAP7_75t_L g781 ( .A(n_649), .Y(n_781) );
AND2x4_ASAP7_75t_L g782 ( .A(n_649), .B(n_675), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_650), .B(n_700), .Y(n_830) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_653), .B(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g725 ( .A(n_653), .B(n_670), .Y(n_725) );
INVx1_ASAP7_75t_L g817 ( .A(n_653), .Y(n_817) );
AND2x2_ASAP7_75t_L g816 ( .A(n_654), .B(n_743), .Y(n_816) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_658), .A2(n_788), .B1(n_790), .B2(n_792), .Y(n_787) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g696 ( .A(n_664), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g732 ( .A(n_664), .Y(n_732) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_664), .Y(n_738) );
INVx2_ASAP7_75t_L g755 ( .A(n_664), .Y(n_755) );
OR2x2_ASAP7_75t_L g776 ( .A(n_664), .B(n_739), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_664), .B(n_734), .Y(n_786) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g753 ( .A(n_666), .B(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_666), .Y(n_807) );
INVx1_ASAP7_75t_L g734 ( .A(n_667), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B(n_676), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_671), .B(n_702), .Y(n_701) );
INVx3_ASAP7_75t_L g739 ( .A(n_671), .Y(n_739) );
AND2x2_ASAP7_75t_L g813 ( .A(n_671), .B(n_814), .Y(n_813) );
AOI211x1_ASAP7_75t_SL g741 ( .A1(n_672), .A2(n_742), .B(n_745), .C(n_752), .Y(n_741) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g798 ( .A(n_674), .B(n_675), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_675), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_675), .Y(n_791) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g706 ( .A(n_678), .Y(n_706) );
NOR2x1p5_ASAP7_75t_L g763 ( .A(n_678), .B(n_764), .Y(n_763) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_679), .B(n_708), .Y(n_707) );
NOR2xp67_ASAP7_75t_SL g780 ( .A(n_679), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g841 ( .A(n_681), .B(n_749), .Y(n_841) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_726), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_684), .B(n_692), .C(n_710), .Y(n_683) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_686), .Y(n_717) );
AND2x2_ASAP7_75t_L g724 ( .A(n_686), .B(n_720), .Y(n_724) );
AND2x4_ASAP7_75t_SL g838 ( .A(n_686), .B(n_700), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_687), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_689), .A2(n_731), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x4_ASAP7_75t_L g820 ( .A(n_691), .B(n_821), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_699), .B2(n_701), .Y(n_693) );
NAND2x1_ASAP7_75t_L g769 ( .A(n_696), .B(n_749), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_696), .B(n_743), .Y(n_779) );
INVx1_ASAP7_75t_L g806 ( .A(n_696), .Y(n_806) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_699), .A2(n_825), .B(n_828), .Y(n_824) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_700), .A2(n_712), .B(n_715), .Y(n_711) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g785 ( .A(n_704), .Y(n_785) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g729 ( .A(n_707), .Y(n_729) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_717), .B1(n_718), .B2(n_722), .C1(n_724), .C2(n_725), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_712), .A2(n_746), .B(n_751), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_713), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g827 ( .A(n_713), .Y(n_827) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_714), .Y(n_833) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
AND2x2_ASAP7_75t_L g797 ( .A(n_719), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g790 ( .A(n_720), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_741), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B1(n_736), .B2(n_740), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVx1_ASAP7_75t_L g747 ( .A(n_733), .Y(n_747) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx4_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OR2x2_ASAP7_75t_L g775 ( .A(n_750), .B(n_767), .Y(n_775) );
OR2x2_ASAP7_75t_L g835 ( .A(n_750), .B(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND5xp2_ASAP7_75t_L g811 ( .A(n_756), .B(n_803), .C(n_812), .D(n_815), .E(n_817), .Y(n_811) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_794), .Y(n_758) );
NAND2xp67_ASAP7_75t_SL g759 ( .A(n_760), .B(n_777), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_765), .B1(n_770), .B2(n_771), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
NAND3xp33_ASAP7_75t_SL g765 ( .A(n_766), .B(n_768), .C(n_769), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g800 ( .A(n_769), .Y(n_800) );
NAND3xp33_ASAP7_75t_SL g771 ( .A(n_772), .B(n_775), .C(n_776), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g793 ( .A(n_774), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_SL g805 ( .A1(n_775), .A2(n_806), .B(n_807), .C(n_808), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .B1(n_782), .B2(n_783), .C(n_787), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_784), .B(n_832), .Y(n_831) );
OR2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g801 ( .A(n_788), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_799), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g804 ( .A(n_798), .Y(n_804) );
AOI211xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B(n_802), .C(n_805), .Y(n_799) );
AOI211x1_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_818), .B(n_824), .C(n_839), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2x1p5_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NAND2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_831), .B1(n_834), .B2(n_838), .Y(n_828) );
INVxp67_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g852 ( .A(n_844), .B(n_853), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx5_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
BUFx10_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_860), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx8_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_885), .Y(n_860) );
AOI31xp33_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_873), .A3(n_874), .B(n_879), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_862), .B(n_887), .Y(n_886) );
AO22x1_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_865), .B1(n_871), .B2(n_872), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_863), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_865), .Y(n_872) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx2_ASAP7_75t_L g888 ( .A(n_873), .Y(n_888) );
INVx1_ASAP7_75t_L g887 ( .A(n_874), .Y(n_887) );
BUFx2_ASAP7_75t_SL g874 ( .A(n_875), .Y(n_874) );
INVx4_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g883 ( .A(n_878), .Y(n_883) );
NOR2xp33_ASAP7_75t_SL g879 ( .A(n_880), .B(n_884), .Y(n_879) );
INVx5_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_888), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
CKINVDCx16_ASAP7_75t_R g891 ( .A(n_892), .Y(n_891) );
endmodule