module real_jpeg_4027_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_89),
.B(n_92),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_1),
.B(n_228),
.C(n_231),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_1),
.A2(n_61),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_1),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_1),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_1),
.A2(n_131),
.B1(n_286),
.B2(n_294),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_2),
.A2(n_63),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_2),
.A2(n_63),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_3),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_141),
.B1(n_208),
.B2(n_211),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_29),
.B1(n_115),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_4),
.A2(n_29),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_4),
.A2(n_29),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_61),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_86),
.B1(n_132),
.B2(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_8),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_12),
.A2(n_56),
.B1(n_133),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_12),
.A2(n_56),
.B1(n_240),
.B2(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_14),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_14),
.A2(n_114),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_14),
.A2(n_114),
.B1(n_237),
.B2(n_240),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_14),
.A2(n_114),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_216),
.B1(n_217),
.B2(n_349),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_18),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_214),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_179),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_20),
.B(n_179),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_118),
.C(n_157),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_21),
.B(n_347),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_21),
.Y(n_350)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_59),
.CI(n_87),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_22),
.B(n_59),
.C(n_87),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B1(n_32),
.B2(n_50),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_23),
.A2(n_30),
.B1(n_32),
.B2(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_24),
.B(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_27),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_27),
.Y(n_323)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_31),
.A2(n_51),
.B(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_31),
.A2(n_174),
.B1(n_247),
.B2(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_41),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_32),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_32),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_32)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_33),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_33),
.Y(n_235)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_35),
.Y(n_317)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_37),
.Y(n_311)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_39),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_39),
.Y(n_239)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_39),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_39),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g306 ( 
.A1(n_57),
.A2(n_307),
.A3(n_309),
.B1(n_312),
.B2(n_316),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_58),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_66),
.B(n_81),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_60),
.B(n_212),
.Y(n_340)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_64),
.Y(n_318)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_66),
.A2(n_206),
.B1(n_207),
.B2(n_212),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_66),
.A2(n_338),
.B(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_67),
.A2(n_82),
.B1(n_233),
.B2(n_236),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_67),
.A2(n_82),
.B1(n_236),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_67),
.A2(n_82),
.B1(n_249),
.B2(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_69),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_75),
.Y(n_231)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_80),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_83),
.Y(n_206)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B1(n_109),
.B2(n_117),
.Y(n_87)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_95),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_110),
.A2(n_171),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_120),
.A3(n_123),
.B1(n_125),
.B2(n_129),
.Y(n_119)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_117),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_118),
.B(n_157),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_130),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_130),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_138),
.B1(n_146),
.B2(n_150),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_131),
.A2(n_150),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_131),
.A2(n_257),
.B(n_259),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_131),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_131),
.A2(n_202),
.B1(n_274),
.B2(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_131),
.A2(n_200),
.B(n_261),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_137),
.Y(n_298)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_160),
.B(n_164),
.Y(n_159)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_143),
.Y(n_258)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_145),
.Y(n_267)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_154),
.Y(n_275)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.C(n_172),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_158),
.A2(n_159),
.B1(n_169),
.B2(n_170),
.Y(n_333)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_172),
.B(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_197),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_213),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_208),
.Y(n_326)
);

INVx5_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_212),
.B(n_234),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_344),
.B(n_348),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_328),
.B(n_343),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_302),
.B(n_327),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_270),
.B(n_301),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_243),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_222),
.B(n_243),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_232),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_234),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_234),
.B(n_313),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_234),
.A2(n_312),
.B(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_256),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_255),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_255),
.C(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_248),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_268),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_282),
.B(n_300),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_281),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_281),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_292),
.B(n_299),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_304),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_320),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_321),
.C(n_324),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_319),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_329),
.B(n_330),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_337),
.C(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_341),
.B2(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_346),
.Y(n_348)
);


endmodule