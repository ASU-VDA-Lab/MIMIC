module fake_jpeg_54_n_606 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_606);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_606;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_58),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_59),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_186)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_61),
.B(n_80),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_63),
.Y(n_194)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_66),
.Y(n_182)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_70),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_27),
.B(n_18),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_8),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_89),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_27),
.B(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_25),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_94),
.B(n_96),
.Y(n_173)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_37),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_97),
.Y(n_213)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_23),
.B(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_99),
.B(n_113),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_112),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_22),
.B(n_7),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_125),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_43),
.B(n_46),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_23),
.B(n_7),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_30),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_52),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_55),
.Y(n_133)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_127),
.B(n_1),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_133),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_44),
.B1(n_51),
.B2(n_34),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_135),
.A2(n_159),
.B1(n_168),
.B2(n_196),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_43),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_137),
.B(n_148),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_48),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_48),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_151),
.B(n_58),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_46),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_156),
.B(n_166),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_69),
.A2(n_51),
.B1(n_44),
.B2(n_34),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_45),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_100),
.A2(n_45),
.B1(n_42),
.B2(n_55),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_60),
.Y(n_172)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_72),
.B(n_42),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_183),
.B(n_184),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_93),
.B(n_36),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_189),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_186),
.A2(n_191),
.B1(n_214),
.B2(n_134),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_91),
.B(n_9),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_62),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_191)
);

HAxp5_ASAP7_75t_SL g192 ( 
.A(n_70),
.B(n_16),
.CON(n_192),
.SN(n_192)
);

OR2x2_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_58),
.Y(n_224)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_107),
.A2(n_110),
.B1(n_119),
.B2(n_114),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_197),
.A2(n_202),
.B1(n_196),
.B2(n_135),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_69),
.A2(n_16),
.B1(n_13),
.B2(n_11),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_63),
.B(n_10),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_206),
.B(n_211),
.Y(n_284)
);

NAND2x1_ASAP7_75t_L g207 ( 
.A(n_125),
.B(n_11),
.Y(n_207)
);

NAND2x1_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_1),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_77),
.B(n_11),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_1),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_71),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_77),
.B(n_11),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_218),
.B(n_182),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_129),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_219),
.B(n_221),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_223),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_224),
.A2(n_242),
.B(n_247),
.Y(n_345)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_225),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_168),
.B1(n_83),
.B2(n_97),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_226),
.A2(n_255),
.B1(n_256),
.B2(n_278),
.Y(n_336)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_227),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_131),
.A2(n_85),
.B1(n_90),
.B2(n_74),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_228),
.Y(n_326)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_230),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_233),
.B(n_244),
.Y(n_304)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_234),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_197),
.A2(n_88),
.B1(n_81),
.B2(n_79),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_235),
.A2(n_243),
.B1(n_139),
.B2(n_239),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_237),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_238),
.B(n_240),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_239),
.B(n_263),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_73),
.Y(n_240)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_131),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_152),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_246),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_155),
.B(n_4),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_145),
.B(n_4),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_266),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_149),
.Y(n_252)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_254),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_164),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_169),
.A2(n_5),
.B1(n_205),
.B2(n_175),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_5),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_264),
.Y(n_307)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_207),
.A2(n_159),
.B(n_212),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_261),
.A2(n_247),
.B(n_295),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_134),
.Y(n_262)
);

INVx13_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_155),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_153),
.B(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_128),
.B(n_132),
.Y(n_266)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_158),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_270),
.Y(n_328)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_193),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_271),
.B(n_272),
.Y(n_340)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_210),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_182),
.B(n_152),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_274),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_215),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_276),
.Y(n_323)
);

BUFx4f_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_282),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_136),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_286),
.Y(n_311)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_285),
.A2(n_287),
.B1(n_289),
.B2(n_291),
.Y(n_346)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_143),
.A2(n_144),
.B1(n_204),
.B2(n_157),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_253),
.B1(n_267),
.B2(n_223),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_177),
.A2(n_188),
.B1(n_201),
.B2(n_198),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_180),
.B(n_143),
.C(n_140),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_140),
.C(n_144),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_154),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_154),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_157),
.Y(n_293)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_167),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_295),
.Y(n_324)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_161),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_309),
.B1(n_332),
.B2(n_335),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_278),
.A2(n_261),
.B1(n_273),
.B2(n_284),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_250),
.A2(n_162),
.B1(n_213),
.B2(n_204),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_313),
.B1(n_320),
.B2(n_351),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_312),
.B(n_319),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_235),
.A2(n_192),
.B1(n_174),
.B2(n_142),
.Y(n_313)
);

OAI22x1_ASAP7_75t_L g317 ( 
.A1(n_224),
.A2(n_136),
.B1(n_142),
.B2(n_163),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_SL g376 ( 
.A1(n_317),
.A2(n_316),
.B(n_324),
.Y(n_376)
);

NAND2x1_ASAP7_75t_L g319 ( 
.A(n_242),
.B(n_163),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_275),
.A2(n_174),
.B1(n_208),
.B2(n_202),
.Y(n_320)
);

AO22x1_ASAP7_75t_SL g329 ( 
.A1(n_243),
.A2(n_139),
.B1(n_208),
.B2(n_239),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_349),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_139),
.B1(n_275),
.B2(n_265),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_249),
.B(n_251),
.C(n_266),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_339),
.C(n_348),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g339 ( 
.A(n_257),
.B(n_247),
.C(n_290),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_342),
.A2(n_326),
.B(n_319),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_282),
.A2(n_260),
.B1(n_268),
.B2(n_271),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_281),
.B1(n_241),
.B2(n_285),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_SL g348 ( 
.A(n_231),
.B(n_248),
.C(n_232),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_225),
.B(n_280),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_227),
.B(n_286),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_347),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_277),
.A2(n_220),
.B1(n_259),
.B2(n_272),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_237),
.B(n_283),
.C(n_245),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_352),
.B(n_263),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_335),
.A2(n_252),
.B1(n_229),
.B2(n_277),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_353),
.A2(n_368),
.B1(n_371),
.B2(n_376),
.Y(n_398)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_358),
.Y(n_417)
);

AOI22x1_ASAP7_75t_SL g360 ( 
.A1(n_309),
.A2(n_246),
.B1(n_292),
.B2(n_230),
.Y(n_360)
);

OA22x2_ASAP7_75t_L g418 ( 
.A1(n_360),
.A2(n_362),
.B1(n_370),
.B2(n_378),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_361),
.B(n_374),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_222),
.B1(n_234),
.B2(n_291),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_349),
.Y(n_363)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_236),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_375),
.Y(n_404)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_315),
.Y(n_367)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_342),
.A2(n_294),
.B1(n_317),
.B2(n_298),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_369),
.A2(n_377),
.B(n_391),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_326),
.A2(n_344),
.B1(n_303),
.B2(n_332),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_298),
.A2(n_345),
.B1(n_308),
.B2(n_329),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_304),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_372),
.B(n_381),
.Y(n_410)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_340),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_319),
.A2(n_346),
.B(n_324),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_300),
.A2(n_323),
.B1(n_329),
.B2(n_339),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_380),
.Y(n_402)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_314),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_386),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_316),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_385),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_312),
.A2(n_307),
.B1(n_316),
.B2(n_338),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_394),
.B1(n_376),
.B2(n_383),
.Y(n_409)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_300),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_325),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_388),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_306),
.B(n_333),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_306),
.B(n_352),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_390),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_334),
.B(n_305),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_346),
.A2(n_301),
.B1(n_302),
.B2(n_299),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_392),
.B(n_393),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_327),
.A2(n_331),
.B1(n_318),
.B2(n_321),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_343),
.B(n_302),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_396),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_331),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_395),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_412),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_377),
.A2(n_325),
.B(n_297),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_400),
.A2(n_357),
.B(n_391),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_297),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_403),
.B(n_408),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

INVx8_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_301),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_387),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_322),
.C(n_299),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_429),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_359),
.A2(n_327),
.B1(n_318),
.B2(n_341),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_414),
.A2(n_362),
.B1(n_381),
.B2(n_380),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_322),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_426),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_337),
.Y(n_425)
);

XNOR2x1_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_430),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_378),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_379),
.B(n_341),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_337),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_341),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_415),
.A2(n_369),
.B(n_377),
.Y(n_434)
);

AO21x1_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_463),
.B(n_448),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_365),
.Y(n_436)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

OA22x2_ASAP7_75t_L g437 ( 
.A1(n_398),
.A2(n_368),
.B1(n_370),
.B2(n_354),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_437),
.B(n_466),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_359),
.B1(n_354),
.B2(n_371),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_439),
.A2(n_440),
.B1(n_448),
.B2(n_454),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_409),
.A2(n_373),
.B1(n_367),
.B2(n_363),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_402),
.Y(n_441)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_443),
.A2(n_456),
.B1(n_458),
.B2(n_464),
.Y(n_481)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_419),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_445),
.B(n_447),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_406),
.A2(n_360),
.B1(n_358),
.B2(n_356),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_446),
.A2(n_459),
.B1(n_461),
.B2(n_423),
.Y(n_468)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_406),
.A2(n_355),
.B1(n_353),
.B2(n_389),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_419),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_449),
.B(n_455),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_453),
.A2(n_415),
.B(n_400),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_432),
.A2(n_433),
.B1(n_421),
.B2(n_417),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_428),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_411),
.A2(n_375),
.B1(n_360),
.B2(n_374),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_411),
.A2(n_372),
.B1(n_364),
.B2(n_355),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_421),
.B1(n_401),
.B2(n_404),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_396),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_460),
.B(n_407),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_404),
.A2(n_388),
.B1(n_390),
.B2(n_382),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_422),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_462),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_426),
.B(n_394),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_424),
.A2(n_366),
.B1(n_385),
.B2(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_431),
.Y(n_469)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_471),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_472),
.A2(n_483),
.B(n_487),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_405),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_475),
.B(n_477),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_424),
.B1(n_420),
.B2(n_423),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_476),
.A2(n_441),
.B1(n_444),
.B2(n_447),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_410),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_416),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_478),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_430),
.B1(n_425),
.B2(n_429),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_446),
.B1(n_464),
.B2(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_434),
.A2(n_418),
.B(n_403),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_413),
.C(n_408),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_486),
.C(n_488),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_418),
.C(n_442),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_453),
.A2(n_418),
.B(n_449),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_442),
.B(n_418),
.C(n_438),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_445),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_489),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_456),
.B(n_436),
.Y(n_490)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_490),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_438),
.B(n_451),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_485),
.Y(n_508)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_451),
.B(n_439),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_492),
.B(n_437),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_450),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_493),
.B(n_497),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_459),
.C(n_466),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_450),
.C(n_454),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_503),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_501),
.B(n_508),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_507),
.A2(n_467),
.B1(n_494),
.B2(n_474),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_488),
.C(n_491),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_514),
.C(n_520),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_437),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_515),
.Y(n_539)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_512),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_437),
.C(n_463),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_437),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_487),
.A2(n_463),
.B(n_443),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g530 ( 
.A(n_516),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_468),
.B(n_435),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_519),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_435),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_479),
.B(n_469),
.C(n_493),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_473),
.B(n_470),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_522),
.B(n_523),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_498),
.A2(n_481),
.B1(n_490),
.B2(n_467),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_524),
.A2(n_527),
.B1(n_507),
.B2(n_516),
.Y(n_548)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_525),
.Y(n_547)
);

FAx1_ASAP7_75t_SL g526 ( 
.A(n_520),
.B(n_495),
.CI(n_469),
.CON(n_526),
.SN(n_526)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_537),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_498),
.A2(n_481),
.B1(n_467),
.B2(n_489),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_506),
.Y(n_529)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_529),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_513),
.A2(n_473),
.B1(n_470),
.B2(n_495),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_532),
.A2(n_543),
.B1(n_512),
.B2(n_509),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_508),
.B(n_505),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_503),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_502),
.B(n_482),
.C(n_484),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_535),
.B(n_538),
.C(n_540),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_523),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_502),
.B(n_482),
.C(n_484),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_474),
.C(n_472),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_542),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_545),
.A2(n_548),
.B1(n_559),
.B2(n_500),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_546),
.A2(n_554),
.B(n_557),
.Y(n_560)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_535),
.Y(n_549)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_515),
.C(n_519),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_550),
.B(n_552),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_521),
.C(n_518),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_530),
.A2(n_499),
.B(n_497),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_514),
.C(n_517),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_556),
.B(n_558),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_536),
.A2(n_499),
.B(n_497),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_501),
.C(n_505),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_529),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_544),
.B(n_552),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_561),
.B(n_562),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_534),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_539),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_566),
.Y(n_578)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_565),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_558),
.B(n_539),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_556),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_567),
.B(n_570),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_557),
.A2(n_509),
.B(n_511),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_554),
.B(n_531),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_572),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_531),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_524),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_573),
.B(n_547),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_576),
.Y(n_588)
);

AOI21x1_ASAP7_75t_L g576 ( 
.A1(n_560),
.A2(n_564),
.B(n_559),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_561),
.B(n_541),
.C(n_527),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_579),
.B(n_580),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_568),
.B(n_572),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_570),
.A2(n_525),
.B1(n_551),
.B2(n_555),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_583),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_569),
.A2(n_526),
.B1(n_551),
.B2(n_541),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_582),
.B(n_555),
.Y(n_585)
);

AOI21xp33_ASAP7_75t_L g595 ( 
.A1(n_585),
.A2(n_591),
.B(n_480),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_563),
.C(n_566),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_587),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_562),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_589),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_574),
.B(n_504),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_578),
.B(n_579),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_592),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g594 ( 
.A1(n_585),
.A2(n_583),
.B(n_586),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_595),
.Y(n_599)
);

OA21x2_ASAP7_75t_L g598 ( 
.A1(n_593),
.A2(n_588),
.B(n_576),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_598),
.A2(n_586),
.B1(n_596),
.B2(n_581),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_597),
.B(n_590),
.C(n_578),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_600),
.B(n_504),
.C(n_528),
.Y(n_602)
);

OAI321xp33_ASAP7_75t_L g603 ( 
.A1(n_601),
.A2(n_602),
.A3(n_599),
.B1(n_526),
.B2(n_528),
.C(n_471),
.Y(n_603)
);

BUFx24_ASAP7_75t_SL g604 ( 
.A(n_603),
.Y(n_604)
);

FAx1_ASAP7_75t_SL g605 ( 
.A(n_604),
.B(n_471),
.CI(n_603),
.CON(n_605),
.SN(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_605),
.B(n_471),
.Y(n_606)
);


endmodule