module fake_jpeg_22980_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_35),
.B(n_39),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_45),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_31),
.Y(n_51)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_36),
.B1(n_19),
.B2(n_16),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_66),
.B(n_38),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_56),
.Y(n_88)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI222xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_18),
.B1(n_16),
.B2(n_22),
.C1(n_25),
.C2(n_19),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_23),
.C(n_31),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_1),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_44),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_44),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_89),
.C(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_80),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_38),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_87),
.B(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_81),
.B1(n_64),
.B2(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_26),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_44),
.B(n_45),
.Y(n_87)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_15),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_52),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_43),
.B1(n_40),
.B2(n_34),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_64),
.B1(n_47),
.B2(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_1),
.Y(n_124)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_34),
.B1(n_19),
.B2(n_17),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_111),
.B1(n_100),
.B2(n_99),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_54),
.B1(n_64),
.B2(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_119),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_121),
.B1(n_125),
.B2(n_128),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_68),
.B(n_62),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_91),
.B(n_92),
.C(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_122),
.Y(n_131)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_2),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_76),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_50),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_79),
.A2(n_95),
.B1(n_74),
.B2(n_88),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_40),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_33),
.B1(n_32),
.B2(n_40),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_135),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_74),
.B1(n_97),
.B2(n_72),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_137),
.B1(n_139),
.B2(n_147),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_148),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_97),
.B1(n_99),
.B2(n_91),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_97),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_103),
.B(n_118),
.Y(n_158)
);

XOR2x2_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_120),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_149),
.Y(n_159)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_150),
.Y(n_163)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_119),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_86),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_102),
.B(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_164),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_106),
.C(n_116),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_148),
.C(n_139),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_161),
.B(n_137),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_103),
.B1(n_121),
.B2(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_114),
.B(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_109),
.B1(n_128),
.B2(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_2),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_146),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_137),
.B(n_140),
.C(n_149),
.D(n_134),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_175),
.C(n_179),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_158),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_133),
.C(n_131),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_131),
.C(n_129),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_181),
.B(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_149),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_155),
.B1(n_163),
.B2(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_191),
.B(n_180),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_163),
.B1(n_140),
.B2(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_175),
.Y(n_195)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_2),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_179),
.C(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_161),
.B1(n_143),
.B2(n_9),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_181),
.B(n_168),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_196),
.B(n_199),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_188),
.B1(n_183),
.B2(n_190),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_188),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_191),
.A2(n_173),
.B(n_14),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_9),
.B(n_11),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_4),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_205),
.C(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_189),
.B(n_187),
.C(n_6),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_210),
.B(n_202),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_198),
.B(n_5),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_207),
.B(n_202),
.C(n_6),
.Y(n_212)
);

AO21x2_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_214),
.B(n_4),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_7),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_5),
.C(n_6),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_7),
.Y(n_220)
);


endmodule