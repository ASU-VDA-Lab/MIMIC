module real_jpeg_32390_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_288;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_105;
wire n_40;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_238;
wire n_67;
wire n_76;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_295;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_206;
wire n_53;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_181;
wire n_102;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_0),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_0),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_34),
.B1(n_94),
.B2(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_3),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_4),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_4),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_4),
.A2(n_111),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_4),
.A2(n_111),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_132),
.B1(n_135),
.B2(n_139),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_139),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_5),
.A2(n_139),
.B1(n_254),
.B2(n_259),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_6),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_6),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_6),
.A2(n_90),
.B1(n_231),
.B2(n_236),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_8),
.A2(n_50),
.A3(n_59),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_8),
.A2(n_51),
.B1(n_118),
.B2(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_8),
.B(n_122),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_8),
.A2(n_25),
.B1(n_253),
.B2(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_11),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_12),
.Y(n_120)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_13),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_13),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_190),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_189),
.Y(n_15)
);

INVxp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_168),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_18),
.B(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_107),
.B2(n_108),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_72),
.B1(n_105),
.B2(n_106),
.Y(n_20)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_22),
.A2(n_23),
.B1(n_49),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_37),
.B2(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_24),
.A2(n_40),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_24),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_282)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_25),
.A2(n_230),
.B1(n_238),
.B2(n_242),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_25),
.A2(n_253),
.B1(n_262),
.B2(n_267),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_30),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_30),
.Y(n_237)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_30),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_33),
.Y(n_226)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_39),
.Y(n_151)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_39),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_44),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_59),
.B(n_66),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_67),
.C(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_51),
.B(n_160),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_51),
.A2(n_197),
.B(n_200),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_51),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_51),
.B(n_97),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_51),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_58),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_59),
.A2(n_124),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_71),
.Y(n_212)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_88),
.B1(n_97),
.B2(n_99),
.Y(n_72)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_73),
.A2(n_97),
.B1(n_176),
.B2(n_246),
.Y(n_245)
);

AO21x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_80),
.B(n_84),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_85),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_89),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_97),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_147),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_121),
.B1(n_131),
.B2(n_140),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_124)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_131),
.A2(n_140),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_158),
.B2(n_159),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.C(n_183),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_169),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_174),
.B(n_184),
.Y(n_294)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_196),
.B1(n_205),
.B2(n_213),
.Y(n_195)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_291),
.B(n_295),
.Y(n_190)
);

OAI21x1_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_249),
.B(n_290),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_228),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_193),
.B(n_228),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_214),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_194),
.A2(n_195),
.B1(n_214),
.B2(n_215),
.Y(n_288)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_223),
.B1(n_224),
.B2(n_227),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_243),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_245),
.C(n_247),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_281),
.B(n_289),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_269),
.B(n_280),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_268),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_268),
.Y(n_280)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_288),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);


endmodule