module real_jpeg_15535_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_173;
wire n_40;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_0),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_0),
.Y(n_149)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_3),
.A2(n_105),
.B1(n_108),
.B2(n_114),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_114),
.B1(n_169),
.B2(n_173),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_3),
.A2(n_114),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_4),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_5),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_53),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_58),
.B1(n_64),
.B2(n_68),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

OAI22x1_ASAP7_75t_L g178 ( 
.A1(n_6),
.A2(n_68),
.B1(n_179),
.B2(n_183),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_7),
.Y(n_142)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_7),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_7),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_8),
.Y(n_172)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_8),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_93),
.B1(n_98),
.B2(n_103),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_118),
.A3(n_123),
.B1(n_124),
.B2(n_127),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_9),
.B(n_71),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_9),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_9),
.B(n_175),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_11),
.Y(n_205)
);

XNOR2x2_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_192),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_191),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp67_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_166),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_16),
.B(n_166),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_69),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_34),
.B1(n_48),
.B2(n_57),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_20),
.A2(n_49),
.B1(n_168),
.B2(n_175),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_20),
.A2(n_168),
.B1(n_175),
.B2(n_218),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_24),
.Y(n_174)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_28),
.Y(n_215)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_32),
.Y(n_123)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_34),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_36),
.Y(n_258)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_43),
.Y(n_140)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_43),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_43),
.Y(n_165)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_43),
.Y(n_237)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_43),
.Y(n_250)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_92),
.B1(n_104),
.B2(n_115),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_103),
.B(n_212),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_103),
.A2(n_211),
.B(n_219),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_103),
.A2(n_138),
.B1(n_245),
.B2(n_248),
.Y(n_244)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

XOR2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_136),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_143),
.B(n_153),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_137),
.A2(n_228),
.B1(n_238),
.B2(n_239),
.Y(n_227)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_178),
.B(n_186),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_138),
.A2(n_229),
.B1(n_248),
.B2(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_142),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_SL g239 ( 
.A(n_156),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_176),
.C(n_177),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_176),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_225),
.B(n_266),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_223),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_194),
.B(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_216),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_216),
.B1(n_217),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_200),
.A3(n_206),
.B1(n_211),
.B2(n_213),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_242),
.B(n_265),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_240),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_240),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_259),
.B(n_264),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);


endmodule