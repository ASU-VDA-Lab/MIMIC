module real_jpeg_26039_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_1),
.A2(n_28),
.B1(n_56),
.B2(n_57),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_1),
.A2(n_54),
.B(n_165),
.C(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_55),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_57),
.B(n_75),
.C(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_1),
.B(n_22),
.C(n_36),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_1),
.B(n_73),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_1),
.B(n_87),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_1),
.B(n_38),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_43),
.B1(n_51),
.B2(n_130),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_40),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_52),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_105),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_105),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_105),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_134),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_132),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_106),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_106),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_83),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_62),
.B2(n_63),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_20),
.A2(n_29),
.B1(n_45),
.B2(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_20),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_20),
.A2(n_45),
.B1(n_189),
.B2(n_247),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_26),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_21),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_21),
.B(n_26),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_21),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_22),
.B(n_231),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_24),
.Y(n_168)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_28),
.A2(n_53),
.B(n_57),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_28),
.A2(n_37),
.B(n_77),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_29),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_30),
.A2(n_66),
.B(n_68),
.Y(n_146)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_31),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_31),
.B(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_31),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_33),
.A2(n_37),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_33),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_38),
.B(n_194),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_39),
.A2(n_68),
.B(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_41),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_41),
.B(n_193),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_59),
.B(n_60),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_49),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_49),
.B(n_61),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_55),
.B(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_57),
.B1(n_75),
.B2(n_77),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_82),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_65),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_70),
.B(n_204),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_78),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_81),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_79),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_125),
.Y(n_158)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_79),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.C(n_99),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_85),
.B(n_92),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_86),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_90),
.A2(n_116),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_90),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_99),
.B1(n_100),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_94),
.B(n_156),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_96),
.B(n_149),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_107),
.B(n_110),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_112),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_124),
.C(n_126),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_113),
.A2(n_114),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_122),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_118),
.B(n_217),
.Y(n_236)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_124),
.A2(n_126),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_124),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_126),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_270),
.B(n_274),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_182),
.B(n_256),
.C(n_269),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_170),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_137),
.B(n_170),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_153),
.B2(n_169),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_151),
.B2(n_152),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_140),
.B(n_152),
.C(n_169),
.Y(n_257)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_143),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_155),
.B(n_162),
.C(n_163),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.C(n_177),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_172),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_255),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_198),
.B(n_254),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_185),
.B(n_195),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_191),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_188),
.B(n_191),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_189),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_249),
.B(n_253),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_240),
.B(n_248),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_221),
.B(n_239),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_220),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_214),
.C(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_228),
.B(n_238),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_234),
.B(n_237),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_245),
.C(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_268),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_266),
.B2(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_267),
.C(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);


endmodule