module fake_jpeg_2962_n_354 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_1),
.B(n_2),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_42),
.A2(n_1),
.B(n_2),
.Y(n_106)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_45),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_8),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_36),
.Y(n_85)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_77),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_78),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_33),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_94),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_23),
.B1(n_36),
.B2(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_98),
.B1(n_117),
.B2(n_71),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_113),
.B1(n_114),
.B2(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_42),
.A2(n_29),
.B1(n_35),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_53),
.A2(n_58),
.B1(n_51),
.B2(n_56),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_102),
.A2(n_101),
.B1(n_86),
.B2(n_92),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_5),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_35),
.B1(n_65),
.B2(n_77),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_45),
.B1(n_37),
.B2(n_16),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_17),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_17),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_112),
.B(n_119),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_46),
.A2(n_35),
.B1(n_66),
.B2(n_69),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_40),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_34),
.B1(n_19),
.B2(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_19),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_34),
.B1(n_16),
.B2(n_24),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_31),
.B1(n_10),
.B2(n_13),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_52),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_4),
.Y(n_141)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_47),
.C(n_67),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_115),
.C(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_81),
.A2(n_127),
.B(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_131),
.B(n_134),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_45),
.B(n_43),
.C(n_49),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_133),
.A2(n_132),
.B(n_157),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_104),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_105),
.B1(n_92),
.B2(n_101),
.Y(n_175)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_142),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_47),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_144),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_11),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_145),
.A2(n_153),
.B(n_132),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

OR2x2_ASAP7_75t_SL g148 ( 
.A(n_97),
.B(n_37),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_12),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_107),
.A2(n_37),
.B1(n_16),
.B2(n_31),
.Y(n_150)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_85),
.B1(n_95),
.B2(n_122),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_82),
.A2(n_37),
.B1(n_16),
.B2(n_7),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_155),
.B1(n_156),
.B2(n_126),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_12),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_5),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_82),
.A2(n_16),
.B1(n_6),
.B2(n_9),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_165),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_164),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_95),
.B(n_6),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_6),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_87),
.Y(n_170)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_124),
.B(n_105),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_175),
.A2(n_180),
.B1(n_194),
.B2(n_197),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_207),
.B(n_138),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_9),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_190),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_184),
.A2(n_186),
.B1(n_196),
.B2(n_203),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_124),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_121),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_100),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_199),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_100),
.B1(n_109),
.B2(n_115),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_9),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_198),
.B(n_154),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_10),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_129),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_176),
.B(n_199),
.Y(n_237)
);

AND2x4_ASAP7_75t_SL g207 ( 
.A(n_146),
.B(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_222),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_237),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_128),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_145),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_217),
.Y(n_258)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_133),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_169),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_166),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_226),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_230),
.B(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_137),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_140),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_224),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_138),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_227),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_138),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_160),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_150),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_229),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_170),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_139),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_209),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_180),
.A2(n_136),
.B(n_155),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_186),
.B(n_195),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_234),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_188),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_196),
.B1(n_184),
.B2(n_202),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_207),
.B1(n_205),
.B2(n_178),
.Y(n_256)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_256),
.B1(n_229),
.B2(n_248),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_207),
.B1(n_182),
.B2(n_178),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_238),
.B1(n_228),
.B2(n_217),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_248),
.A2(n_264),
.B(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_195),
.B(n_188),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_207),
.C(n_178),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_212),
.C(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_181),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_235),
.B(n_221),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_212),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_270),
.C(n_271),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_213),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_214),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_241),
.B(n_222),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_225),
.B(n_226),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_277),
.A2(n_282),
.B(n_268),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_214),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_280),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_247),
.A2(n_246),
.B1(n_244),
.B2(n_261),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_281),
.A2(n_285),
.B1(n_230),
.B2(n_251),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_259),
.C(n_256),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_284),
.C(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_237),
.C(n_211),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_211),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_215),
.C(n_220),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_287),
.B(n_257),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_264),
.B1(n_263),
.B2(n_254),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_289),
.A2(n_304),
.B1(n_197),
.B2(n_240),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_283),
.C(n_270),
.Y(n_306)
);

XOR2x1_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_257),
.Y(n_293)
);

OAI321xp33_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_195),
.A3(n_231),
.B1(n_218),
.B2(n_183),
.C(n_266),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_249),
.B(n_219),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_296),
.B(n_298),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_243),
.B(n_221),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_210),
.B(n_223),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_262),
.B(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_300),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_269),
.C(n_271),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_308),
.C(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_284),
.C(n_287),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_278),
.C(n_234),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_318),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_281),
.B1(n_275),
.B2(n_286),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_311),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_245),
.B1(n_236),
.B2(n_252),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_296),
.A2(n_245),
.B1(n_252),
.B2(n_216),
.Y(n_316)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_289),
.A2(n_297),
.B1(n_295),
.B2(n_291),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_200),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_303),
.B1(n_293),
.B2(n_304),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_323),
.B1(n_319),
.B2(n_311),
.Y(n_335)
);

NOR2x1_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_206),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_299),
.B(n_297),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_329),
.B(n_310),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_291),
.B1(n_305),
.B2(n_292),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_326),
.C(n_327),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_302),
.C(n_305),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_240),
.C(n_181),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_332),
.A2(n_334),
.B1(n_336),
.B2(n_337),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_335),
.B(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

AOI321xp33_ASAP7_75t_L g336 ( 
.A1(n_324),
.A2(n_306),
.A3(n_314),
.B1(n_313),
.B2(n_317),
.C(n_316),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_325),
.A2(n_314),
.B1(n_315),
.B2(n_208),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_338),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_326),
.C(n_327),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_342),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_344),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_333),
.B(n_323),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_337),
.B(n_320),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_339),
.A2(n_322),
.B(n_206),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_343),
.C(n_341),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_348),
.A2(n_172),
.B1(n_204),
.B2(n_347),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_349),
.A2(n_350),
.B(n_345),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_204),
.C(n_172),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_172),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_353),
.B(n_204),
.Y(n_354)
);


endmodule