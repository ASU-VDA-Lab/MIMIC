module real_jpeg_6571_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_59),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_54),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_2),
.A2(n_54),
.B1(n_119),
.B2(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_2),
.A2(n_54),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_2),
.A2(n_222),
.B(n_225),
.C(n_228),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_2),
.B(n_84),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_42),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.C(n_266),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_2),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_2),
.B(n_260),
.C(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_2),
.B(n_93),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_27),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_3),
.A2(n_27),
.B1(n_99),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_3),
.A2(n_27),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_5),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_78),
.B1(n_161),
.B2(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_6),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_8),
.Y(n_102)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_8),
.Y(n_224)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_206),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_205),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_186),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_15),
.B(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_154),
.C(n_170),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_154),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_85),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_17),
.B(n_86),
.C(n_117),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_56),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_18),
.A2(n_19),
.B1(n_56),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_18),
.A2(n_19),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_18),
.A2(n_19),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_19),
.B(n_230),
.C(n_274),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_19),
.B(n_300),
.C(n_302),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B1(n_51),
.B2(n_52),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_21),
.B(n_42),
.Y(n_181)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_24),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_25),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_25),
.Y(n_199)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_26),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_26),
.Y(n_261)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_30),
.B(n_51),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_31),
.B(n_53),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_31),
.A2(n_42),
.B1(n_157),
.B2(n_197),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_42),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_37),
.Y(n_265)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_40),
.Y(n_159)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_42),
.A2(n_157),
.B(n_163),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_53),
.B(n_319),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_54),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_56),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_65),
.B1(n_73),
.B2(n_81),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_58),
.A2(n_82),
.B(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_62),
.Y(n_267)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_65),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_66),
.A2(n_176),
.B1(n_231),
.B2(n_234),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_66),
.A2(n_176),
.B1(n_231),
.B2(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_68),
.Y(n_233)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_72),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_74),
.B(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_77),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_116),
.B1(n_117),
.B2(n_153),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_86),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_86),
.B(n_200),
.C(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_86),
.A2(n_153),
.B1(n_200),
.B2(n_308),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_92),
.B1(n_111),
.B2(n_115),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_87),
.A2(n_92),
.B1(n_111),
.B2(n_115),
.Y(n_185)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_92),
.A2(n_111),
.B(n_115),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_95),
.Y(n_287)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_103)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_98),
.Y(n_226)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_104),
.Y(n_228)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_116),
.A2(n_117),
.B1(n_180),
.B2(n_258),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_116),
.B(n_258),
.C(n_282),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_116),
.A2(n_117),
.B1(n_318),
.B2(n_320),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_117),
.B(n_185),
.C(n_318),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_125),
.B1(n_140),
.B2(n_149),
.Y(n_117)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_118),
.A2(n_125),
.B1(n_140),
.B2(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_125),
.B(n_140),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_140),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_135),
.B2(n_137),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_136),
.Y(n_292)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_140),
.Y(n_275)
);

AOI22x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_165),
.B2(n_169),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_169),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_166),
.B(n_176),
.Y(n_293)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_182),
.C(n_185),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_173),
.A2(n_180),
.B1(n_258),
.B2(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_173),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_180),
.A2(n_258),
.B1(n_259),
.B2(n_268),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_180),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_185),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_185),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_185),
.A2(n_215),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_203),
.B2(n_204),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_194),
.B1(n_195),
.B2(n_202),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_200),
.B(n_201),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_200),
.Y(n_201)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_200),
.A2(n_304),
.B1(n_305),
.B2(n_308),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_200),
.Y(n_308)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_236),
.B(n_347),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_209),
.B(n_211),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.C(n_219),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_217),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_219),
.B(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_220),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_221),
.A2(n_229),
.B1(n_230),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_221),
.Y(n_326)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_229),
.A2(n_230),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_253),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_233),
.Y(n_246)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_328),
.B(n_344),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_312),
.B(n_327),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_297),
.B(n_311),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_279),
.B(n_296),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_270),
.B(n_278),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_255),
.B(n_269),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_252),
.B(n_254),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_248),
.A2(n_256),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_257),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_306),
.C(n_308),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_281),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_295),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_293),
.B2(n_294),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_294),
.Y(n_300)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_310),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_310),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_302),
.B1(n_303),
.B2(n_309),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_314),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_323),
.C(n_324),
.Y(n_337)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_338),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_337),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_336),
.C(n_340),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_338),
.A2(n_345),
.B(n_346),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_341),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);


endmodule