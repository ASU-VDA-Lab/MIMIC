module fake_ariane_1895_n_2463 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_387, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_381, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_389, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_382, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_393, n_359, n_155, n_127, n_2463);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_387;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_2463;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_1298;
wire n_737;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_645;
wire n_559;
wire n_2233;
wire n_2370;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_432;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_612;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_1833;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_1884;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_762;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_436;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_489;
wire n_2294;
wire n_2274;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_471;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_501;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1733;
wire n_1856;
wire n_463;
wire n_1524;
wire n_640;
wire n_1258;
wire n_2016;
wire n_1476;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_586;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_1659;
wire n_885;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1959;
wire n_1290;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_493;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_556;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_1663;
wire n_919;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_1720;
wire n_663;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_406;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_2372;
wire n_1533;
wire n_1806;
wire n_671;
wire n_1470;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1477;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_1591;
wire n_664;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_537;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_2081;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_2361;
wire n_1001;
wire n_1722;
wire n_1313;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_803;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_457;
wire n_2063;
wire n_1925;
wire n_782;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_284),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_145),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_170),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_308),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_162),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_93),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_176),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_321),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_187),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_262),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_120),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_70),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_302),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_280),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_256),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_283),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_388),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_189),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_108),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_317),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_296),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_288),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_268),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_304),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_61),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_92),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_378),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_5),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_88),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_6),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_56),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_300),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_244),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_285),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_356),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_100),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_193),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_67),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_29),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_278),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_88),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_117),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_365),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_19),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_113),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_358),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_326),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_167),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_58),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_99),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_312),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_393),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_260),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_293),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_359),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_92),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_258),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_367),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_250),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_137),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_384),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_135),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_7),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_214),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_17),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_154),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_93),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_7),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_153),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_267),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_279),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_325),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_112),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_179),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_352),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_218),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_332),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_224),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_328),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_166),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_381),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_175),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_299),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_112),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_281),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_131),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_94),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_90),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_220),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_118),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_341),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_121),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_197),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_313),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_183),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_140),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_10),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_12),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_368),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_232),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_307),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_38),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_54),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_226),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_178),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_297),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_215),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_257),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_166),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_319),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_24),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_354),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_336),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_180),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_316),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_301),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_298),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_331),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_111),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_94),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_31),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_294),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_150),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_152),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_343),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_338),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_119),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_123),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_122),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_286),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_177),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_391),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_222),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_208),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_202),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_122),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_238),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_188),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_383),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_104),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_355),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_18),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_109),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_305),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_17),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_182),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_75),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_69),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_27),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_13),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_234),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_67),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_324),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_246),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_75),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_361),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_113),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_128),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_241),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_357),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_273),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_375),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_134),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_231),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_30),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_309),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_185),
.Y(n_569)
);

BUFx8_ASAP7_75t_SL g570 ( 
.A(n_207),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_107),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_247),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_327),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_23),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_382),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_120),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_85),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_369),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_37),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_339),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_190),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_132),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_20),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_287),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_290),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_235),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_165),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_353),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_377),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_2),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_282),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_276),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_372),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_289),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_69),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_184),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_380),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_104),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_57),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_87),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_142),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_347),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_379),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_225),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_242),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_192),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_346),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_85),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_248),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_108),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_342),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_194),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_271),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_50),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_72),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_243),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_323),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_306),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_27),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_337),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_44),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_71),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_340),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_29),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_363),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_255),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_37),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_50),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_98),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_270),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_149),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_171),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_49),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_76),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_275),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_154),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_344),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_36),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_291),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_144),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_295),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_79),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_386),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_263),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_261),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_216),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_90),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_335),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_292),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_4),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_303),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_251),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_240),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_385),
.Y(n_654)
);

CKINVDCx14_ASAP7_75t_R g655 ( 
.A(n_371),
.Y(n_655)
);

CKINVDCx14_ASAP7_75t_R g656 ( 
.A(n_65),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_0),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_390),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_236),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_71),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_62),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_330),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_274),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_191),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_272),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_33),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_233),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_28),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_266),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_265),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_42),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_376),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_4),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_264),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_23),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_345),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_165),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_348),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_45),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_161),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_259),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_320),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_209),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_26),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_329),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_366),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_161),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_77),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_11),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_362),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_227),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_101),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_318),
.Y(n_693)
);

BUFx10_ASAP7_75t_L g694 ( 
.A(n_245),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_310),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_201),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_204),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_200),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_5),
.Y(n_699)
);

CKINVDCx16_ASAP7_75t_R g700 ( 
.A(n_143),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_35),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_22),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_252),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_315),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_22),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_72),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_34),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_11),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_14),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_21),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_81),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_374),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_206),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_81),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_42),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_364),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_351),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_389),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_210),
.Y(n_719)
);

CKINVDCx16_ASAP7_75t_R g720 ( 
.A(n_333),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_60),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_314),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_114),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_0),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_87),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_148),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_40),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_370),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_15),
.Y(n_729)
);

CKINVDCx16_ASAP7_75t_R g730 ( 
.A(n_322),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_84),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_91),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_153),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_91),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_269),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_148),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_157),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_350),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_277),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_146),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_467),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_441),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_441),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_587),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_587),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_600),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_467),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_600),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_406),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_715),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_715),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_724),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_480),
.B(n_1),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_570),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_724),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_397),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_407),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_450),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_456),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_463),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_467),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_467),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_487),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_488),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_413),
.B(n_1),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_492),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_503),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_504),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_521),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_700),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_531),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_538),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_689),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_467),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_498),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_547),
.Y(n_776)
);

BUFx8_ASAP7_75t_SL g777 ( 
.A(n_425),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_473),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_559),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_595),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_598),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_530),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_427),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_656),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_601),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_608),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_610),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_621),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_576),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_461),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_624),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_618),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_582),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_636),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_443),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_638),
.Y(n_796)
);

INVxp33_ASAP7_75t_SL g797 ( 
.A(n_728),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_647),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_657),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_687),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_692),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_465),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_498),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_701),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_705),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_706),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_465),
.B(n_2),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_615),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_707),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_631),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_453),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_710),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_464),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_498),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_529),
.B(n_629),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

INVxp33_ASAP7_75t_L g817 ( 
.A(n_428),
.Y(n_817)
);

INVxp33_ASAP7_75t_L g818 ( 
.A(n_428),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_438),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_725),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_498),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_734),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_438),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_448),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_720),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_498),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_642),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_730),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_448),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_550),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_411),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_449),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_449),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_469),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_550),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_469),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_699),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_458),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_599),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_398),
.Y(n_840)
);

INVxp33_ASAP7_75t_SL g841 ( 
.A(n_398),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_568),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_550),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_599),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_673),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_668),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_581),
.Y(n_847)
);

CKINVDCx14_ASAP7_75t_R g848 ( 
.A(n_655),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_550),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_668),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_550),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_408),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_529),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_629),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_637),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_540),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_411),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_649),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_408),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_458),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_408),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_605),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_605),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_605),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_673),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_694),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_673),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_694),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_459),
.Y(n_869)
);

INVxp67_ASAP7_75t_SL g870 ( 
.A(n_459),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_535),
.Y(n_871)
);

CKINVDCx16_ASAP7_75t_R g872 ( 
.A(n_694),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_535),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_429),
.B(n_3),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_402),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_404),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_409),
.Y(n_877)
);

INVxp67_ASAP7_75t_SL g878 ( 
.A(n_585),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_585),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_696),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_400),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_410),
.Y(n_882)
);

BUFx10_ASAP7_75t_L g883 ( 
.A(n_626),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_412),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_414),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_417),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_719),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_738),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_400),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_460),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_420),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_462),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_424),
.Y(n_893)
);

XNOR2x1_ASAP7_75t_L g894 ( 
.A(n_401),
.B(n_3),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_686),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_466),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_686),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_432),
.Y(n_898)
);

INVxp33_ASAP7_75t_L g899 ( 
.A(n_440),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_434),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_697),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_437),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_401),
.Y(n_903)
);

INVxp67_ASAP7_75t_SL g904 ( 
.A(n_697),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_446),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_447),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_395),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_551),
.B(n_6),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_395),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_451),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_419),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_470),
.Y(n_912)
);

INVxp33_ASAP7_75t_L g913 ( 
.A(n_440),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_475),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_419),
.Y(n_915)
);

INVxp33_ASAP7_75t_SL g916 ( 
.A(n_426),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_472),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_426),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_476),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_482),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_396),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_632),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_491),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_495),
.Y(n_924)
);

INVxp33_ASAP7_75t_SL g925 ( 
.A(n_430),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_430),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_500),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_501),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_431),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_396),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_399),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_506),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_509),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_518),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_431),
.Y(n_935)
);

INVxp33_ASAP7_75t_L g936 ( 
.A(n_475),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_519),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_524),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_541),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_543),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_546),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_558),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_563),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_572),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_481),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_578),
.Y(n_946)
);

CKINVDCx14_ASAP7_75t_R g947 ( 
.A(n_399),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_626),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_468),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_484),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_584),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_486),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_588),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_490),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_594),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_609),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_613),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_436),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_616),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_630),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_635),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_639),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_481),
.Y(n_963)
);

CKINVDCx14_ASAP7_75t_R g964 ( 
.A(n_403),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_648),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_659),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_667),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_497),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_670),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_499),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_510),
.Y(n_971)
);

CKINVDCx16_ASAP7_75t_R g972 ( 
.A(n_458),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_674),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_682),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_690),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_691),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_512),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_698),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_522),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_523),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_703),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_739),
.Y(n_982)
);

INVxp33_ASAP7_75t_SL g983 ( 
.A(n_436),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_439),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_502),
.B(n_8),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_439),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_525),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_442),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_403),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_442),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_526),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_444),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_405),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_502),
.Y(n_994)
);

BUFx10_ASAP7_75t_L g995 ( 
.A(n_405),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_444),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_445),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_445),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_679),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_679),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_646),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_680),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_680),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_684),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_646),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_458),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_684),
.Y(n_1007)
);

CKINVDCx14_ASAP7_75t_R g1008 ( 
.A(n_416),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_688),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_688),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_542),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_702),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_544),
.B(n_8),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_702),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_708),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_458),
.Y(n_1016)
);

INVxp33_ASAP7_75t_L g1017 ( 
.A(n_474),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_545),
.B(n_9),
.Y(n_1018)
);

INVxp33_ASAP7_75t_SL g1019 ( 
.A(n_708),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_474),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_474),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_709),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_709),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_711),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_778),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_774),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_778),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_782),
.Y(n_1028)
);

INVxp33_ASAP7_75t_SL g1029 ( 
.A(n_754),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_830),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_851),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_756),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1006),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_758),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_759),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_852),
.B(n_948),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_760),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_783),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_852),
.B(n_452),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_763),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_764),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_852),
.B(n_415),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_795),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_766),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_767),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_972),
.B(n_532),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_922),
.B(n_773),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_811),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_1017),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_813),
.Y(n_1050)
);

INVxp33_ASAP7_75t_SL g1051 ( 
.A(n_790),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_880),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_768),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_880),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_769),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_771),
.Y(n_1056)
);

BUFx10_ASAP7_75t_L g1057 ( 
.A(n_790),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_782),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_842),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_772),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_847),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_789),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_855),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_831),
.Y(n_1064)
);

INVxp67_ASAP7_75t_SL g1065 ( 
.A(n_1017),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_776),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_888),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_779),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_858),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_887),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_888),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_780),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_777),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_777),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_781),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_789),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_840),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_793),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_770),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_785),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_797),
.B(n_536),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_793),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_810),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_786),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_808),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_749),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_837),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_797),
.B(n_597),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_907),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1006),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_889),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_889),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_787),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_831),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1020),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_788),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_791),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_907),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_909),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_909),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_794),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_796),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_947),
.B(n_607),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_810),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_798),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_911),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_921),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_799),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1020),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_827),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_947),
.B(n_625),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_980),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_911),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_800),
.Y(n_1114)
);

INVxp67_ASAP7_75t_SL g1115 ( 
.A(n_871),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_991),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_921),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_827),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_801),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_804),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_805),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_806),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_809),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_930),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_848),
.B(n_964),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_930),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_R g1127 ( 
.A(n_848),
.B(n_964),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_812),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_816),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_820),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_931),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_822),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_742),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_918),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_743),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_871),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_918),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_931),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_895),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_744),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_929),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_929),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_895),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_989),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_784),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_989),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_745),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_993),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_935),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_993),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_890),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_935),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_892),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_984),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_746),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_984),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_741),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_896),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_748),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_949),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_750),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_751),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_990),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_950),
.Y(n_1164)
);

INVxp67_ASAP7_75t_SL g1165 ( 
.A(n_901),
.Y(n_1165)
);

INVxp67_ASAP7_75t_SL g1166 ( 
.A(n_901),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_752),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1021),
.B(n_644),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_741),
.Y(n_1169)
);

BUFx10_ASAP7_75t_L g1170 ( 
.A(n_792),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_755),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_990),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_997),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_997),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_952),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_994),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1000),
.Y(n_1177)
);

INVxp33_ASAP7_75t_SL g1178 ( 
.A(n_792),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_954),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_994),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_747),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_747),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_968),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_970),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_761),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1005),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_971),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1008),
.B(n_416),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_1000),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1005),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_1016),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_857),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1004),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_857),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_977),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1008),
.B(n_418),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_979),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_869),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_869),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_859),
.B(n_418),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_987),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_873),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_881),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1001),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1011),
.Y(n_1205)
);

INVxp33_ASAP7_75t_L g1206 ( 
.A(n_903),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_R g1207 ( 
.A(n_828),
.B(n_454),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_828),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_865),
.B(n_455),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1112),
.B(n_872),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1176),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1133),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1135),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1064),
.B(n_1094),
.Y(n_1214)
);

AND2x2_ASAP7_75t_SL g1215 ( 
.A(n_1081),
.B(n_765),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1151),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1180),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1140),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1147),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1116),
.B(n_867),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1186),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1155),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1159),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1191),
.B(n_870),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1033),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1190),
.Y(n_1226)
);

NAND2xp33_ASAP7_75t_SL g1227 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1047),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_1064),
.B(n_861),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1161),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1192),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1025),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_1073),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1115),
.B(n_862),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1162),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1049),
.B(n_1065),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1090),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1090),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1204),
.B(n_878),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1085),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1167),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1153),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_SL g1243 ( 
.A(n_1086),
.B(n_825),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1136),
.B(n_863),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1194),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1171),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1198),
.Y(n_1247)
);

BUFx12f_ASAP7_75t_L g1248 ( 
.A(n_1074),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1158),
.Y(n_1249)
);

BUFx8_ASAP7_75t_L g1250 ( 
.A(n_1092),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1087),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_R g1252 ( 
.A(n_1160),
.B(n_757),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1199),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1202),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1095),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1032),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1038),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1139),
.B(n_864),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1095),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1109),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1034),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1143),
.B(n_866),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1109),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1164),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1035),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1206),
.B(n_817),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1037),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1040),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1157),
.Y(n_1269)
);

NOR2x1_ASAP7_75t_L g1270 ( 
.A(n_1103),
.B(n_868),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1036),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1165),
.B(n_904),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1175),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1179),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1169),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1206),
.B(n_817),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1183),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1184),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1043),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1041),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1048),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1187),
.Y(n_1283)
);

INVxp33_ASAP7_75t_L g1284 ( 
.A(n_1088),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1089),
.A2(n_894),
.B1(n_908),
.B2(n_874),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1044),
.Y(n_1286)
);

INVxp33_ASAP7_75t_SL g1287 ( 
.A(n_1195),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1166),
.B(n_815),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1077),
.B(n_818),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1169),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1197),
.B(n_985),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1045),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1181),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1134),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1039),
.B(n_986),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1053),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1026),
.B(n_899),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_1057),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1055),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1181),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1056),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1060),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1182),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1066),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1030),
.B(n_899),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1025),
.Y(n_1307)
);

NAND2xp33_ASAP7_75t_L g1308 ( 
.A(n_1098),
.B(n_474),
.Y(n_1308)
);

AND2x6_ASAP7_75t_L g1309 ( 
.A(n_1042),
.B(n_474),
.Y(n_1309)
);

BUFx8_ASAP7_75t_L g1310 ( 
.A(n_1106),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1068),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1185),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1185),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1201),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1111),
.B(n_1188),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1031),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1072),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1075),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1080),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1084),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1050),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1046),
.B(n_913),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1027),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1093),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1096),
.B(n_992),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1097),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1101),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1102),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1105),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1108),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1114),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1205),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1119),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1120),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1059),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1121),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1122),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1123),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1128),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1196),
.A2(n_841),
.B1(n_925),
.B2(n_916),
.Y(n_1340)
);

AND3x2_ASAP7_75t_L g1341 ( 
.A(n_1079),
.B(n_1203),
.C(n_1145),
.Y(n_1341)
);

INVxp33_ASAP7_75t_SL g1342 ( 
.A(n_1099),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1129),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1168),
.B(n_913),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1130),
.B(n_936),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1061),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1132),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1200),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1209),
.B(n_996),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1057),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1100),
.B(n_995),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1107),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1117),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1124),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1126),
.B(n_998),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1131),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1063),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1057),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1138),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1144),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1146),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1148),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1170),
.B(n_818),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1069),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1150),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1170),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1208),
.B(n_999),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1051),
.A2(n_841),
.B1(n_925),
.B2(n_916),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1170),
.Y(n_1369)
);

XOR2xp5_ASAP7_75t_L g1370 ( 
.A(n_1052),
.B(n_1004),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1266),
.B(n_1070),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1316),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1212),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1213),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1225),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1218),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1219),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1211),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1222),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1232),
.A2(n_1137),
.B1(n_1141),
.B2(n_1134),
.Y(n_1380)
);

AND3x1_ASAP7_75t_L g1381 ( 
.A(n_1368),
.B(n_753),
.C(n_1013),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1225),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1358),
.B(n_933),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1322),
.B(n_936),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1215),
.A2(n_1178),
.B1(n_983),
.B2(n_1019),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1223),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1216),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1230),
.Y(n_1388)
);

XOR2x2_ASAP7_75t_SL g1389 ( 
.A(n_1285),
.B(n_894),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1277),
.B(n_915),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1235),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1232),
.A2(n_1141),
.B1(n_1142),
.B2(n_1137),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1289),
.B(n_958),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_SL g1394 ( 
.A(n_1274),
.Y(n_1394)
);

AND2x6_ASAP7_75t_L g1395 ( 
.A(n_1358),
.B(n_555),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1255),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1358),
.B(n_995),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1241),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1246),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1242),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1256),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1211),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1228),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1211),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1306),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1210),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1306),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1272),
.B(n_983),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1322),
.B(n_995),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1228),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1215),
.A2(n_1019),
.B1(n_807),
.B2(n_721),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1358),
.B(n_933),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1261),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1350),
.B(n_1002),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1265),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1363),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1267),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1211),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1285),
.B(n_988),
.C(n_1014),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1344),
.B(n_1207),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1288),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1217),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1237),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1268),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1217),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1217),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1281),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1286),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1217),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1272),
.B(n_1348),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1238),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1292),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1296),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1307),
.A2(n_1149),
.B1(n_1152),
.B2(n_1142),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1299),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1260),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1301),
.Y(n_1437)
);

XNOR2xp5_ASAP7_75t_L g1438 ( 
.A(n_1370),
.B(n_1054),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1307),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1302),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1284),
.B(n_1029),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1288),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1284),
.B(n_883),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1304),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1220),
.B(n_819),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1311),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1317),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1318),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1319),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1344),
.B(n_757),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1226),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1331),
.Y(n_1452)
);

BUFx6f_ASAP7_75t_L g1453 ( 
.A(n_1226),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1333),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1239),
.B(n_1236),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1336),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1338),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1240),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1350),
.B(n_1003),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1269),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1328),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1328),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1251),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1329),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1271),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1276),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1329),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1273),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1334),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1226),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1239),
.B(n_914),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1334),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1345),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1226),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1300),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1343),
.Y(n_1476)
);

AND2x6_ASAP7_75t_L g1477 ( 
.A(n_1366),
.B(n_555),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1343),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1236),
.B(n_1224),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1303),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1323),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1224),
.B(n_945),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1324),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1245),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1326),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1330),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1347),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1312),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1340),
.A2(n_721),
.B1(n_723),
.B2(n_711),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1323),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1247),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1253),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1221),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1231),
.Y(n_1494)
);

AND2x6_ASAP7_75t_L g1495 ( 
.A(n_1369),
.B(n_555),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1294),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_SL g1497 ( 
.A(n_1274),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1231),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1254),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1254),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1320),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1345),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1280),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1315),
.A2(n_1018),
.B1(n_722),
.B2(n_876),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1320),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1315),
.B(n_963),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1279),
.B(n_1283),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1354),
.A2(n_856),
.B1(n_802),
.B2(n_1007),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1273),
.B(n_1001),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1291),
.A2(n_877),
.B1(n_882),
.B2(n_875),
.Y(n_1510)
);

AND2x6_ASAP7_75t_L g1511 ( 
.A(n_1422),
.B(n_1354),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1375),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1408),
.B(n_1287),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1408),
.B(n_1287),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1410),
.B(n_1091),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1389),
.A2(n_1327),
.B1(n_1337),
.B2(n_1320),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1468),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1503),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1473),
.B(n_1297),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1356),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1468),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1420),
.A2(n_1264),
.B1(n_1278),
.B2(n_1249),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1373),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1502),
.B(n_1356),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1422),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1374),
.Y(n_1526)
);

BUFx10_ASAP7_75t_L g1527 ( 
.A(n_1394),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1376),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1502),
.B(n_1342),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1445),
.B(n_1393),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_R g1531 ( 
.A(n_1387),
.B(n_1314),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1403),
.B(n_1332),
.C(n_1346),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1403),
.A2(n_1291),
.B1(n_1353),
.B2(n_1359),
.C(n_1352),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1422),
.Y(n_1534)
);

AND2x6_ASAP7_75t_L g1535 ( 
.A(n_1422),
.B(n_1214),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1479),
.B(n_1297),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1382),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1377),
.A2(n_1337),
.B1(n_1339),
.B2(n_1327),
.Y(n_1538)
);

NAND2x1_ASAP7_75t_L g1539 ( 
.A(n_1425),
.B(n_1327),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1463),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1425),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1379),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1390),
.B(n_1507),
.Y(n_1543)
);

OAI21xp33_ASAP7_75t_L g1544 ( 
.A1(n_1385),
.A2(n_1342),
.B(n_1357),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1421),
.B(n_1275),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1386),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1388),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1391),
.A2(n_1337),
.B1(n_1339),
.B2(n_1327),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1384),
.B(n_1305),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1387),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1503),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_1463),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1371),
.B(n_1257),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1421),
.B(n_1275),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1455),
.B(n_1305),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1430),
.B(n_1409),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1396),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1398),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1482),
.B(n_1214),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1399),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1405),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1401),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1471),
.B(n_1234),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1430),
.B(n_1362),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1461),
.A2(n_1360),
.B1(n_1365),
.B2(n_1361),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1501),
.A2(n_1308),
.B(n_1295),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1442),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1439),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1506),
.B(n_1234),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1425),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1416),
.B(n_1351),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1413),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1490),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1405),
.Y(n_1574)
);

BUFx10_ASAP7_75t_L g1575 ( 
.A(n_1394),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1415),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1425),
.B(n_1337),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1406),
.B(n_1113),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1400),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1400),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1429),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1417),
.A2(n_1339),
.B1(n_1325),
.B2(n_1245),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1442),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1497),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1416),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1424),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_SL g1587 ( 
.A(n_1497),
.B(n_1364),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1481),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1429),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1429),
.B(n_1339),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1458),
.B(n_1257),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1427),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1407),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1407),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1383),
.B(n_1325),
.Y(n_1595)
);

INVxp33_ASAP7_75t_L g1596 ( 
.A(n_1438),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1429),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1383),
.B(n_1229),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1428),
.A2(n_1245),
.B1(n_1309),
.B2(n_937),
.Y(n_1599)
);

XNOR2xp5_ASAP7_75t_L g1600 ( 
.A(n_1380),
.B(n_1067),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1432),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1509),
.B(n_1244),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1433),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1435),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1381),
.A2(n_1355),
.B1(n_1270),
.B2(n_1295),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_SL g1606 ( 
.A(n_1414),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1450),
.B(n_1351),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1412),
.Y(n_1608)
);

INVxp33_ASAP7_75t_L g1609 ( 
.A(n_1392),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1412),
.Y(n_1610)
);

OR2x6_ASAP7_75t_L g1611 ( 
.A(n_1434),
.B(n_1282),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1453),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1512),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1536),
.B(n_1555),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1519),
.B(n_1458),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1529),
.B(n_1355),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1513),
.B(n_1149),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1549),
.B(n_1321),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1518),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1609),
.A2(n_1419),
.B1(n_1154),
.B2(n_1156),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1518),
.Y(n_1621)
);

AND2x2_ASAP7_75t_SL g1622 ( 
.A(n_1516),
.B(n_1308),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1609),
.A2(n_1154),
.B1(n_1156),
.B2(n_1152),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1595),
.B(n_1437),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1512),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1529),
.B(n_1321),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1537),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1551),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1513),
.B(n_1335),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1537),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1557),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1514),
.B(n_1335),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1557),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1514),
.B(n_1163),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1595),
.A2(n_1172),
.B1(n_1174),
.B2(n_1163),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1545),
.B(n_1367),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1561),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_SL g1638 ( 
.A(n_1550),
.B(n_1233),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1545),
.B(n_1367),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1561),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1172),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1530),
.B(n_1440),
.Y(n_1642)
);

INVx4_ASAP7_75t_L g1643 ( 
.A(n_1535),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1554),
.B(n_1414),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1174),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1574),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1574),
.Y(n_1647)
);

AND2x2_ASAP7_75t_SL g1648 ( 
.A(n_1516),
.B(n_1453),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1520),
.B(n_1459),
.Y(n_1649)
);

OAI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1544),
.A2(n_1173),
.B1(n_1489),
.B2(n_1411),
.C(n_1441),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1520),
.B(n_1459),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1554),
.B(n_1591),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1593),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1552),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1593),
.Y(n_1655)
);

OR2x6_ASAP7_75t_L g1656 ( 
.A(n_1598),
.B(n_1453),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1551),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1522),
.B(n_1441),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_L g1659 ( 
.A(n_1541),
.B(n_1378),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1535),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1563),
.B(n_1444),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1556),
.B(n_1446),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1553),
.B(n_1243),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1540),
.B(n_1177),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1532),
.B(n_1227),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1525),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1556),
.A2(n_1397),
.B(n_1443),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1594),
.Y(n_1668)
);

NOR2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1580),
.B(n_1298),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1594),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1543),
.B(n_1447),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1525),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1515),
.B(n_1177),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1559),
.B(n_1448),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1525),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1569),
.B(n_1602),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1642),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1614),
.B(n_1567),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1621),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1629),
.B(n_1567),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1643),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1642),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1654),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1641),
.A2(n_1600),
.B1(n_1372),
.B2(n_1193),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_R g1686 ( 
.A(n_1638),
.B(n_1531),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1618),
.B(n_1583),
.Y(n_1687)
);

OR2x6_ASAP7_75t_SL g1688 ( 
.A(n_1615),
.B(n_1294),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1645),
.B(n_1649),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1583),
.Y(n_1690)
);

AO221x1_ASAP7_75t_L g1691 ( 
.A1(n_1672),
.A2(n_1565),
.B1(n_1534),
.B2(n_1525),
.C(n_1453),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1621),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1662),
.A2(n_1397),
.B(n_1577),
.Y(n_1693)
);

AND2x6_ASAP7_75t_SL g1694 ( 
.A(n_1673),
.B(n_1611),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1617),
.B(n_1596),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1634),
.B(n_1596),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1643),
.B(n_1581),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1671),
.B(n_1585),
.Y(n_1698)
);

NOR2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1580),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1664),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1661),
.B(n_1585),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1622),
.B(n_1564),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1676),
.B(n_1579),
.Y(n_1703)
);

A2O1A1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1667),
.A2(n_1564),
.B(n_1571),
.C(n_1605),
.Y(n_1704)
);

NOR2x1p5_ASAP7_75t_L g1705 ( 
.A(n_1657),
.B(n_1248),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1625),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1624),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1669),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1674),
.A2(n_1590),
.B(n_1577),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1613),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1622),
.B(n_1571),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1625),
.Y(n_1712)
);

NOR2xp67_ASAP7_75t_L g1713 ( 
.A(n_1619),
.B(n_1584),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1624),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1613),
.Y(n_1715)
);

BUFx4f_ASAP7_75t_L g1716 ( 
.A(n_1624),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1620),
.A2(n_1193),
.B1(n_1189),
.B2(n_1611),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1632),
.B(n_1598),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1627),
.Y(n_1719)
);

OR2x6_ASAP7_75t_L g1720 ( 
.A(n_1644),
.B(n_1611),
.Y(n_1720)
);

NAND2xp33_ASAP7_75t_SL g1721 ( 
.A(n_1686),
.B(n_1531),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1689),
.B(n_1648),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1686),
.B(n_1648),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1680),
.B(n_1672),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_SL g1725 ( 
.A(n_1699),
.B(n_1669),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1678),
.B(n_1658),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_SL g1728 ( 
.A(n_1703),
.B(n_1252),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1701),
.B(n_1672),
.Y(n_1729)
);

NAND2xp33_ASAP7_75t_SL g1730 ( 
.A(n_1681),
.B(n_1665),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1681),
.B(n_1660),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1677),
.B(n_1663),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1698),
.B(n_1652),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1690),
.B(n_1716),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1716),
.B(n_1672),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1695),
.B(n_1675),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1683),
.B(n_1626),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1684),
.B(n_1616),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1695),
.B(n_1696),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1700),
.B(n_1517),
.Y(n_1740)
);

NAND2xp33_ASAP7_75t_SL g1741 ( 
.A(n_1681),
.B(n_1660),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_R g1742 ( 
.A(n_1720),
.B(n_1252),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1714),
.B(n_1521),
.Y(n_1743)
);

AND2x4_ASAP7_75t_SL g1744 ( 
.A(n_1681),
.B(n_1656),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1696),
.B(n_1675),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1718),
.B(n_1524),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1704),
.B(n_1675),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1704),
.B(n_1675),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1688),
.B(n_1189),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1679),
.B(n_1675),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1679),
.B(n_1587),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1692),
.B(n_1619),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1692),
.B(n_1711),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1707),
.B(n_1524),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1711),
.B(n_1628),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1707),
.B(n_1523),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_SL g1757 ( 
.A(n_1717),
.B(n_1071),
.Y(n_1757)
);

NAND2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1708),
.B(n_1606),
.Y(n_1758)
);

NAND2xp33_ASAP7_75t_SL g1759 ( 
.A(n_1705),
.B(n_1606),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1682),
.B(n_1584),
.Y(n_1760)
);

NAND2xp33_ASAP7_75t_SL g1761 ( 
.A(n_1682),
.B(n_1636),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_SL g1762 ( 
.A(n_1697),
.B(n_1639),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1697),
.B(n_1628),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1697),
.B(n_1666),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1732),
.B(n_1702),
.Y(n_1765)
);

NAND2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1747),
.B(n_1702),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1744),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1730),
.A2(n_1691),
.B(n_1693),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1721),
.A2(n_1742),
.B1(n_1728),
.B2(n_1762),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1759),
.Y(n_1770)
);

BUFx2_ASAP7_75t_SL g1771 ( 
.A(n_1751),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1729),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1730),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1748),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1744),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1724),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1731),
.A2(n_1709),
.B(n_1590),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1737),
.B(n_1710),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1727),
.B(n_1715),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1731),
.A2(n_1548),
.B(n_1538),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1741),
.A2(n_1548),
.B(n_1538),
.Y(n_1782)
);

O2A1O1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1739),
.A2(n_1650),
.B(n_1533),
.C(n_1443),
.Y(n_1783)
);

BUFx8_ASAP7_75t_L g1784 ( 
.A(n_1721),
.Y(n_1784)
);

AND2x2_ASAP7_75t_SL g1785 ( 
.A(n_1757),
.B(n_1685),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1754),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1764),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1749),
.B(n_1496),
.Y(n_1788)
);

CKINVDCx16_ASAP7_75t_R g1789 ( 
.A(n_1725),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1756),
.Y(n_1790)
);

CKINVDCx8_ASAP7_75t_R g1791 ( 
.A(n_1758),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1750),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1741),
.A2(n_1761),
.B(n_1755),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1736),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1746),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1745),
.B(n_1753),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1743),
.Y(n_1797)
);

AOI222xp33_ASAP7_75t_L g1798 ( 
.A1(n_1722),
.A2(n_1685),
.B1(n_1635),
.B2(n_1623),
.C1(n_845),
.C2(n_731),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1760),
.B(n_1713),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1752),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1733),
.B(n_1719),
.Y(n_1801)
);

INVx5_ASAP7_75t_L g1802 ( 
.A(n_1723),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1734),
.A2(n_1504),
.B(n_1510),
.C(n_1227),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1735),
.A2(n_1539),
.B(n_1666),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1763),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1740),
.Y(n_1807)
);

INVx4_ASAP7_75t_L g1808 ( 
.A(n_1744),
.Y(n_1808)
);

CKINVDCx11_ASAP7_75t_R g1809 ( 
.A(n_1721),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1732),
.B(n_1712),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1747),
.Y(n_1811)
);

BUFx12f_ASAP7_75t_L g1812 ( 
.A(n_1732),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1797),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1765),
.B(n_1720),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1790),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1768),
.A2(n_1712),
.B(n_1706),
.Y(n_1816)
);

AO31x2_ASAP7_75t_L g1817 ( 
.A1(n_1774),
.A2(n_1706),
.A3(n_1630),
.B(n_1631),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1797),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1783),
.A2(n_1803),
.B(n_1785),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1793),
.A2(n_1720),
.B(n_1666),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1790),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1807),
.Y(n_1822)
);

O2A1O1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1798),
.A2(n_1508),
.B(n_1588),
.C(n_926),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1789),
.A2(n_1582),
.B1(n_1028),
.B2(n_1058),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1799),
.A2(n_1568),
.B(n_1573),
.C(n_1349),
.Y(n_1825)
);

OAI21x1_ASAP7_75t_L g1826 ( 
.A1(n_1777),
.A2(n_1630),
.B(n_1627),
.Y(n_1826)
);

O2A1O1Ixp33_ASAP7_75t_SL g1827 ( 
.A1(n_1788),
.A2(n_1009),
.B(n_1012),
.C(n_1010),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_SL g1828 ( 
.A1(n_1769),
.A2(n_1015),
.B(n_1023),
.C(n_1022),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1805),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1776),
.B(n_1778),
.C(n_1794),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1812),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1781),
.A2(n_1640),
.B(n_1631),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1765),
.B(n_1527),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1771),
.B(n_1694),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1807),
.B(n_937),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1770),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1773),
.A2(n_1582),
.B(n_1659),
.Y(n_1837)
);

BUFx12f_ASAP7_75t_L g1838 ( 
.A(n_1770),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1791),
.B(n_1773),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1786),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1785),
.A2(n_845),
.B(n_967),
.C(n_962),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1812),
.A2(n_1028),
.B1(n_1058),
.B2(n_1027),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1786),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1782),
.A2(n_1655),
.B(n_1640),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1766),
.A2(n_1511),
.B(n_1309),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1766),
.A2(n_1670),
.B(n_1655),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1795),
.B(n_962),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1804),
.A2(n_1659),
.B(n_1656),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1779),
.B(n_967),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1800),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_L g1851 ( 
.A1(n_1766),
.A2(n_1670),
.B(n_1637),
.Y(n_1851)
);

OAI22x1_ASAP7_75t_L g1852 ( 
.A1(n_1802),
.A2(n_1062),
.B1(n_1104),
.B2(n_1083),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1774),
.A2(n_1656),
.B(n_1534),
.Y(n_1853)
);

O2A1O1Ixp33_ASAP7_75t_SL g1854 ( 
.A1(n_1792),
.A2(n_1791),
.B(n_1780),
.C(n_1771),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1811),
.A2(n_1534),
.B(n_1566),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1779),
.B(n_969),
.Y(n_1856)
);

O2A1O1Ixp33_ASAP7_75t_SL g1857 ( 
.A1(n_1792),
.A2(n_1806),
.B(n_1024),
.C(n_1772),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_SL g1858 ( 
.A1(n_1806),
.A2(n_1612),
.B(n_1589),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1795),
.B(n_1578),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1796),
.A2(n_1083),
.B1(n_1104),
.B2(n_1062),
.Y(n_1860)
);

A2O1A1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1802),
.A2(n_969),
.B(n_976),
.C(n_729),
.Y(n_1861)
);

OAI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1772),
.A2(n_1637),
.B(n_1633),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1805),
.B(n_976),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1802),
.A2(n_1566),
.B(n_1581),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1801),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1767),
.A2(n_1646),
.B(n_1633),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1810),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1802),
.A2(n_1597),
.B(n_1589),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1801),
.B(n_884),
.Y(n_1869)
);

OAI21x1_ASAP7_75t_SL g1870 ( 
.A1(n_1800),
.A2(n_1528),
.B(n_1526),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1810),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1800),
.B(n_1250),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1802),
.A2(n_729),
.B(n_726),
.C(n_727),
.Y(n_1873)
);

AOI221x1_ASAP7_75t_L g1874 ( 
.A1(n_1787),
.A2(n_829),
.B1(n_832),
.B2(n_824),
.C(n_823),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1796),
.A2(n_1612),
.B(n_1597),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1809),
.A2(n_1118),
.B1(n_1110),
.B2(n_1078),
.Y(n_1876)
);

OAI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1775),
.A2(n_1511),
.B(n_1309),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1787),
.B(n_1527),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1787),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1809),
.B(n_1250),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1865),
.Y(n_1881)
);

OR2x6_ASAP7_75t_L g1882 ( 
.A(n_1858),
.B(n_1775),
.Y(n_1882)
);

OAI21x1_ASAP7_75t_L g1883 ( 
.A1(n_1816),
.A2(n_1767),
.B(n_1647),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1870),
.A2(n_1767),
.B(n_1647),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1850),
.Y(n_1885)
);

OAI21x1_ASAP7_75t_L g1886 ( 
.A1(n_1819),
.A2(n_1653),
.B(n_1646),
.Y(n_1886)
);

CKINVDCx16_ASAP7_75t_R g1887 ( 
.A(n_1839),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1819),
.A2(n_1787),
.B1(n_1118),
.B2(n_1110),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1871),
.B(n_1787),
.Y(n_1889)
);

AO31x2_ASAP7_75t_L g1890 ( 
.A1(n_1853),
.A2(n_1808),
.A3(n_1775),
.B(n_762),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1831),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1824),
.A2(n_1076),
.B1(n_1082),
.B2(n_1608),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1867),
.Y(n_1893)
);

BUFx2_ASAP7_75t_SL g1894 ( 
.A(n_1836),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1815),
.B(n_1808),
.Y(n_1895)
);

INVx8_ASAP7_75t_L g1896 ( 
.A(n_1838),
.Y(n_1896)
);

A2O1A1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1841),
.A2(n_726),
.B(n_727),
.C(n_723),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_SL g1898 ( 
.A1(n_1836),
.A2(n_1808),
.B(n_1784),
.Y(n_1898)
);

OR2x6_ASAP7_75t_L g1899 ( 
.A(n_1820),
.B(n_1784),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1830),
.A2(n_1835),
.B(n_1847),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_SL g1901 ( 
.A1(n_1839),
.A2(n_1784),
.B(n_854),
.Y(n_1901)
);

INVx4_ASAP7_75t_L g1902 ( 
.A(n_1878),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_R g1903 ( 
.A(n_1880),
.B(n_1575),
.Y(n_1903)
);

OAI21x1_ASAP7_75t_L g1904 ( 
.A1(n_1855),
.A2(n_1668),
.B(n_1546),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1843),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1813),
.Y(n_1906)
);

OAI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1832),
.A2(n_1547),
.B(n_1542),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1879),
.Y(n_1908)
);

A2O1A1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1823),
.A2(n_1834),
.B(n_1825),
.C(n_1872),
.Y(n_1909)
);

AO21x2_ASAP7_75t_L g1910 ( 
.A1(n_1835),
.A2(n_834),
.B(n_833),
.Y(n_1910)
);

O2A1O1Ixp33_ASAP7_75t_L g1911 ( 
.A1(n_1828),
.A2(n_1827),
.B(n_1873),
.C(n_1861),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1824),
.A2(n_733),
.B1(n_736),
.B2(n_732),
.C(n_731),
.Y(n_1912)
);

AO21x2_ASAP7_75t_L g1913 ( 
.A1(n_1847),
.A2(n_839),
.B(n_836),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1840),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1821),
.B(n_1829),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1849),
.B(n_761),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1818),
.Y(n_1917)
);

OAI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1844),
.A2(n_1560),
.B(n_1558),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_L g1919 ( 
.A1(n_1864),
.A2(n_1572),
.B(n_1562),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1822),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1854),
.A2(n_1570),
.B(n_1541),
.Y(n_1921)
);

OAI21x1_ASAP7_75t_L g1922 ( 
.A1(n_1866),
.A2(n_1826),
.B(n_1846),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1869),
.B(n_762),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1817),
.Y(n_1924)
);

BUFx8_ASAP7_75t_SL g1925 ( 
.A(n_1833),
.Y(n_1925)
);

O2A1O1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1857),
.A2(n_886),
.B(n_891),
.C(n_885),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1852),
.A2(n_736),
.B1(n_737),
.B2(n_733),
.C(n_732),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1863),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1887),
.A2(n_1876),
.B1(n_1842),
.B2(n_1856),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1888),
.A2(n_1860),
.B1(n_1814),
.B2(n_1859),
.Y(n_1930)
);

AOI221xp5_ASAP7_75t_L g1931 ( 
.A1(n_1888),
.A2(n_737),
.B1(n_554),
.B2(n_557),
.C(n_552),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1896),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1902),
.B(n_1817),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1896),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1912),
.A2(n_1310),
.B1(n_1837),
.B2(n_1610),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1905),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1899),
.A2(n_1848),
.B(n_1868),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_SL g1938 ( 
.A1(n_1900),
.A2(n_1899),
.B1(n_1901),
.B2(n_1310),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1902),
.B(n_1817),
.Y(n_1939)
);

OR2x6_ASAP7_75t_L g1940 ( 
.A(n_1899),
.B(n_1882),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1909),
.A2(n_1875),
.B1(n_1845),
.B2(n_1511),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1906),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1894),
.A2(n_1877),
.B1(n_1511),
.B2(n_560),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1917),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1915),
.B(n_1908),
.Y(n_1945)
);

INVx4_ASAP7_75t_SL g1946 ( 
.A(n_1890),
.Y(n_1946)
);

NAND2x1p5_ASAP7_75t_L g1947 ( 
.A(n_1928),
.B(n_1851),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1915),
.B(n_1862),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1882),
.A2(n_1877),
.B1(n_565),
.B2(n_567),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1896),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_1925),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1924),
.Y(n_1952)
);

CKINVDCx9p33_ASAP7_75t_R g1953 ( 
.A(n_1898),
.Y(n_1953)
);

OAI21x1_ASAP7_75t_L g1954 ( 
.A1(n_1922),
.A2(n_1874),
.B(n_853),
.Y(n_1954)
);

AO21x2_ASAP7_75t_L g1955 ( 
.A1(n_1923),
.A2(n_846),
.B(n_844),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1912),
.A2(n_1586),
.B1(n_1592),
.B2(n_1576),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1920),
.Y(n_1957)
);

AOI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1927),
.A2(n_574),
.B1(n_577),
.B2(n_571),
.C(n_549),
.Y(n_1958)
);

INVx4_ASAP7_75t_L g1959 ( 
.A(n_1932),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1951),
.B(n_1891),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1936),
.Y(n_1961)
);

AOI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1929),
.A2(n_1923),
.B(n_1900),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1940),
.B(n_1885),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1935),
.A2(n_1892),
.B1(n_1913),
.B2(n_1910),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1942),
.Y(n_1965)
);

NAND3xp33_ASAP7_75t_L g1966 ( 
.A(n_1931),
.B(n_1927),
.C(n_1911),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1944),
.Y(n_1967)
);

OAI221xp5_ASAP7_75t_L g1968 ( 
.A1(n_1935),
.A2(n_1897),
.B1(n_1892),
.B2(n_1911),
.C(n_1889),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1951),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1952),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1948),
.A2(n_1885),
.B(n_1919),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1957),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1945),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1933),
.B(n_1881),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1939),
.B(n_1908),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1937),
.A2(n_1884),
.B(n_1895),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1947),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1955),
.A2(n_1913),
.B1(n_1910),
.B2(n_1928),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1947),
.B(n_1893),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1952),
.Y(n_1980)
);

AND2x4_ASAP7_75t_SL g1981 ( 
.A(n_1940),
.B(n_1882),
.Y(n_1981)
);

AOI222xp33_ASAP7_75t_L g1982 ( 
.A1(n_1930),
.A2(n_883),
.B1(n_850),
.B2(n_583),
.C1(n_590),
.C2(n_619),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1940),
.B(n_1916),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1955),
.A2(n_1914),
.B1(n_1904),
.B2(n_1886),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1961),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_R g1986 ( 
.A(n_1960),
.B(n_1903),
.Y(n_1986)
);

XNOR2xp5_ASAP7_75t_L g1987 ( 
.A(n_1969),
.B(n_1981),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1981),
.B(n_1932),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1971),
.Y(n_1989)
);

NAND2xp33_ASAP7_75t_R g1990 ( 
.A(n_1963),
.B(n_1903),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1973),
.B(n_1930),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1961),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1969),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1971),
.Y(n_1994)
);

OR2x6_ASAP7_75t_L g1995 ( 
.A(n_1959),
.B(n_1950),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1963),
.B(n_1950),
.Y(n_1996)
);

NAND2xp33_ASAP7_75t_SL g1997 ( 
.A(n_1959),
.B(n_1934),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1965),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1963),
.B(n_1938),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1965),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1967),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1983),
.Y(n_2002)
);

XNOR2xp5_ASAP7_75t_L g2003 ( 
.A(n_1966),
.B(n_1943),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1959),
.B(n_1946),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_R g2005 ( 
.A(n_1963),
.B(n_1341),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_R g2006 ( 
.A(n_1962),
.B(n_1341),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_R g2007 ( 
.A(n_1962),
.B(n_1575),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1967),
.B(n_1949),
.Y(n_2008)
);

NAND2xp33_ASAP7_75t_R g2009 ( 
.A(n_1976),
.B(n_1953),
.Y(n_2009)
);

OR2x6_ASAP7_75t_L g2010 ( 
.A(n_1966),
.B(n_1975),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1968),
.B(n_1958),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1972),
.Y(n_2012)
);

OR2x6_ASAP7_75t_L g2013 ( 
.A(n_1975),
.B(n_1926),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1974),
.B(n_1977),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1972),
.B(n_1941),
.Y(n_2015)
);

NAND2xp33_ASAP7_75t_SL g2016 ( 
.A(n_1977),
.B(n_1953),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_1979),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_2010),
.B(n_1970),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1996),
.B(n_1946),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1985),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1985),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2001),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1988),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1995),
.B(n_1970),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2001),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1995),
.B(n_1980),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1992),
.Y(n_2027)
);

OR2x2_ASAP7_75t_SL g2028 ( 
.A(n_2008),
.B(n_1980),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_1993),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_2013),
.A2(n_1987),
.B1(n_1991),
.B2(n_1988),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2013),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2003),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_2004),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2004),
.B(n_1946),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_2002),
.B(n_1978),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_2011),
.A2(n_1964),
.B1(n_1982),
.B2(n_1984),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2014),
.B(n_1890),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_2000),
.B(n_1954),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2029),
.B(n_2012),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_2036),
.A2(n_2006),
.B1(n_2007),
.B2(n_1999),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2031),
.B(n_2015),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2031),
.B(n_1998),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2023),
.B(n_1989),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2023),
.B(n_1994),
.Y(n_2044)
);

OAI21xp33_ASAP7_75t_L g2045 ( 
.A1(n_2017),
.A2(n_2009),
.B(n_1956),
.Y(n_2045)
);

NAND3xp33_ASAP7_75t_L g2046 ( 
.A(n_2018),
.B(n_2016),
.C(n_1997),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2023),
.B(n_1986),
.Y(n_2047)
);

OR2x6_ASAP7_75t_SL g2048 ( 
.A(n_2030),
.B(n_2032),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_2018),
.B(n_2035),
.C(n_2026),
.Y(n_2049)
);

OAI21xp33_ASAP7_75t_L g2050 ( 
.A1(n_2017),
.A2(n_1956),
.B(n_614),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2035),
.B(n_1926),
.Y(n_2051)
);

NAND4xp25_ASAP7_75t_L g2052 ( 
.A(n_2017),
.B(n_1990),
.C(n_2005),
.D(n_1921),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_2017),
.B(n_1921),
.Y(n_2053)
);

OA21x2_ASAP7_75t_L g2054 ( 
.A1(n_2032),
.A2(n_1883),
.B(n_1907),
.Y(n_2054)
);

NOR2x1_ASAP7_75t_L g2055 ( 
.A(n_2047),
.B(n_2027),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2042),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2043),
.B(n_2033),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2039),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2044),
.B(n_2033),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2048),
.A2(n_2028),
.B1(n_2035),
.B2(n_2027),
.Y(n_2060)
);

AOI31xp33_ASAP7_75t_SL g2061 ( 
.A1(n_2040),
.A2(n_2041),
.A3(n_2051),
.B(n_2046),
.Y(n_2061)
);

OAI211xp5_ASAP7_75t_L g2062 ( 
.A1(n_2045),
.A2(n_2021),
.B(n_2022),
.C(n_2020),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2054),
.Y(n_2063)
);

NAND2x1_ASAP7_75t_L g2064 ( 
.A(n_2057),
.B(n_2024),
.Y(n_2064)
);

NOR2x1_ASAP7_75t_L g2065 ( 
.A(n_2061),
.B(n_2049),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2055),
.B(n_2050),
.Y(n_2066)
);

NAND4xp25_ASAP7_75t_L g2067 ( 
.A(n_2058),
.B(n_2050),
.C(n_2052),
.D(n_2021),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_2056),
.B(n_2060),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_2059),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_2060),
.A2(n_2054),
.B1(n_2053),
.B2(n_2037),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2069),
.B(n_2024),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2068),
.Y(n_2072)
);

INVxp67_ASAP7_75t_SL g2073 ( 
.A(n_2065),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_2066),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2064),
.Y(n_2075)
);

OAI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2073),
.A2(n_2070),
.B1(n_2072),
.B2(n_2062),
.C(n_2074),
.Y(n_2076)
);

OAI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_2074),
.A2(n_2067),
.B1(n_2063),
.B2(n_2028),
.Y(n_2077)
);

CKINVDCx16_ASAP7_75t_R g2078 ( 
.A(n_2071),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2078),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2076),
.B(n_2071),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2079),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_2080),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_2079),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2083),
.B(n_2075),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_2082),
.B(n_2062),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_2084),
.A2(n_2077),
.B(n_2081),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2085),
.B(n_2026),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2084),
.B(n_2020),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_2086),
.A2(n_2025),
.B(n_2022),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2087),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2088),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2087),
.A2(n_2034),
.B1(n_2025),
.B2(n_2019),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2091),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2090),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2089),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2092),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2094),
.A2(n_2096),
.B1(n_2095),
.B2(n_2093),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2093),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2093),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2094),
.A2(n_1349),
.B(n_2034),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2093),
.Y(n_2101)
);

OAI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_2094),
.A2(n_2019),
.B(n_2037),
.Y(n_2102)
);

OAI211xp5_ASAP7_75t_SL g2103 ( 
.A1(n_2096),
.A2(n_898),
.B(n_900),
.C(n_893),
.Y(n_2103)
);

BUFx2_ASAP7_75t_L g2104 ( 
.A(n_2093),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2094),
.A2(n_2019),
.B(n_2038),
.Y(n_2105)
);

NOR2x1_ASAP7_75t_SL g2106 ( 
.A(n_2094),
.B(n_2038),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2093),
.Y(n_2107)
);

XOR2xp5_ASAP7_75t_L g2108 ( 
.A(n_2096),
.B(n_819),
.Y(n_2108)
);

OAI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_2096),
.A2(n_627),
.B1(n_628),
.B2(n_622),
.C(n_579),
.Y(n_2109)
);

AOI221xp5_ASAP7_75t_L g2110 ( 
.A1(n_2094),
.A2(n_640),
.B1(n_650),
.B2(n_634),
.C(n_633),
.Y(n_2110)
);

OAI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_2104),
.A2(n_661),
.B(n_666),
.C(n_660),
.Y(n_2111)
);

OAI211xp5_ASAP7_75t_L g2112 ( 
.A1(n_2098),
.A2(n_675),
.B(n_677),
.C(n_671),
.Y(n_2112)
);

INVxp67_ASAP7_75t_L g2113 ( 
.A(n_2108),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2097),
.A2(n_740),
.B(n_902),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_2099),
.A2(n_1452),
.B1(n_1454),
.B2(n_1449),
.Y(n_2115)
);

O2A1O1Ixp5_ASAP7_75t_L g2116 ( 
.A1(n_2101),
.A2(n_1229),
.B(n_1457),
.C(n_1456),
.Y(n_2116)
);

OAI32xp33_ASAP7_75t_L g2117 ( 
.A1(n_2107),
.A2(n_1601),
.A3(n_1604),
.B1(n_1603),
.B2(n_1492),
.Y(n_2117)
);

NOR4xp25_ASAP7_75t_L g2118 ( 
.A(n_2109),
.B(n_906),
.C(n_910),
.D(n_905),
.Y(n_2118)
);

OAI32xp33_ASAP7_75t_L g2119 ( 
.A1(n_2105),
.A2(n_1491),
.A3(n_919),
.B1(n_920),
.B2(n_917),
.Y(n_2119)
);

OAI211xp5_ASAP7_75t_L g2120 ( 
.A1(n_2110),
.A2(n_923),
.B(n_924),
.C(n_912),
.Y(n_2120)
);

NOR3xp33_ASAP7_75t_L g2121 ( 
.A(n_2103),
.B(n_1258),
.C(n_1244),
.Y(n_2121)
);

OAI211xp5_ASAP7_75t_SL g2122 ( 
.A1(n_2100),
.A2(n_928),
.B(n_932),
.C(n_927),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_2102),
.Y(n_2123)
);

OAI211xp5_ASAP7_75t_SL g2124 ( 
.A1(n_2106),
.A2(n_938),
.B(n_939),
.C(n_934),
.Y(n_2124)
);

INVxp67_ASAP7_75t_SL g2125 ( 
.A(n_2104),
.Y(n_2125)
);

AOI211xp5_ASAP7_75t_SL g2126 ( 
.A1(n_2097),
.A2(n_1262),
.B(n_1258),
.C(n_941),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2104),
.B(n_940),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_2097),
.A2(n_943),
.B(n_942),
.Y(n_2128)
);

NOR3xp33_ASAP7_75t_L g2129 ( 
.A(n_2104),
.B(n_1262),
.C(n_946),
.Y(n_2129)
);

AOI21xp5_ASAP7_75t_L g2130 ( 
.A1(n_2097),
.A2(n_951),
.B(n_944),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2104),
.Y(n_2131)
);

AOI321xp33_ASAP7_75t_L g2132 ( 
.A1(n_2097),
.A2(n_953),
.A3(n_956),
.B1(n_959),
.B2(n_957),
.C(n_955),
.Y(n_2132)
);

AOI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2097),
.A2(n_965),
.B1(n_966),
.B2(n_961),
.C(n_960),
.Y(n_2133)
);

AOI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_2097),
.A2(n_975),
.B1(n_978),
.B2(n_974),
.C(n_973),
.Y(n_2134)
);

INVxp67_ASAP7_75t_L g2135 ( 
.A(n_2104),
.Y(n_2135)
);

OAI211xp5_ASAP7_75t_L g2136 ( 
.A1(n_2104),
.A2(n_982),
.B(n_981),
.C(n_422),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2104),
.B(n_883),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2104),
.A2(n_1485),
.B1(n_1486),
.B2(n_1483),
.Y(n_2138)
);

AOI22x1_ASAP7_75t_L g2139 ( 
.A1(n_2104),
.A2(n_1464),
.B1(n_1467),
.B2(n_1462),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2104),
.B(n_873),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2097),
.A2(n_897),
.B1(n_879),
.B2(n_1487),
.C(n_423),
.Y(n_2141)
);

AOI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_2097),
.A2(n_897),
.B1(n_879),
.B2(n_423),
.C(n_433),
.Y(n_2142)
);

AOI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_2097),
.A2(n_433),
.B1(n_435),
.B2(n_422),
.C(n_421),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_2097),
.A2(n_435),
.B(n_421),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2097),
.A2(n_681),
.B(n_678),
.Y(n_2145)
);

NOR3xp33_ASAP7_75t_L g2146 ( 
.A(n_2104),
.B(n_803),
.C(n_775),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2104),
.B(n_9),
.Y(n_2147)
);

AOI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_2097),
.A2(n_681),
.B(n_678),
.Y(n_2148)
);

OAI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_2104),
.A2(n_1472),
.B1(n_1476),
.B2(n_1469),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2104),
.Y(n_2150)
);

OAI211xp5_ASAP7_75t_L g2151 ( 
.A1(n_2104),
.A2(n_685),
.B(n_693),
.C(n_683),
.Y(n_2151)
);

AOI21x1_ASAP7_75t_L g2152 ( 
.A1(n_2104),
.A2(n_803),
.B(n_775),
.Y(n_2152)
);

NAND4xp25_ASAP7_75t_SL g2153 ( 
.A(n_2098),
.B(n_13),
.C(n_10),
.D(n_12),
.Y(n_2153)
);

NOR3xp33_ASAP7_75t_L g2154 ( 
.A(n_2104),
.B(n_821),
.C(n_814),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_SL g2155 ( 
.A1(n_2104),
.A2(n_14),
.B(n_15),
.Y(n_2155)
);

OAI22xp33_ASAP7_75t_SL g2156 ( 
.A1(n_2125),
.A2(n_2150),
.B1(n_2135),
.B2(n_2131),
.Y(n_2156)
);

NAND5xp2_ASAP7_75t_L g2157 ( 
.A(n_2126),
.B(n_19),
.C(n_16),
.D(n_18),
.E(n_20),
.Y(n_2157)
);

OAI311xp33_ASAP7_75t_L g2158 ( 
.A1(n_2137),
.A2(n_1493),
.A3(n_24),
.B1(n_16),
.C1(n_21),
.Y(n_2158)
);

OAI211xp5_ASAP7_75t_SL g2159 ( 
.A1(n_2127),
.A2(n_28),
.B(n_25),
.C(n_26),
.Y(n_2159)
);

OAI21xp33_ASAP7_75t_L g2160 ( 
.A1(n_2155),
.A2(n_685),
.B(n_683),
.Y(n_2160)
);

OA22x2_ASAP7_75t_L g2161 ( 
.A1(n_2123),
.A2(n_695),
.B1(n_704),
.B2(n_693),
.Y(n_2161)
);

XNOR2xp5_ASAP7_75t_L g2162 ( 
.A(n_2147),
.B(n_25),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2123),
.A2(n_1511),
.B1(n_1395),
.B2(n_1478),
.Y(n_2163)
);

OAI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2111),
.A2(n_704),
.B1(n_712),
.B2(n_695),
.Y(n_2164)
);

OAI211xp5_ASAP7_75t_SL g2165 ( 
.A1(n_2140),
.A2(n_2113),
.B(n_2141),
.C(n_2136),
.Y(n_2165)
);

OAI211xp5_ASAP7_75t_SL g2166 ( 
.A1(n_2142),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_2132),
.B(n_712),
.Y(n_2167)
);

A2O1A1Ixp33_ASAP7_75t_L g2168 ( 
.A1(n_2144),
.A2(n_716),
.B(n_717),
.C(n_713),
.Y(n_2168)
);

NOR3xp33_ASAP7_75t_L g2169 ( 
.A(n_2124),
.B(n_821),
.C(n_814),
.Y(n_2169)
);

NAND4xp25_ASAP7_75t_L g2170 ( 
.A(n_2116),
.B(n_34),
.C(n_32),
.D(n_33),
.Y(n_2170)
);

AOI211xp5_ASAP7_75t_L g2171 ( 
.A1(n_2153),
.A2(n_716),
.B(n_717),
.C(n_713),
.Y(n_2171)
);

AOI322xp5_ASAP7_75t_L g2172 ( 
.A1(n_2129),
.A2(n_735),
.A3(n_718),
.B1(n_1599),
.B2(n_835),
.C1(n_826),
.C2(n_849),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2128),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2152),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_2145),
.A2(n_735),
.B(n_718),
.Y(n_2175)
);

NAND3xp33_ASAP7_75t_L g2176 ( 
.A(n_2143),
.B(n_835),
.C(n_826),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2121),
.Y(n_2177)
);

AOI211xp5_ASAP7_75t_L g2178 ( 
.A1(n_2112),
.A2(n_849),
.B(n_843),
.C(n_1494),
.Y(n_2178)
);

AOI221xp5_ASAP7_75t_L g2179 ( 
.A1(n_2118),
.A2(n_843),
.B1(n_477),
.B2(n_478),
.C(n_471),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2114),
.B(n_35),
.Y(n_2180)
);

AOI221xp5_ASAP7_75t_L g2181 ( 
.A1(n_2119),
.A2(n_483),
.B1(n_485),
.B2(n_479),
.C(n_457),
.Y(n_2181)
);

AOI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_2151),
.A2(n_1395),
.B1(n_1535),
.B2(n_1495),
.Y(n_2182)
);

AOI211xp5_ASAP7_75t_L g2183 ( 
.A1(n_2148),
.A2(n_1499),
.B(n_1500),
.C(n_1498),
.Y(n_2183)
);

AOI221xp5_ASAP7_75t_L g2184 ( 
.A1(n_2149),
.A2(n_494),
.B1(n_496),
.B2(n_493),
.C(n_489),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2120),
.Y(n_2185)
);

AOI221xp5_ASAP7_75t_L g2186 ( 
.A1(n_2122),
.A2(n_508),
.B1(n_511),
.B2(n_507),
.C(n_505),
.Y(n_2186)
);

O2A1O1Ixp5_ASAP7_75t_L g2187 ( 
.A1(n_2130),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2115),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2154),
.A2(n_515),
.B1(n_516),
.B2(n_514),
.C(n_513),
.Y(n_2189)
);

AOI211xp5_ASAP7_75t_SL g2190 ( 
.A1(n_2146),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_2190)
);

OAI31xp33_ASAP7_75t_L g2191 ( 
.A1(n_2139),
.A2(n_1599),
.A3(n_44),
.B(n_41),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_2138),
.A2(n_1395),
.B1(n_1535),
.B2(n_1495),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2117),
.A2(n_527),
.B1(n_528),
.B2(n_520),
.C(n_517),
.Y(n_2193)
);

OAI21xp33_ASAP7_75t_L g2194 ( 
.A1(n_2133),
.A2(n_534),
.B(n_533),
.Y(n_2194)
);

AOI211xp5_ASAP7_75t_SL g2195 ( 
.A1(n_2134),
.A2(n_46),
.B(n_43),
.C(n_45),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2135),
.A2(n_539),
.B1(n_548),
.B2(n_537),
.Y(n_2196)
);

AOI221xp5_ASAP7_75t_SL g2197 ( 
.A1(n_2135),
.A2(n_47),
.B1(n_43),
.B2(n_46),
.C(n_48),
.Y(n_2197)
);

AOI211xp5_ASAP7_75t_L g2198 ( 
.A1(n_2150),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2150),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2125),
.A2(n_1395),
.B1(n_1535),
.B2(n_1495),
.Y(n_2200)
);

AOI211xp5_ASAP7_75t_L g2201 ( 
.A1(n_2150),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_2201)
);

AOI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_2125),
.A2(n_556),
.B(n_553),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2125),
.B(n_51),
.Y(n_2203)
);

AOI211xp5_ASAP7_75t_L g2204 ( 
.A1(n_2150),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2125),
.B(n_55),
.Y(n_2205)
);

OAI31xp33_ASAP7_75t_SL g2206 ( 
.A1(n_2150),
.A2(n_57),
.A3(n_55),
.B(n_56),
.Y(n_2206)
);

NOR3xp33_ASAP7_75t_L g2207 ( 
.A(n_2125),
.B(n_562),
.C(n_561),
.Y(n_2207)
);

NOR4xp25_ASAP7_75t_L g2208 ( 
.A(n_2150),
.B(n_60),
.C(n_58),
.D(n_59),
.Y(n_2208)
);

O2A1O1Ixp33_ASAP7_75t_SL g2209 ( 
.A1(n_2150),
.A2(n_62),
.B(n_59),
.C(n_61),
.Y(n_2209)
);

AOI221xp5_ASAP7_75t_L g2210 ( 
.A1(n_2125),
.A2(n_566),
.B1(n_575),
.B2(n_573),
.C(n_569),
.Y(n_2210)
);

OAI211xp5_ASAP7_75t_L g2211 ( 
.A1(n_2125),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_2211)
);

AOI221xp5_ASAP7_75t_L g2212 ( 
.A1(n_2125),
.A2(n_620),
.B1(n_672),
.B2(n_580),
.C(n_586),
.Y(n_2212)
);

NAND4xp25_ASAP7_75t_L g2213 ( 
.A(n_2150),
.B(n_66),
.C(n_63),
.D(n_64),
.Y(n_2213)
);

AOI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2125),
.A2(n_592),
.B(n_589),
.Y(n_2214)
);

AND5x1_ASAP7_75t_L g2215 ( 
.A(n_2141),
.B(n_66),
.C(n_68),
.D(n_70),
.E(n_73),
.Y(n_2215)
);

AOI221xp5_ASAP7_75t_L g2216 ( 
.A1(n_2125),
.A2(n_641),
.B1(n_669),
.B2(n_665),
.C(n_593),
.Y(n_2216)
);

NOR3xp33_ASAP7_75t_L g2217 ( 
.A(n_2125),
.B(n_602),
.C(n_596),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_L g2218 ( 
.A1(n_2135),
.A2(n_604),
.B1(n_606),
.B2(n_603),
.Y(n_2218)
);

AOI211xp5_ASAP7_75t_SL g2219 ( 
.A1(n_2135),
.A2(n_74),
.B(n_68),
.C(n_73),
.Y(n_2219)
);

OAI21xp33_ASAP7_75t_L g2220 ( 
.A1(n_2125),
.A2(n_612),
.B(n_611),
.Y(n_2220)
);

CKINVDCx16_ASAP7_75t_R g2221 ( 
.A(n_2150),
.Y(n_2221)
);

XNOR2xp5_ASAP7_75t_L g2222 ( 
.A(n_2162),
.B(n_74),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2221),
.Y(n_2223)
);

INVxp67_ASAP7_75t_SL g2224 ( 
.A(n_2156),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2199),
.Y(n_2225)
);

NOR2x1_ASAP7_75t_L g2226 ( 
.A(n_2203),
.B(n_76),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_2213),
.A2(n_2160),
.B1(n_2205),
.B2(n_2188),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2206),
.B(n_77),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2161),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_2207),
.A2(n_1395),
.B1(n_1495),
.B2(n_1477),
.Y(n_2230)
);

NOR2x2_ASAP7_75t_L g2231 ( 
.A(n_2215),
.B(n_78),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2187),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2217),
.A2(n_1495),
.B1(n_1477),
.B2(n_1309),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2209),
.Y(n_2234)
);

INVxp67_ASAP7_75t_SL g2235 ( 
.A(n_2167),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2157),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2174),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2211),
.Y(n_2238)
);

AOI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_2159),
.A2(n_1477),
.B1(n_1309),
.B2(n_623),
.Y(n_2239)
);

NOR2xp67_ASAP7_75t_L g2240 ( 
.A(n_2180),
.B(n_78),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2196),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2218),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2198),
.A2(n_643),
.B1(n_645),
.B2(n_617),
.Y(n_2243)
);

OR3x2_ASAP7_75t_L g2244 ( 
.A(n_2170),
.B(n_79),
.C(n_80),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2164),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2165),
.A2(n_1477),
.B1(n_652),
.B2(n_654),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2197),
.A2(n_1477),
.B1(n_658),
.B2(n_662),
.Y(n_2247)
);

NOR2x1_ASAP7_75t_L g2248 ( 
.A(n_2168),
.B(n_80),
.Y(n_2248)
);

NOR2x1_ASAP7_75t_L g2249 ( 
.A(n_2202),
.B(n_82),
.Y(n_2249)
);

NOR3xp33_ASAP7_75t_L g2250 ( 
.A(n_2220),
.B(n_663),
.C(n_651),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2171),
.Y(n_2251)
);

INVxp33_ASAP7_75t_SL g2252 ( 
.A(n_2173),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2185),
.A2(n_676),
.B1(n_664),
.B2(n_1505),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2177),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2214),
.Y(n_2255)
);

NOR2x1_ASAP7_75t_L g2256 ( 
.A(n_2176),
.B(n_82),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2166),
.A2(n_2204),
.B1(n_2201),
.B2(n_2194),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2208),
.Y(n_2258)
);

NOR2x1p5_ASAP7_75t_L g2259 ( 
.A(n_2219),
.B(n_83),
.Y(n_2259)
);

AOI22xp5_ASAP7_75t_L g2260 ( 
.A1(n_2210),
.A2(n_1402),
.B1(n_1404),
.B2(n_1378),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2195),
.B(n_83),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2190),
.B(n_84),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2169),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2212),
.A2(n_1404),
.B1(n_1418),
.B2(n_1402),
.Y(n_2264)
);

AOI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_2216),
.A2(n_2184),
.B1(n_2186),
.B2(n_2183),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2178),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2179),
.A2(n_1426),
.B1(n_1451),
.B2(n_1418),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2181),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2182),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2175),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2193),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2189),
.A2(n_2163),
.B1(n_2158),
.B2(n_2192),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2200),
.Y(n_2273)
);

NAND4xp25_ASAP7_75t_L g2274 ( 
.A(n_2225),
.B(n_2172),
.C(n_2191),
.D(n_95),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_R g2275 ( 
.A(n_2223),
.B(n_2258),
.Y(n_2275)
);

NOR3xp33_ASAP7_75t_SL g2276 ( 
.A(n_2224),
.B(n_86),
.C(n_89),
.Y(n_2276)
);

NOR2x1_ASAP7_75t_L g2277 ( 
.A(n_2234),
.B(n_555),
.Y(n_2277)
);

NAND3xp33_ASAP7_75t_SL g2278 ( 
.A(n_2237),
.B(n_86),
.C(n_89),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2259),
.Y(n_2279)
);

O2A1O1Ixp33_ASAP7_75t_L g2280 ( 
.A1(n_2252),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2232),
.B(n_555),
.Y(n_2281)
);

AOI21xp5_ASAP7_75t_L g2282 ( 
.A1(n_2228),
.A2(n_2262),
.B(n_2222),
.Y(n_2282)
);

NAND3xp33_ASAP7_75t_SL g2283 ( 
.A(n_2254),
.B(n_96),
.C(n_97),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2231),
.Y(n_2284)
);

NAND2x1p5_ASAP7_75t_L g2285 ( 
.A(n_2226),
.B(n_1426),
.Y(n_2285)
);

NAND4xp75_ASAP7_75t_L g2286 ( 
.A(n_2240),
.B(n_98),
.C(n_99),
.D(n_100),
.Y(n_2286)
);

NOR2x1_ASAP7_75t_L g2287 ( 
.A(n_2249),
.B(n_564),
.Y(n_2287)
);

NAND3x1_ASAP7_75t_L g2288 ( 
.A(n_2248),
.B(n_101),
.C(n_102),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_2236),
.B(n_102),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_R g2290 ( 
.A(n_2238),
.B(n_103),
.Y(n_2290)
);

NAND4xp75_ASAP7_75t_L g2291 ( 
.A(n_2240),
.B(n_103),
.C(n_105),
.D(n_106),
.Y(n_2291)
);

INVx1_ASAP7_75t_SL g2292 ( 
.A(n_2261),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2244),
.Y(n_2293)
);

AND3x4_ASAP7_75t_L g2294 ( 
.A(n_2256),
.B(n_105),
.C(n_106),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_L g2295 ( 
.A(n_2229),
.B(n_107),
.Y(n_2295)
);

XOR2x2_ASAP7_75t_L g2296 ( 
.A(n_2227),
.B(n_109),
.Y(n_2296)
);

BUFx2_ASAP7_75t_L g2297 ( 
.A(n_2235),
.Y(n_2297)
);

NAND2x1p5_ASAP7_75t_SL g2298 ( 
.A(n_2241),
.B(n_110),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2255),
.B(n_110),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2270),
.B(n_111),
.Y(n_2300)
);

OAI211xp5_ASAP7_75t_L g2301 ( 
.A1(n_2247),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2242),
.B(n_115),
.Y(n_2302)
);

OR3x2_ASAP7_75t_L g2303 ( 
.A(n_2251),
.B(n_116),
.C(n_117),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2239),
.Y(n_2304)
);

NOR3xp33_ASAP7_75t_L g2305 ( 
.A(n_2268),
.B(n_118),
.C(n_119),
.Y(n_2305)
);

NAND2xp33_ASAP7_75t_L g2306 ( 
.A(n_2250),
.B(n_2243),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_2245),
.B(n_121),
.Y(n_2307)
);

OR4x2_ASAP7_75t_L g2308 ( 
.A(n_2257),
.B(n_123),
.C(n_124),
.D(n_125),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2271),
.B(n_124),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2272),
.B(n_564),
.Y(n_2310)
);

NAND4xp75_ASAP7_75t_L g2311 ( 
.A(n_2263),
.B(n_2266),
.C(n_2253),
.D(n_2273),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2269),
.Y(n_2312)
);

HB1xp67_ASAP7_75t_L g2313 ( 
.A(n_2246),
.Y(n_2313)
);

AOI221xp5_ASAP7_75t_L g2314 ( 
.A1(n_2265),
.A2(n_564),
.B1(n_591),
.B2(n_653),
.C(n_838),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2260),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2264),
.Y(n_2316)
);

AOI31xp33_ASAP7_75t_L g2317 ( 
.A1(n_2267),
.A2(n_126),
.A3(n_127),
.B(n_128),
.Y(n_2317)
);

NOR3x1_ASAP7_75t_L g2318 ( 
.A(n_2230),
.B(n_2233),
.C(n_129),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2223),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_R g2320 ( 
.A(n_2319),
.B(n_129),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_R g2321 ( 
.A(n_2297),
.B(n_130),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_R g2322 ( 
.A(n_2293),
.B(n_130),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_R g2323 ( 
.A(n_2279),
.B(n_131),
.Y(n_2323)
);

XNOR2xp5_ASAP7_75t_L g2324 ( 
.A(n_2284),
.B(n_132),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2275),
.B(n_133),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_SL g2326 ( 
.A(n_2276),
.B(n_2290),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2312),
.B(n_564),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_R g2328 ( 
.A(n_2278),
.B(n_133),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_R g2329 ( 
.A(n_2283),
.B(n_2300),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2292),
.B(n_564),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2309),
.B(n_591),
.Y(n_2331)
);

NAND2xp33_ASAP7_75t_L g2332 ( 
.A(n_2305),
.B(n_134),
.Y(n_2332)
);

XNOR2xp5_ASAP7_75t_L g2333 ( 
.A(n_2296),
.B(n_135),
.Y(n_2333)
);

NAND3xp33_ASAP7_75t_SL g2334 ( 
.A(n_2282),
.B(n_136),
.C(n_137),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_R g2335 ( 
.A(n_2295),
.B(n_136),
.Y(n_2335)
);

XNOR2xp5_ASAP7_75t_L g2336 ( 
.A(n_2298),
.B(n_138),
.Y(n_2336)
);

NAND2xp33_ASAP7_75t_SL g2337 ( 
.A(n_2299),
.B(n_138),
.Y(n_2337)
);

NAND2xp33_ASAP7_75t_SL g2338 ( 
.A(n_2294),
.B(n_139),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_R g2339 ( 
.A(n_2306),
.B(n_139),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_R g2340 ( 
.A(n_2289),
.B(n_140),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_R g2341 ( 
.A(n_2304),
.B(n_141),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_R g2342 ( 
.A(n_2313),
.B(n_2307),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_2280),
.B(n_591),
.Y(n_2343)
);

NOR3xp33_ASAP7_75t_SL g2344 ( 
.A(n_2311),
.B(n_141),
.C(n_142),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_R g2345 ( 
.A(n_2307),
.B(n_143),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2287),
.B(n_144),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_R g2347 ( 
.A(n_2316),
.B(n_2302),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_R g2348 ( 
.A(n_2302),
.B(n_2303),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_SL g2349 ( 
.A(n_2286),
.B(n_591),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_R g2350 ( 
.A(n_2308),
.B(n_145),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2285),
.B(n_146),
.Y(n_2351)
);

XNOR2xp5_ASAP7_75t_L g2352 ( 
.A(n_2288),
.B(n_147),
.Y(n_2352)
);

NAND2xp33_ASAP7_75t_SL g2353 ( 
.A(n_2315),
.B(n_147),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_R g2354 ( 
.A(n_2291),
.B(n_149),
.Y(n_2354)
);

XNOR2xp5_ASAP7_75t_L g2355 ( 
.A(n_2277),
.B(n_150),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2317),
.B(n_591),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_R g2357 ( 
.A(n_2318),
.B(n_151),
.Y(n_2357)
);

XNOR2xp5_ASAP7_75t_L g2358 ( 
.A(n_2274),
.B(n_151),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2301),
.B(n_653),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_R g2360 ( 
.A(n_2310),
.B(n_152),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_R g2361 ( 
.A(n_2281),
.B(n_155),
.Y(n_2361)
);

OAI31xp33_ASAP7_75t_SL g2362 ( 
.A1(n_2352),
.A2(n_2314),
.A3(n_156),
.B(n_157),
.Y(n_2362)
);

A2O1A1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2325),
.A2(n_155),
.B(n_156),
.C(n_158),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2336),
.Y(n_2364)
);

NOR2x1p5_ASAP7_75t_L g2365 ( 
.A(n_2334),
.B(n_158),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2333),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2324),
.Y(n_2367)
);

NAND3x1_ASAP7_75t_L g2368 ( 
.A(n_2346),
.B(n_159),
.C(n_160),
.Y(n_2368)
);

NAND3x1_ASAP7_75t_L g2369 ( 
.A(n_2351),
.B(n_159),
.C(n_160),
.Y(n_2369)
);

OR2x2_ASAP7_75t_L g2370 ( 
.A(n_2326),
.B(n_162),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_2342),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2350),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2345),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2347),
.B(n_163),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2338),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_L g2376 ( 
.A(n_2337),
.B(n_163),
.Y(n_2376)
);

NOR3xp33_ASAP7_75t_L g2377 ( 
.A(n_2331),
.B(n_164),
.C(n_167),
.Y(n_2377)
);

AND3x1_ASAP7_75t_L g2378 ( 
.A(n_2344),
.B(n_2349),
.C(n_2348),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2355),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2320),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2358),
.Y(n_2381)
);

NOR3xp33_ASAP7_75t_L g2382 ( 
.A(n_2327),
.B(n_164),
.C(n_168),
.Y(n_2382)
);

NAND3xp33_ASAP7_75t_L g2383 ( 
.A(n_2332),
.B(n_653),
.C(n_838),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_2329),
.Y(n_2384)
);

NAND5xp2_ASAP7_75t_L g2385 ( 
.A(n_2354),
.B(n_2357),
.C(n_2328),
.D(n_2335),
.E(n_2360),
.Y(n_2385)
);

XOR2xp5_ASAP7_75t_L g2386 ( 
.A(n_2356),
.B(n_168),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_SL g2387 ( 
.A(n_2330),
.B(n_169),
.C(n_170),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2339),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2353),
.A2(n_653),
.B1(n_838),
.B2(n_860),
.Y(n_2389)
);

NAND2x1p5_ASAP7_75t_L g2390 ( 
.A(n_2371),
.B(n_2359),
.Y(n_2390)
);

NOR2x1_ASAP7_75t_L g2391 ( 
.A(n_2384),
.B(n_2343),
.Y(n_2391)
);

OAI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2372),
.A2(n_2321),
.B1(n_2322),
.B2(n_2341),
.C(n_2323),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2365),
.Y(n_2393)
);

A2O1A1Ixp33_ASAP7_75t_L g2394 ( 
.A1(n_2366),
.A2(n_2340),
.B(n_2361),
.C(n_169),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2373),
.B(n_171),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2388),
.Y(n_2396)
);

CKINVDCx5p33_ASAP7_75t_R g2397 ( 
.A(n_2380),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2375),
.B(n_1890),
.Y(n_2398)
);

NOR3xp33_ASAP7_75t_SL g2399 ( 
.A(n_2385),
.B(n_172),
.C(n_173),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2370),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2374),
.Y(n_2401)
);

INVxp33_ASAP7_75t_L g2402 ( 
.A(n_2376),
.Y(n_2402)
);

CKINVDCx12_ASAP7_75t_R g2403 ( 
.A(n_2364),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2367),
.B(n_1918),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2379),
.B(n_174),
.Y(n_2405)
);

BUFx2_ASAP7_75t_L g2406 ( 
.A(n_2369),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2381),
.Y(n_2407)
);

OAI211xp5_ASAP7_75t_SL g2408 ( 
.A1(n_2362),
.A2(n_653),
.B(n_186),
.C(n_195),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2378),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_2387),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2386),
.Y(n_2411)
);

AOI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2403),
.A2(n_2368),
.B1(n_2377),
.B2(n_2382),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2407),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2406),
.Y(n_2414)
);

OAI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2396),
.A2(n_2383),
.B(n_2389),
.Y(n_2415)
);

NOR2xp67_ASAP7_75t_L g2416 ( 
.A(n_2392),
.B(n_2363),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_2400),
.B(n_2393),
.Y(n_2417)
);

AOI222xp33_ASAP7_75t_L g2418 ( 
.A1(n_2409),
.A2(n_838),
.B1(n_860),
.B2(n_1245),
.C1(n_1475),
.C2(n_1423),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2410),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2390),
.Y(n_2420)
);

NAND3xp33_ASAP7_75t_L g2421 ( 
.A(n_2397),
.B(n_860),
.C(n_1259),
.Y(n_2421)
);

OA21x2_ASAP7_75t_L g2422 ( 
.A1(n_2411),
.A2(n_181),
.B(n_196),
.Y(n_2422)
);

OAI21xp33_ASAP7_75t_L g2423 ( 
.A1(n_2402),
.A2(n_2399),
.B(n_2391),
.Y(n_2423)
);

OAI22x1_ASAP7_75t_L g2424 ( 
.A1(n_2401),
.A2(n_1488),
.B1(n_1480),
.B2(n_1475),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2394),
.A2(n_860),
.B1(n_1451),
.B2(n_1484),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2413),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2417),
.Y(n_2427)
);

OAI22xp5_ASAP7_75t_SL g2428 ( 
.A1(n_2420),
.A2(n_2395),
.B1(n_2405),
.B2(n_2408),
.Y(n_2428)
);

OAI22xp5_ASAP7_75t_SL g2429 ( 
.A1(n_2414),
.A2(n_2405),
.B1(n_2404),
.B2(n_2398),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_2419),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2422),
.Y(n_2431)
);

OAI22xp33_ASAP7_75t_SL g2432 ( 
.A1(n_2412),
.A2(n_198),
.B1(n_199),
.B2(n_203),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2423),
.Y(n_2433)
);

A2O1A1Ixp33_ASAP7_75t_SL g2434 ( 
.A1(n_2415),
.A2(n_1484),
.B(n_1474),
.C(n_1470),
.Y(n_2434)
);

BUFx2_ASAP7_75t_SL g2435 ( 
.A(n_2416),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_2426),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2435),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2427),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2431),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2430),
.Y(n_2440)
);

AND3x4_ASAP7_75t_L g2441 ( 
.A(n_2428),
.B(n_2425),
.C(n_2424),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2440),
.A2(n_2433),
.B1(n_2429),
.B2(n_2432),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2436),
.A2(n_2421),
.B1(n_2434),
.B2(n_2418),
.Y(n_2443)
);

AOI31xp33_ASAP7_75t_L g2444 ( 
.A1(n_2438),
.A2(n_205),
.A3(n_211),
.B(n_212),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_2439),
.A2(n_1465),
.B1(n_1423),
.B2(n_1431),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2442),
.Y(n_2446)
);

HB1xp67_ASAP7_75t_L g2447 ( 
.A(n_2443),
.Y(n_2447)
);

OAI22x1_ASAP7_75t_L g2448 ( 
.A1(n_2444),
.A2(n_2437),
.B1(n_2441),
.B2(n_219),
.Y(n_2448)
);

XNOR2xp5_ASAP7_75t_L g2449 ( 
.A(n_2445),
.B(n_213),
.Y(n_2449)
);

AOI21xp33_ASAP7_75t_SL g2450 ( 
.A1(n_2446),
.A2(n_217),
.B(n_221),
.Y(n_2450)
);

AOI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2447),
.A2(n_1313),
.B(n_1293),
.Y(n_2451)
);

AOI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2448),
.A2(n_1313),
.B1(n_1293),
.B2(n_1290),
.C(n_1263),
.Y(n_2452)
);

AOI22xp33_ASAP7_75t_L g2453 ( 
.A1(n_2452),
.A2(n_2449),
.B1(n_1488),
.B2(n_1480),
.Y(n_2453)
);

AOI222xp33_ASAP7_75t_L g2454 ( 
.A1(n_2450),
.A2(n_2451),
.B1(n_1263),
.B2(n_1313),
.C1(n_1290),
.C2(n_1293),
.Y(n_2454)
);

AOI222xp33_ASAP7_75t_L g2455 ( 
.A1(n_2452),
.A2(n_1263),
.B1(n_1290),
.B2(n_1293),
.C1(n_1313),
.C2(n_1466),
.Y(n_2455)
);

AO21x2_ASAP7_75t_L g2456 ( 
.A1(n_2450),
.A2(n_223),
.B(n_228),
.Y(n_2456)
);

OAI222xp33_ASAP7_75t_L g2457 ( 
.A1(n_2453),
.A2(n_1466),
.B1(n_1465),
.B2(n_1460),
.C1(n_1436),
.C2(n_1431),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2456),
.B(n_229),
.Y(n_2458)
);

XNOR2xp5_ASAP7_75t_L g2459 ( 
.A(n_2454),
.B(n_230),
.Y(n_2459)
);

OAI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2458),
.A2(n_2455),
.B(n_1460),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2460),
.A2(n_2459),
.B1(n_2457),
.B2(n_1290),
.Y(n_2461)
);

AOI221xp5_ASAP7_75t_L g2462 ( 
.A1(n_2461),
.A2(n_1263),
.B1(n_1436),
.B2(n_249),
.C(n_253),
.Y(n_2462)
);

AOI211xp5_ASAP7_75t_L g2463 ( 
.A1(n_2462),
.A2(n_237),
.B(n_239),
.C(n_254),
.Y(n_2463)
);


endmodule