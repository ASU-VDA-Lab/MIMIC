module fake_ibex_1616_n_2387 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_688, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_673, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_679, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_672, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_675, n_463, n_624, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_2387);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_688;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_673;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_679;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_672;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_2387;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_1308;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2151;
wire n_1391;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_876;
wire n_711;
wire n_1840;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_787;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_2090;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_1445;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_745;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_1649;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_1549;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_1040;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_2256;
wire n_737;
wire n_1571;
wire n_1980;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_1591;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_2006;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2358;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_817;
wire n_2193;
wire n_2095;
wire n_951;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_863;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_895;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_972;
wire n_1815;
wire n_1917;
wire n_1444;
wire n_920;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_991;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2344;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_2141;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_1259;
wire n_2108;
wire n_1001;
wire n_2143;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_1124;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_934;
wire n_775;
wire n_950;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_1167;
wire n_818;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_1632;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_1329;
wire n_2337;
wire n_854;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_1092;
wire n_1808;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_918;
wire n_2056;
wire n_1913;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_1472;
wire n_1365;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_866;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_867;
wire n_983;
wire n_1417;
wire n_2282;
wire n_970;
wire n_921;
wire n_1534;
wire n_908;
wire n_1346;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_1854;
wire n_1506;

BUFx3_ASAP7_75t_L g696 ( 
.A(n_207),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_647),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_92),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_636),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_364),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_366),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_299),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_473),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_50),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_375),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_689),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_578),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_660),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_337),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_540),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_597),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_261),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_93),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_47),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_684),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_638),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_662),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_669),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_622),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_29),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_671),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_668),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_49),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_559),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_486),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_531),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_315),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_688),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_282),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_654),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_373),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_489),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_302),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_536),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_419),
.Y(n_736)
);

BUFx10_ASAP7_75t_L g737 ( 
.A(n_47),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_252),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_525),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_692),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_297),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_150),
.Y(n_742)
);

BUFx5_ASAP7_75t_L g743 ( 
.A(n_224),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_670),
.Y(n_744)
);

CKINVDCx16_ASAP7_75t_R g745 ( 
.A(n_650),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_544),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_684),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_62),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_676),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_42),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_352),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_656),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_434),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_440),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_595),
.Y(n_755)
);

CKINVDCx16_ASAP7_75t_R g756 ( 
.A(n_434),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_516),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_372),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_334),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_209),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_588),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_280),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_186),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_300),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_285),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_33),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_105),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_205),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_330),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_121),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_584),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_644),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_629),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_169),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_102),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_160),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_657),
.Y(n_777)
);

BUFx5_ASAP7_75t_L g778 ( 
.A(n_687),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_658),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_312),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_18),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_70),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_225),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_284),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_514),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_133),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_265),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_679),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_340),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_472),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_458),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_46),
.Y(n_792)
);

BUFx5_ASAP7_75t_L g793 ( 
.A(n_39),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_98),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_653),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_601),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_601),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_634),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_594),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_555),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_231),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_624),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_661),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_126),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_320),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_649),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_382),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_659),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_677),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_179),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_556),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_532),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_174),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_150),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_639),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_75),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_333),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_76),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_354),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_461),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_495),
.Y(n_821)
);

BUFx5_ASAP7_75t_L g822 ( 
.A(n_273),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_678),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_69),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_353),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_552),
.Y(n_826)
);

CKINVDCx16_ASAP7_75t_R g827 ( 
.A(n_168),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_631),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_173),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_665),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_5),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_558),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_459),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_597),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_158),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_671),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_557),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_520),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_685),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_674),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_625),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_682),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_643),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_630),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_273),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_172),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_689),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_446),
.Y(n_848)
);

BUFx5_ASAP7_75t_L g849 ( 
.A(n_146),
.Y(n_849)
);

BUFx5_ASAP7_75t_L g850 ( 
.A(n_694),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_321),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_553),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_229),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_641),
.Y(n_854)
);

BUFx5_ASAP7_75t_L g855 ( 
.A(n_582),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_554),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_670),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_591),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_672),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_673),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_643),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_640),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_683),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_691),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_559),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_120),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_278),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_687),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_399),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_646),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_82),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_298),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_526),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_642),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_452),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_107),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_126),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_383),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_101),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_680),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_666),
.Y(n_881)
);

INVxp67_ASAP7_75t_SL g882 ( 
.A(n_85),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_165),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_614),
.Y(n_884)
);

CKINVDCx16_ASAP7_75t_R g885 ( 
.A(n_602),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_397),
.Y(n_886)
);

CKINVDCx16_ASAP7_75t_R g887 ( 
.A(n_599),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_242),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_651),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_590),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_263),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_596),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_328),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_46),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_313),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_464),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_187),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_27),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_158),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_581),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_252),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_144),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_33),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_36),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_626),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_94),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_442),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_227),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_589),
.Y(n_909)
);

CKINVDCx12_ASAP7_75t_R g910 ( 
.A(n_309),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_603),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_253),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_420),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_335),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_645),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_599),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_294),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_119),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_466),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_278),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_389),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_675),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_681),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_627),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_196),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_587),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_531),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_586),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_59),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_516),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_551),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_302),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_65),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_399),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_569),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_693),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_392),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_170),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_365),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_633),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_426),
.Y(n_941)
);

BUFx10_ASAP7_75t_L g942 ( 
.A(n_664),
.Y(n_942)
);

CKINVDCx14_ASAP7_75t_R g943 ( 
.A(n_315),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_279),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_652),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_42),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_137),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_25),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_686),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_628),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_46),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_129),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_462),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_663),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_648),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_593),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_511),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_25),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_374),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_695),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_85),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_693),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_600),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_649),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_611),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_623),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_386),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_632),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_637),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_439),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_477),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_151),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_243),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_667),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_247),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_78),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_644),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_635),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_265),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_666),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_404),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_676),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_199),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_588),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_327),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_84),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_275),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_407),
.Y(n_988)
);

INVxp67_ASAP7_75t_L g989 ( 
.A(n_528),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_655),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_640),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_13),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_660),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_180),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_431),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_532),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_573),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_585),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_148),
.Y(n_999)
);

CKINVDCx14_ASAP7_75t_R g1000 ( 
.A(n_116),
.Y(n_1000)
);

CKINVDCx14_ASAP7_75t_R g1001 ( 
.A(n_474),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_690),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_502),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_95),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_177),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_568),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_274),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_542),
.Y(n_1008)
);

BUFx10_ASAP7_75t_L g1009 ( 
.A(n_580),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_53),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_455),
.Y(n_1011)
);

BUFx5_ASAP7_75t_L g1012 ( 
.A(n_600),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_583),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_698),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_791),
.Y(n_1015)
);

INVxp33_ASAP7_75t_L g1016 ( 
.A(n_701),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_879),
.Y(n_1017)
);

CKINVDCx16_ASAP7_75t_R g1018 ( 
.A(n_756),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_943),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_713),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_906),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_1000),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_876),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_934),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_789),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_759),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_794),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_827),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_813),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_1001),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_910),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_700),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_769),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_907),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_696),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_702),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_709),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_712),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_705),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_784),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_734),
.Y(n_1041)
);

CKINVDCx16_ASAP7_75t_R g1042 ( 
.A(n_716),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_753),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_714),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_706),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_825),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_762),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_764),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_696),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_721),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_724),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_780),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_781),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_945),
.B(n_0),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_914),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_728),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_786),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1012),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_787),
.Y(n_1059)
);

INVxp33_ASAP7_75t_L g1060 ( 
.A(n_965),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_732),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_728),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_737),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_730),
.Y(n_1064)
);

INVxp67_ASAP7_75t_SL g1065 ( 
.A(n_736),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_738),
.Y(n_1066)
);

CKINVDCx16_ASAP7_75t_R g1067 ( 
.A(n_745),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_804),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_807),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_741),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_742),
.Y(n_1071)
);

CKINVDCx16_ASAP7_75t_R g1072 ( 
.A(n_885),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_748),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_820),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_887),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_750),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_754),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_758),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_778),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_833),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_815),
.B(n_0),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_838),
.B(n_1),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_938),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_760),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_948),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_859),
.B(n_1),
.Y(n_1086)
);

INVx6_ASAP7_75t_L g1087 ( 
.A(n_1045),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_1063),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1035),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_1064),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_1034),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_1063),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1058),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1034),
.B(n_1049),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1016),
.B(n_737),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1014),
.B(n_788),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1020),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1056),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1060),
.B(n_816),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1065),
.Y(n_1100)
);

OA21x2_ASAP7_75t_L g1101 ( 
.A1(n_1079),
.A2(n_1038),
.B(n_1037),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1065),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1023),
.B(n_911),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1015),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1049),
.B(n_766),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1017),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_1021),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1062),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1064),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1018),
.A2(n_768),
.B1(n_770),
.B2(n_767),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_1064),
.Y(n_1111)
);

CKINVDCx8_ASAP7_75t_R g1112 ( 
.A(n_1025),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1041),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1032),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1043),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1047),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1048),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1052),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1036),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1053),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1057),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1059),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1028),
.B(n_763),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1022),
.B(n_775),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1027),
.B(n_776),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1068),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1029),
.B(n_763),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1024),
.B(n_727),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1069),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1074),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1080),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1081),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1082),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1086),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1054),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1039),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1042),
.B(n_810),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1044),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1050),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1051),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1061),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1066),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1070),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_1071),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1073),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1031),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1076),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_1077),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1078),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1084),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1030),
.B(n_782),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1075),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1026),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1033),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1040),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1046),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1055),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1085),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1083),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1020),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1016),
.B(n_810),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1014),
.B(n_989),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1064),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1035),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1035),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1058),
.A2(n_783),
.B(n_751),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1034),
.B(n_792),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1034),
.B(n_755),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1064),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1034),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1035),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1063),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1063),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1035),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1034),
.B(n_812),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1063),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1064),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1034),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1016),
.B(n_848),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1064),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1034),
.B(n_805),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1058),
.A2(n_783),
.B(n_751),
.Y(n_1183)
);

AND2x6_ASAP7_75t_L g1184 ( 
.A(n_1063),
.B(n_848),
.Y(n_1184)
);

CKINVDCx8_ASAP7_75t_R g1185 ( 
.A(n_1018),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_L g1186 ( 
.A(n_1019),
.B(n_743),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1035),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1035),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1020),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1063),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1064),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1064),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1035),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1035),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1045),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1035),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1026),
.A2(n_1007),
.B1(n_729),
.B2(n_777),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1045),
.Y(n_1198)
);

INVxp33_ASAP7_75t_SL g1199 ( 
.A(n_1019),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1018),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1035),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1064),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1063),
.B(n_743),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1035),
.Y(n_1204)
);

AND2x6_ASAP7_75t_L g1205 ( 
.A(n_1063),
.B(n_921),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1035),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1020),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1016),
.B(n_814),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1091),
.B(n_1171),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1101),
.Y(n_1210)
);

AND3x2_ASAP7_75t_L g1211 ( 
.A(n_1097),
.B(n_1208),
.C(n_1161),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1094),
.B(n_743),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1104),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1167),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_SL g1215 ( 
.A(n_1159),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1107),
.Y(n_1216)
);

BUFx4f_ASAP7_75t_L g1217 ( 
.A(n_1147),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1091),
.A2(n_818),
.B1(n_819),
.B2(n_817),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1132),
.B(n_824),
.Y(n_1219)
);

AND2x6_ASAP7_75t_L g1220 ( 
.A(n_1102),
.B(n_944),
.Y(n_1220)
);

BUFx4f_ASAP7_75t_L g1221 ( 
.A(n_1147),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1189),
.B(n_704),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1183),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1207),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_1171),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1197),
.B(n_882),
.C(n_765),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1162),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1126),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_1200),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1133),
.B(n_829),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1179),
.B(n_831),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1180),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1184),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1122),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1089),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1122),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1092),
.B(n_835),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1112),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1087),
.Y(n_1239)
);

AND2x6_ASAP7_75t_L g1240 ( 
.A(n_1123),
.B(n_944),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1129),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1105),
.B(n_793),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1098),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1184),
.Y(n_1244)
);

INVxp33_ASAP7_75t_L g1245 ( 
.A(n_1095),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1168),
.B(n_801),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1131),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1173),
.B(n_846),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1099),
.Y(n_1249)
);

AND2x6_ASAP7_75t_L g1250 ( 
.A(n_1100),
.B(n_1010),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1165),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1205),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1141),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1088),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1135),
.A2(n_1172),
.B1(n_1175),
.B2(n_1166),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1187),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1188),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1185),
.Y(n_1258)
);

INVx4_ASAP7_75t_SL g1259 ( 
.A(n_1137),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1182),
.B(n_845),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1193),
.Y(n_1261)
);

CKINVDCx6p67_ASAP7_75t_R g1262 ( 
.A(n_1159),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_1174),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1194),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_L g1265 ( 
.A(n_1146),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1196),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1201),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1103),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1204),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1142),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1114),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1206),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1169),
.Y(n_1273)
);

INVx5_ASAP7_75t_L g1274 ( 
.A(n_1177),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1143),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1108),
.B(n_793),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1190),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1119),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1150),
.Y(n_1279)
);

BUFx4f_ASAP7_75t_L g1280 ( 
.A(n_1144),
.Y(n_1280)
);

NOR3xp33_ASAP7_75t_L g1281 ( 
.A(n_1110),
.B(n_894),
.C(n_869),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1116),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1154),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1127),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1195),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1176),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_R g1287 ( 
.A(n_1199),
.B(n_866),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1124),
.B(n_939),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1115),
.A2(n_871),
.B1(n_872),
.B2(n_851),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1152),
.B(n_867),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_L g1291 ( 
.A(n_1153),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1157),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1113),
.B(n_822),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1125),
.B(n_961),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1198),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1149),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1117),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1155),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1148),
.B(n_961),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1156),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1128),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1128),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_L g1303 ( 
.A(n_1136),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1134),
.B(n_891),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1158),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1118),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1120),
.B(n_1005),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1121),
.A2(n_875),
.B1(n_878),
.B2(n_877),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1130),
.B(n_1011),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1138),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1093),
.A2(n_883),
.B1(n_888),
.B2(n_886),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1096),
.B(n_849),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1203),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1139),
.B(n_893),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1163),
.B(n_849),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1140),
.B(n_895),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1186),
.B(n_902),
.C(n_897),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1145),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1160),
.B(n_1151),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1090),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1090),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1109),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1111),
.B(n_730),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1202),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1164),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1178),
.B(n_697),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1178),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1181),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1181),
.Y(n_1330)
);

AND2x6_ASAP7_75t_L g1331 ( 
.A(n_1191),
.B(n_730),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1192),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1202),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

AND2x6_ASAP7_75t_L g1335 ( 
.A(n_1102),
.B(n_730),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1097),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1102),
.A2(n_899),
.B1(n_901),
.B2(n_898),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1106),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1167),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1167),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1091),
.B(n_746),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_SL g1342 ( 
.A(n_1112),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_1184),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1094),
.B(n_849),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1091),
.B(n_746),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1184),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1101),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1097),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1189),
.Y(n_1349)
);

XOR2x2_ASAP7_75t_SL g1350 ( 
.A(n_1110),
.B(n_795),
.Y(n_1350)
);

INVx8_ASAP7_75t_L g1351 ( 
.A(n_1215),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1245),
.B(n_925),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1348),
.Y(n_1353)
);

O2A1O1Ixp5_ASAP7_75t_L g1354 ( 
.A1(n_1294),
.A2(n_908),
.B(n_912),
.C(n_904),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1255),
.B(n_929),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1219),
.B(n_932),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1233),
.B(n_937),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1224),
.B(n_802),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1282),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1230),
.B(n_951),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1347),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1214),
.A2(n_1334),
.B(n_1223),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1222),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1235),
.A2(n_837),
.B1(n_840),
.B2(n_828),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1244),
.B(n_1252),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1249),
.B(n_970),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1209),
.A2(n_981),
.B1(n_985),
.B2(n_976),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1218),
.A2(n_987),
.B1(n_988),
.B2(n_986),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1252),
.B(n_999),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1279),
.A2(n_884),
.B1(n_889),
.B2(n_865),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_SL g1372 ( 
.A(n_1239),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1343),
.B(n_1346),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1243),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1227),
.A2(n_707),
.B1(n_711),
.B2(n_708),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1251),
.B(n_1004),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1256),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1257),
.B(n_1261),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1264),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1266),
.B(n_1267),
.Y(n_1380)
);

INVxp33_ASAP7_75t_SL g1381 ( 
.A(n_1296),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1271),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1341),
.B(n_1345),
.Y(n_1383)
);

AND2x6_ASAP7_75t_L g1384 ( 
.A(n_1318),
.B(n_774),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1242),
.A2(n_917),
.B(n_913),
.Y(n_1385)
);

OAI22x1_ASAP7_75t_L g1386 ( 
.A1(n_1350),
.A2(n_719),
.B1(n_720),
.B2(n_718),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1269),
.B(n_1272),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1290),
.B(n_918),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1284),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1306),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1220),
.B(n_920),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1270),
.B(n_790),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1232),
.A2(n_725),
.B1(n_726),
.B2(n_722),
.Y(n_1393)
);

NOR3xp33_ASAP7_75t_L g1394 ( 
.A(n_1226),
.B(n_881),
.C(n_880),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1220),
.B(n_933),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1298),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1262),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1339),
.A2(n_947),
.B(n_946),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1211),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1338),
.B(n_952),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1337),
.A2(n_958),
.B1(n_959),
.B2(n_953),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1285),
.Y(n_1402)
);

INVx8_ASAP7_75t_L g1403 ( 
.A(n_1240),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1212),
.A2(n_973),
.B(n_975),
.C(n_967),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1281),
.B(n_1316),
.C(n_1314),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1344),
.A2(n_983),
.B(n_992),
.C(n_979),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1292),
.B(n_1002),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1303),
.B(n_735),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1295),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1310),
.B(n_739),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1268),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1250),
.B(n_994),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1250),
.B(n_995),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1278),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1297),
.B(n_747),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1275),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1340),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1287),
.Y(n_1418)
);

AND2x6_ASAP7_75t_L g1419 ( 
.A(n_1258),
.B(n_774),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1259),
.B(n_699),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1323),
.Y(n_1421)
);

INVx8_ASAP7_75t_L g1422 ( 
.A(n_1240),
.Y(n_1422)
);

A2O1A1Ixp33_ASAP7_75t_L g1423 ( 
.A1(n_1276),
.A2(n_717),
.B(n_723),
.C(n_715),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_SL g1424 ( 
.A(n_1229),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1283),
.B(n_773),
.C(n_772),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1308),
.B(n_796),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1238),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1248),
.Y(n_1428)
);

NAND2x1_ASAP7_75t_L g1429 ( 
.A(n_1335),
.B(n_774),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1273),
.A2(n_803),
.B1(n_806),
.B2(n_800),
.Y(n_1430)
);

AND2x6_ASAP7_75t_SL g1431 ( 
.A(n_1342),
.B(n_731),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1280),
.B(n_808),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1237),
.B(n_1305),
.C(n_1289),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1217),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1323),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1221),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1323),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1319),
.A2(n_740),
.B1(n_744),
.B2(n_733),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1286),
.B(n_811),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1293),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1300),
.B(n_2),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1246),
.A2(n_752),
.B(n_771),
.C(n_749),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1311),
.B(n_826),
.C(n_823),
.Y(n_1443)
);

AND2x2_ASAP7_75t_SL g1444 ( 
.A(n_1265),
.B(n_703),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1286),
.B(n_839),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1291),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1260),
.B(n_843),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1228),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1213),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1216),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1307),
.B(n_1309),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1288),
.B(n_856),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1317),
.B(n_857),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1301),
.A2(n_1013),
.B1(n_860),
.B2(n_862),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1302),
.B(n_858),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1327),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1312),
.B(n_863),
.Y(n_1457)
);

NOR3xp33_ASAP7_75t_L g1458 ( 
.A(n_1304),
.B(n_1254),
.C(n_1277),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1315),
.B(n_864),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1263),
.B(n_779),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1263),
.B(n_868),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1299),
.A2(n_797),
.B1(n_798),
.B2(n_785),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1274),
.B(n_870),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1234),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1313),
.B(n_873),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1236),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1241),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1327),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1247),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1321),
.B(n_890),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1324),
.B(n_892),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1326),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1328),
.A2(n_809),
.B(n_821),
.C(n_799),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1329),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1322),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1331),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1330),
.A2(n_832),
.B(n_834),
.C(n_830),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1333),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1320),
.B(n_900),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1332),
.A2(n_896),
.B1(n_903),
.B2(n_853),
.Y(n_1480)
);

INVx8_ASAP7_75t_L g1481 ( 
.A(n_1325),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1225),
.A2(n_919),
.B1(n_922),
.B2(n_915),
.C(n_909),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1255),
.B(n_924),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1348),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1231),
.B(n_926),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1255),
.B(n_927),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1231),
.B(n_928),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1255),
.B(n_930),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1255),
.B(n_935),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1210),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1255),
.B(n_936),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1336),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1210),
.Y(n_1493)
);

BUFx5_ASAP7_75t_L g1494 ( 
.A(n_1323),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1231),
.B(n_949),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1255),
.B(n_950),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1349),
.B(n_3),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1255),
.B(n_954),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1231),
.A2(n_956),
.B1(n_960),
.B2(n_955),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1255),
.B(n_964),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1255),
.B(n_966),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1231),
.A2(n_969),
.B1(n_971),
.B2(n_968),
.Y(n_1502)
);

INVxp67_ASAP7_75t_L g1503 ( 
.A(n_1224),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1253),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1255),
.B(n_974),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1224),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1231),
.A2(n_978),
.B1(n_982),
.B2(n_977),
.Y(n_1507)
);

NAND3x1_ASAP7_75t_L g1508 ( 
.A(n_1226),
.B(n_842),
.C(n_841),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1255),
.B(n_984),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1231),
.B(n_991),
.C(n_990),
.Y(n_1510)
);

NOR2xp67_ASAP7_75t_L g1511 ( 
.A(n_1349),
.B(n_4),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1255),
.B(n_993),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1381),
.B(n_997),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1351),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1362),
.A2(n_847),
.B(n_844),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1417),
.A2(n_854),
.B(n_852),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1363),
.B(n_996),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1351),
.Y(n_1518)
);

NAND2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1504),
.B(n_853),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1377),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1379),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1383),
.B(n_916),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1389),
.B(n_923),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1398),
.A2(n_940),
.B(n_931),
.Y(n_1524)
);

NOR3xp33_ASAP7_75t_L g1525 ( 
.A(n_1433),
.B(n_963),
.C(n_962),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1369),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1378),
.B(n_980),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1394),
.A2(n_1009),
.B1(n_942),
.B2(n_941),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1369),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1405),
.A2(n_998),
.B(n_1003),
.C(n_957),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1354),
.A2(n_1008),
.B(n_1006),
.C(n_757),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1380),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1406),
.A2(n_757),
.B(n_761),
.C(n_710),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1358),
.B(n_761),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1414),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1387),
.B(n_836),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1388),
.B(n_905),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1396),
.A2(n_855),
.B1(n_1012),
.B2(n_850),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1440),
.A2(n_855),
.B(n_850),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1428),
.B(n_5),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1385),
.A2(n_972),
.B(n_861),
.C(n_874),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1371),
.A2(n_1012),
.B1(n_855),
.B2(n_972),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1369),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1359),
.A2(n_5),
.B(n_6),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1403),
.Y(n_1546)
);

BUFx4f_ASAP7_75t_L g1547 ( 
.A(n_1403),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1386),
.A2(n_874),
.B1(n_861),
.B2(n_8),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1484),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_L g1550 ( 
.A(n_1434),
.B(n_874),
.Y(n_1550)
);

AOI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1410),
.A2(n_874),
.B(n_6),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1361),
.A2(n_7),
.B(n_9),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1490),
.A2(n_9),
.B(n_10),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1493),
.A2(n_11),
.B(n_12),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1492),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1423),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1441),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1442),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1465),
.A2(n_22),
.B(n_23),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1364),
.B(n_24),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1451),
.B(n_24),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1376),
.A2(n_26),
.B(n_27),
.Y(n_1562)
);

AO22x1_ASAP7_75t_L g1563 ( 
.A1(n_1419),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_1563)
);

AOI21xp33_ASAP7_75t_L g1564 ( 
.A1(n_1352),
.A2(n_28),
.B(n_29),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1422),
.B(n_30),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1392),
.B(n_32),
.Y(n_1566)
);

OAI21xp33_ASAP7_75t_L g1567 ( 
.A1(n_1356),
.A2(n_31),
.B(n_32),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1457),
.A2(n_34),
.B(n_35),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1459),
.A2(n_34),
.B(n_35),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1451),
.B(n_35),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1360),
.A2(n_37),
.B(n_38),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1415),
.A2(n_38),
.B(n_39),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1473),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1422),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1372),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1397),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1454),
.B(n_45),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1510),
.B(n_45),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1438),
.A2(n_47),
.B(n_44),
.C(n_45),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1444),
.B(n_48),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_L g1581 ( 
.A(n_1494),
.B(n_52),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1355),
.B(n_51),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1427),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1497),
.B(n_53),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1511),
.B(n_54),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1483),
.B(n_54),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1486),
.B(n_55),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1400),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1488),
.B(n_57),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1489),
.B(n_58),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1491),
.B(n_58),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1478),
.A2(n_58),
.B(n_59),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1407),
.B(n_59),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1391),
.A2(n_60),
.B(n_61),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1368),
.B(n_1499),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1395),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1477),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1502),
.B(n_67),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1421),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1366),
.B(n_66),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1456),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1496),
.B(n_1498),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1448),
.A2(n_1450),
.B(n_1449),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1468),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1482),
.B(n_68),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1446),
.B(n_69),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1418),
.B(n_70),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1425),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1609)
);

AND2x4_ASAP7_75t_SL g1610 ( 
.A(n_1436),
.B(n_74),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1505),
.B(n_77),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1402),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1509),
.B(n_79),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1512),
.B(n_79),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1409),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1464),
.A2(n_1467),
.B(n_1466),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1426),
.B(n_1367),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1412),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1413),
.A2(n_1443),
.B(n_1401),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1462),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1447),
.A2(n_83),
.B(n_84),
.Y(n_1621)
);

NOR2xp67_ASAP7_75t_L g1622 ( 
.A(n_1436),
.B(n_1399),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1475),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1460),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1469),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1384),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1507),
.B(n_86),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1452),
.A2(n_87),
.B(n_88),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1485),
.B(n_89),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1416),
.B(n_91),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_R g1631 ( 
.A(n_1431),
.B(n_90),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1453),
.A2(n_94),
.B(n_95),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1480),
.B(n_95),
.C(n_96),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1429),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1487),
.B(n_96),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1435),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1474),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1495),
.B(n_97),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1420),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1437),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1375),
.B(n_99),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1393),
.B(n_99),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1420),
.B(n_100),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1508),
.A2(n_102),
.B(n_103),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1365),
.A2(n_102),
.B(n_103),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1458),
.B(n_104),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1373),
.A2(n_106),
.B(n_107),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1437),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1470),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1430),
.B(n_108),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1357),
.A2(n_108),
.B(n_109),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1439),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1445),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1479),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1370),
.A2(n_110),
.B(n_111),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1455),
.B(n_112),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1471),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1463),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1476),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1408),
.B(n_115),
.C(n_114),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1411),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1461),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1419),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1472),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1432),
.Y(n_1665)
);

OR2x6_ASAP7_75t_L g1666 ( 
.A(n_1481),
.B(n_116),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1481),
.B(n_117),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1381),
.B(n_118),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1390),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1390),
.Y(n_1670)
);

NOR3xp33_ASAP7_75t_L g1671 ( 
.A(n_1433),
.B(n_124),
.C(n_123),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1403),
.B(n_122),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1381),
.B(n_123),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1363),
.B(n_125),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1403),
.B(n_127),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1362),
.A2(n_127),
.B(n_128),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1390),
.Y(n_1677)
);

NOR2xp67_ASAP7_75t_R g1678 ( 
.A(n_1504),
.B(n_130),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1405),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1362),
.A2(n_134),
.B(n_135),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1378),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1504),
.B(n_137),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1381),
.B(n_138),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1381),
.B(n_139),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1351),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1362),
.A2(n_138),
.B(n_139),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1381),
.B(n_140),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1504),
.B(n_140),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1363),
.B(n_141),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1381),
.B(n_142),
.Y(n_1690)
);

CKINVDCx8_ASAP7_75t_R g1691 ( 
.A(n_1351),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1404),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1403),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1390),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1398),
.A2(n_146),
.B(n_147),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1369),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1381),
.B(n_148),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1398),
.A2(n_149),
.B(n_151),
.Y(n_1698)
);

AND2x2_ASAP7_75t_SL g1699 ( 
.A(n_1504),
.B(n_149),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1390),
.Y(n_1700)
);

NAND2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1504),
.B(n_152),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1405),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_1702)
);

NOR3xp33_ASAP7_75t_L g1703 ( 
.A(n_1433),
.B(n_156),
.C(n_155),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1403),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1381),
.B(n_154),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1353),
.B(n_155),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1405),
.B(n_157),
.C(n_159),
.Y(n_1707)
);

BUFx4f_ASAP7_75t_L g1708 ( 
.A(n_1351),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1363),
.B(n_160),
.Y(n_1709)
);

BUFx4f_ASAP7_75t_L g1710 ( 
.A(n_1351),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1390),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1374),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1421),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1362),
.A2(n_161),
.B(n_162),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1363),
.B(n_163),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1381),
.B(n_163),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1362),
.A2(n_164),
.B(n_165),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1353),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1363),
.B(n_166),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1363),
.B(n_167),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1369),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1398),
.A2(n_167),
.B(n_168),
.Y(n_1722)
);

CKINVDCx10_ASAP7_75t_R g1723 ( 
.A(n_1424),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1353),
.B(n_167),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1363),
.B(n_168),
.Y(n_1725)
);

NOR2x1_ASAP7_75t_R g1726 ( 
.A(n_1484),
.B(n_169),
.Y(n_1726)
);

A2O1A1Ixp33_ASAP7_75t_L g1727 ( 
.A1(n_1405),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_1727)
);

CKINVDCx14_ASAP7_75t_R g1728 ( 
.A(n_1353),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1362),
.A2(n_175),
.B(n_176),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1421),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1353),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1381),
.B(n_175),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1363),
.B(n_178),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_1353),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1398),
.A2(n_181),
.B(n_182),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1390),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1381),
.B(n_181),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1382),
.B(n_183),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1363),
.B(n_184),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1363),
.B(n_185),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1374),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1383),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1363),
.B(n_188),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1398),
.A2(n_189),
.B(n_190),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1363),
.B(n_191),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1506),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1381),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1383),
.A2(n_195),
.B1(n_192),
.B2(n_194),
.Y(n_1748)
);

AO22x1_ASAP7_75t_L g1749 ( 
.A1(n_1381),
.A2(n_197),
.B1(n_198),
.B2(n_196),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1398),
.A2(n_200),
.B(n_201),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1504),
.B(n_201),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1363),
.B(n_202),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1363),
.B(n_203),
.Y(n_1753)
);

O2A1O1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1404),
.A2(n_205),
.B(n_203),
.C(n_204),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1381),
.B(n_205),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1381),
.B(n_206),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1506),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1421),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1381),
.B(n_208),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1506),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1381),
.B(n_210),
.Y(n_1761)
);

NAND2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1504),
.B(n_210),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1381),
.B(n_212),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1405),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1363),
.B(n_214),
.Y(n_1765)
);

AND3x2_ASAP7_75t_L g1766 ( 
.A(n_1414),
.B(n_214),
.C(n_215),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1381),
.B(n_216),
.Y(n_1767)
);

O2A1O1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1404),
.A2(n_217),
.B(n_215),
.C(n_216),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1404),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1363),
.B(n_218),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1363),
.B(n_219),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1631),
.B(n_220),
.C(n_221),
.Y(n_1772)
);

CKINVDCx6p67_ASAP7_75t_R g1773 ( 
.A(n_1723),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1691),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1708),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_R g1776 ( 
.A(n_1708),
.B(n_222),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1699),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1602),
.A2(n_223),
.B(n_224),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1609),
.A2(n_226),
.B(n_227),
.Y(n_1779)
);

O2A1O1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1530),
.A2(n_229),
.B(n_226),
.C(n_228),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1532),
.B(n_228),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1540),
.A2(n_228),
.B(n_230),
.Y(n_1782)
);

OR2x6_ASAP7_75t_L g1783 ( 
.A(n_1565),
.B(n_230),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1712),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1583),
.B(n_232),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1710),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1595),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1666),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1666),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1685),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1531),
.A2(n_238),
.B(n_239),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1535),
.B(n_239),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1520),
.B(n_240),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1521),
.B(n_240),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1728),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1669),
.B(n_241),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1581),
.A2(n_241),
.B(n_242),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1537),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1580),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1670),
.B(n_243),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1757),
.B(n_244),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1616),
.A2(n_245),
.B(n_246),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1741),
.Y(n_1803)
);

A2O1A1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1571),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1677),
.B(n_248),
.Y(n_1805)
);

A2O1A1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1568),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1538),
.A2(n_249),
.B(n_250),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1569),
.A2(n_254),
.B(n_251),
.C(n_253),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1666),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1746),
.B(n_254),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1513),
.B(n_254),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1694),
.B(n_255),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1700),
.B(n_256),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1565),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1673),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1711),
.B(n_257),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1718),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1736),
.B(n_257),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1683),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_SL g1820 ( 
.A1(n_1542),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_1820)
);

BUFx12f_ASAP7_75t_L g1821 ( 
.A(n_1731),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1657),
.B(n_261),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1575),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_SL g1824 ( 
.A(n_1734),
.B(n_262),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1760),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1546),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1636),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1559),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1541),
.B(n_264),
.Y(n_1829)
);

A2O1A1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1572),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_1830)
);

OAI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1593),
.A2(n_266),
.B(n_267),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1693),
.B(n_267),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1549),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1649),
.B(n_268),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1704),
.B(n_268),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1704),
.Y(n_1836)
);

OR2x6_ASAP7_75t_L g1837 ( 
.A(n_1672),
.B(n_269),
.Y(n_1837)
);

OAI21xp33_ASAP7_75t_L g1838 ( 
.A1(n_1567),
.A2(n_269),
.B(n_270),
.Y(n_1838)
);

AOI22x1_ASAP7_75t_L g1839 ( 
.A1(n_1519),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1601),
.B(n_270),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1636),
.Y(n_1841)
);

OR2x6_ASAP7_75t_L g1842 ( 
.A(n_1672),
.B(n_1675),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1682),
.B(n_467),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1551),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1536),
.A2(n_277),
.B(n_279),
.Y(n_1845)
);

OAI22x1_ASAP7_75t_SL g1846 ( 
.A1(n_1514),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_1846)
);

BUFx12f_ASAP7_75t_L g1847 ( 
.A(n_1518),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1675),
.B(n_280),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1687),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1659),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1675),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1534),
.B(n_286),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1617),
.B(n_287),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1601),
.B(n_288),
.Y(n_1854)
);

AND2x6_ASAP7_75t_L g1855 ( 
.A(n_1663),
.B(n_288),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1555),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1733),
.B(n_289),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1547),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_SL g1859 ( 
.A1(n_1605),
.A2(n_1703),
.B(n_1671),
.C(n_1698),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1586),
.A2(n_289),
.B(n_290),
.Y(n_1860)
);

OR2x6_ASAP7_75t_L g1861 ( 
.A(n_1701),
.B(n_290),
.Y(n_1861)
);

OR2x6_ASAP7_75t_L g1862 ( 
.A(n_1762),
.B(n_291),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1604),
.B(n_291),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1561),
.B(n_291),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1587),
.A2(n_292),
.B(n_293),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1589),
.A2(n_292),
.B(n_293),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1533),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1682),
.B(n_468),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1561),
.B(n_295),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1590),
.A2(n_296),
.B(n_298),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1603),
.B(n_298),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1688),
.B(n_468),
.Y(n_1872)
);

OR2x6_ASAP7_75t_L g1873 ( 
.A(n_1688),
.B(n_300),
.Y(n_1873)
);

INVx5_ASAP7_75t_L g1874 ( 
.A(n_1663),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1591),
.A2(n_301),
.B(n_302),
.Y(n_1875)
);

BUFx12f_ASAP7_75t_L g1876 ( 
.A(n_1576),
.Y(n_1876)
);

O2A1O1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1597),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1668),
.B(n_303),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1600),
.B(n_304),
.Y(n_1879)
);

O2A1O1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1684),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_1880)
);

AND2x4_ASAP7_75t_SL g1881 ( 
.A(n_1751),
.B(n_308),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1751),
.B(n_469),
.Y(n_1882)
);

AND2x2_ASAP7_75t_SL g1883 ( 
.A(n_1610),
.B(n_310),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1690),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1611),
.A2(n_311),
.B(n_313),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1619),
.A2(n_311),
.B(n_314),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1697),
.A2(n_1716),
.B1(n_1732),
.B2(n_1705),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1738),
.B(n_469),
.Y(n_1888)
);

AO21x1_ASAP7_75t_L g1889 ( 
.A1(n_1545),
.A2(n_471),
.B(n_470),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1613),
.A2(n_316),
.B(n_317),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1747),
.A2(n_1527),
.B1(n_1543),
.B2(n_1606),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1755),
.B(n_317),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1614),
.A2(n_318),
.B(n_319),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1756),
.B(n_318),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1560),
.B(n_318),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1650),
.B(n_319),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1582),
.A2(n_320),
.B(n_321),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_SL g1898 ( 
.A(n_1644),
.B(n_320),
.C(n_321),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1612),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1615),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1692),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1515),
.A2(n_323),
.B(n_325),
.Y(n_1902)
);

AOI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1737),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1525),
.B(n_326),
.Y(n_1904)
);

OR2x6_ASAP7_75t_L g1905 ( 
.A(n_1563),
.B(n_329),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1528),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_1906)
);

OR2x6_ASAP7_75t_SL g1907 ( 
.A(n_1726),
.B(n_331),
.Y(n_1907)
);

O2A1O1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1763),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1664),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1622),
.B(n_335),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1767),
.B(n_336),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1759),
.B(n_473),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1624),
.B(n_337),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1625),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1729),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1761),
.A2(n_341),
.B1(n_338),
.B2(n_339),
.Y(n_1916)
);

A2O1A1Ixp33_ASAP7_75t_SL g1917 ( 
.A1(n_1695),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1522),
.B(n_344),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1639),
.B(n_1618),
.Y(n_1919)
);

OA22x2_ASAP7_75t_L g1920 ( 
.A1(n_1766),
.A2(n_347),
.B1(n_345),
.B2(n_346),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1674),
.B(n_345),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1526),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1637),
.B(n_346),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1517),
.B(n_348),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_SL g1925 ( 
.A1(n_1557),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1665),
.B(n_1689),
.Y(n_1926)
);

A2O1A1Ixp33_ASAP7_75t_SL g1927 ( 
.A1(n_1722),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1664),
.Y(n_1928)
);

OAI21xp33_ASAP7_75t_SL g1929 ( 
.A1(n_1553),
.A2(n_352),
.B(n_354),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1588),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1524),
.A2(n_355),
.B(n_356),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_R g1932 ( 
.A(n_1713),
.B(n_356),
.Y(n_1932)
);

BUFx2_ASAP7_75t_SL g1933 ( 
.A(n_1566),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_R g1934 ( 
.A(n_1713),
.B(n_356),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1749),
.B(n_357),
.Y(n_1935)
);

NOR3xp33_ASAP7_75t_L g1936 ( 
.A(n_1579),
.B(n_1564),
.C(n_1707),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1678),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1709),
.B(n_357),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_SL g1939 ( 
.A1(n_1735),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_1939)
);

CKINVDCx11_ASAP7_75t_R g1940 ( 
.A(n_1646),
.Y(n_1940)
);

BUFx2_ASAP7_75t_L g1941 ( 
.A(n_1526),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1715),
.B(n_358),
.Y(n_1942)
);

INVx2_ASAP7_75t_SL g1943 ( 
.A(n_1550),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1730),
.B(n_475),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1719),
.B(n_360),
.Y(n_1945)
);

INVx3_ASAP7_75t_SL g1946 ( 
.A(n_1730),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1720),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1725),
.B(n_363),
.Y(n_1948)
);

NOR2x1_ASAP7_75t_L g1949 ( 
.A(n_1706),
.B(n_364),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1584),
.A2(n_365),
.B(n_366),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1585),
.A2(n_367),
.B(n_368),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1529),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1656),
.A2(n_368),
.B(n_369),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1662),
.B(n_369),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1654),
.B(n_369),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1577),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_1956)
);

INVx5_ASAP7_75t_L g1957 ( 
.A(n_1758),
.Y(n_1957)
);

NOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1724),
.B(n_370),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1598),
.A2(n_373),
.B(n_374),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1660),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1739),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1667),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1740),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1743),
.B(n_378),
.Y(n_1964)
);

AO22x1_ASAP7_75t_L g1965 ( 
.A1(n_1574),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1745),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1661),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1529),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1643),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1752),
.B(n_384),
.Y(n_1970)
);

INVx4_ASAP7_75t_L g1971 ( 
.A(n_1544),
.Y(n_1971)
);

NAND2xp33_ASAP7_75t_SL g1972 ( 
.A(n_1548),
.B(n_385),
.Y(n_1972)
);

INVx5_ASAP7_75t_L g1973 ( 
.A(n_1544),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1753),
.A2(n_390),
.B1(n_387),
.B2(n_388),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1696),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1676),
.A2(n_390),
.B(n_391),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1516),
.A2(n_392),
.B(n_393),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1721),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1765),
.B(n_393),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1630),
.B(n_394),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1770),
.B(n_395),
.Y(n_1981)
);

A2O1A1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1754),
.A2(n_397),
.B(n_395),
.C(n_396),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1623),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1771),
.B(n_1570),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1607),
.A2(n_399),
.B1(n_396),
.B2(n_398),
.Y(n_1985)
);

INVx1_ASAP7_75t_SL g1986 ( 
.A(n_1652),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1681),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1680),
.A2(n_398),
.B(n_400),
.Y(n_1988)
);

O2A1O1Ixp33_ASAP7_75t_SL g1989 ( 
.A1(n_1744),
.A2(n_401),
.B(n_398),
.C(n_400),
.Y(n_1989)
);

OR2x6_ASAP7_75t_L g1990 ( 
.A(n_1620),
.B(n_401),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1641),
.B(n_401),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1686),
.A2(n_402),
.B(n_403),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1653),
.B(n_403),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1642),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1750),
.B(n_476),
.Y(n_1995)
);

OAI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1742),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1768),
.A2(n_411),
.B(n_409),
.C(n_410),
.Y(n_1997)
);

A2O1A1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1769),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1523),
.B(n_412),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1627),
.B(n_412),
.Y(n_2000)
);

O2A1O1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1558),
.A2(n_1658),
.B(n_1556),
.C(n_1573),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1748),
.B(n_414),
.Y(n_2002)
);

INVxp67_ASAP7_75t_SL g2003 ( 
.A(n_1655),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1608),
.B(n_415),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1596),
.Y(n_2005)
);

A2O1A1Ixp33_ASAP7_75t_L g2006 ( 
.A1(n_1621),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1594),
.B(n_418),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1562),
.B(n_420),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1876),
.Y(n_2009)
);

OR2x6_ASAP7_75t_L g2010 ( 
.A(n_1842),
.B(n_1651),
.Y(n_2010)
);

OAI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1842),
.A2(n_1764),
.B1(n_1679),
.B2(n_1727),
.Y(n_2011)
);

INVx4_ASAP7_75t_SL g2012 ( 
.A(n_1783),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1837),
.A2(n_1702),
.B1(n_1633),
.B2(n_1539),
.Y(n_2013)
);

OAI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_1887),
.A2(n_1635),
.B(n_1629),
.Y(n_2014)
);

NOR2xp67_ASAP7_75t_L g2015 ( 
.A(n_1858),
.B(n_1638),
.Y(n_2015)
);

OAI22x1_ASAP7_75t_L g2016 ( 
.A1(n_1848),
.A2(n_1578),
.B1(n_1633),
.B2(n_1626),
.Y(n_2016)
);

OA21x2_ASAP7_75t_L g2017 ( 
.A1(n_1915),
.A2(n_1717),
.B(n_1714),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1873),
.B(n_1628),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1773),
.Y(n_2019)
);

BUFx4_ASAP7_75t_SL g2020 ( 
.A(n_1786),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1891),
.A2(n_1632),
.B(n_1552),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1847),
.Y(n_2022)
);

AOI21x1_ASAP7_75t_SL g2023 ( 
.A1(n_1848),
.A2(n_1829),
.B(n_1904),
.Y(n_2023)
);

O2A1O1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_1859),
.A2(n_1592),
.B(n_1647),
.C(n_1645),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_1798),
.Y(n_2025)
);

INVx5_ASAP7_75t_L g2026 ( 
.A(n_1837),
.Y(n_2026)
);

BUFx2_ASAP7_75t_L g2027 ( 
.A(n_1928),
.Y(n_2027)
);

CKINVDCx20_ASAP7_75t_R g2028 ( 
.A(n_1833),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_2001),
.A2(n_1554),
.B(n_1634),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1784),
.Y(n_2030)
);

AO22x2_ASAP7_75t_L g2031 ( 
.A1(n_1871),
.A2(n_1599),
.B1(n_1648),
.B2(n_1640),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1775),
.Y(n_2032)
);

AO31x2_ASAP7_75t_L g2033 ( 
.A1(n_1889),
.A2(n_423),
.A3(n_421),
.B(n_422),
.Y(n_2033)
);

A2O1A1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1797),
.A2(n_426),
.B(n_424),
.C(n_425),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1883),
.A2(n_1862),
.B1(n_1861),
.B2(n_1972),
.Y(n_2035)
);

OAI22x1_ASAP7_75t_L g2036 ( 
.A1(n_1814),
.A2(n_428),
.B1(n_425),
.B2(n_427),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1990),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_2037)
);

AND2x4_ASAP7_75t_L g2038 ( 
.A(n_1774),
.B(n_430),
.Y(n_2038)
);

CKINVDCx20_ASAP7_75t_R g2039 ( 
.A(n_1776),
.Y(n_2039)
);

AOI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2003),
.A2(n_432),
.B(n_433),
.Y(n_2040)
);

NOR2xp67_ASAP7_75t_L g2041 ( 
.A(n_1826),
.B(n_1836),
.Y(n_2041)
);

O2A1O1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_1912),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1935),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1871),
.B(n_437),
.Y(n_2044)
);

AOI21x1_ASAP7_75t_SL g2045 ( 
.A1(n_2008),
.A2(n_438),
.B(n_440),
.Y(n_2045)
);

NAND3xp33_ASAP7_75t_SL g2046 ( 
.A(n_1824),
.B(n_441),
.C(n_442),
.Y(n_2046)
);

AO32x2_ASAP7_75t_L g2047 ( 
.A1(n_1788),
.A2(n_444),
.A3(n_441),
.B1(n_443),
.B2(n_445),
.Y(n_2047)
);

AO21x2_ASAP7_75t_L g2048 ( 
.A1(n_1886),
.A2(n_441),
.B(n_443),
.Y(n_2048)
);

OAI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1936),
.A2(n_444),
.B(n_445),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_1817),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1881),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1777),
.A2(n_1851),
.B1(n_1789),
.B2(n_1809),
.Y(n_2052)
);

AO21x1_ASAP7_75t_L g2053 ( 
.A1(n_1995),
.A2(n_448),
.B(n_449),
.Y(n_2053)
);

BUFx12f_ASAP7_75t_L g2054 ( 
.A(n_1821),
.Y(n_2054)
);

AO31x2_ASAP7_75t_L g2055 ( 
.A1(n_1782),
.A2(n_451),
.A3(n_448),
.B(n_450),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1932),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1940),
.B(n_450),
.Y(n_2057)
);

AO21x1_ASAP7_75t_L g2058 ( 
.A1(n_1923),
.A2(n_453),
.B(n_454),
.Y(n_2058)
);

INVx2_ASAP7_75t_SL g2059 ( 
.A(n_1790),
.Y(n_2059)
);

AO31x2_ASAP7_75t_L g2060 ( 
.A1(n_1987),
.A2(n_458),
.A3(n_456),
.B(n_457),
.Y(n_2060)
);

AOI211x1_ASAP7_75t_L g2061 ( 
.A1(n_1772),
.A2(n_1843),
.B(n_1872),
.C(n_1868),
.Y(n_2061)
);

O2A1O1Ixp33_ASAP7_75t_L g2062 ( 
.A1(n_1901),
.A2(n_461),
.B(n_459),
.C(n_460),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1961),
.B(n_459),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1966),
.B(n_460),
.Y(n_2064)
);

INVx4_ASAP7_75t_L g2065 ( 
.A(n_1795),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1832),
.B(n_1835),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_1929),
.A2(n_463),
.B(n_465),
.C(n_478),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1907),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1823),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1931),
.A2(n_463),
.B(n_465),
.C(n_478),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1937),
.B(n_479),
.Y(n_2071)
);

AOI221x1_ASAP7_75t_L g2072 ( 
.A1(n_1838),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.C(n_483),
.Y(n_2072)
);

INVx4_ASAP7_75t_L g2073 ( 
.A(n_1909),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1905),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_1853),
.A2(n_484),
.B(n_485),
.Y(n_2075)
);

OAI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_1960),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_2076)
);

NOR2xp67_ASAP7_75t_L g2077 ( 
.A(n_1825),
.B(n_488),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_1984),
.A2(n_490),
.B(n_491),
.Y(n_2078)
);

AO21x1_ASAP7_75t_L g2079 ( 
.A1(n_1923),
.A2(n_492),
.B(n_493),
.Y(n_2079)
);

AOI21xp5_ASAP7_75t_SL g2080 ( 
.A1(n_1898),
.A2(n_492),
.B(n_494),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1934),
.B(n_496),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_SL g2082 ( 
.A1(n_1839),
.A2(n_496),
.B(n_497),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_1917),
.A2(n_498),
.B(n_499),
.Y(n_2083)
);

OAI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1938),
.A2(n_498),
.B(n_499),
.Y(n_2084)
);

INVx3_ASAP7_75t_SL g2085 ( 
.A(n_1856),
.Y(n_2085)
);

OAI21x1_ASAP7_75t_L g2086 ( 
.A1(n_1952),
.A2(n_500),
.B(n_501),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1927),
.A2(n_500),
.B(n_502),
.Y(n_2087)
);

AO22x2_ASAP7_75t_L g2088 ( 
.A1(n_1882),
.A2(n_2007),
.B1(n_1933),
.B2(n_1955),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1895),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_2089)
);

AO32x2_ASAP7_75t_L g2090 ( 
.A1(n_1947),
.A2(n_508),
.A3(n_506),
.B1(n_507),
.B2(n_509),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1910),
.B(n_507),
.Y(n_2091)
);

AOI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1939),
.A2(n_508),
.B(n_509),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1811),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_2093)
);

OAI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_1942),
.A2(n_512),
.B(n_513),
.Y(n_2094)
);

BUFx2_ASAP7_75t_SL g2095 ( 
.A(n_1855),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1822),
.A2(n_518),
.B1(n_515),
.B2(n_517),
.Y(n_2096)
);

NOR2xp67_ASAP7_75t_L g2097 ( 
.A(n_1835),
.B(n_515),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1914),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_1968),
.A2(n_518),
.B(n_519),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1899),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_1930),
.A2(n_2005),
.B(n_1989),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1946),
.Y(n_2102)
);

BUFx10_ASAP7_75t_L g2103 ( 
.A(n_1910),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1913),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1820),
.A2(n_1925),
.B(n_1926),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1957),
.Y(n_2106)
);

OAI21x1_ASAP7_75t_L g2107 ( 
.A1(n_1975),
.A2(n_524),
.B(n_525),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_1810),
.B(n_527),
.Y(n_2108)
);

AOI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1791),
.A2(n_529),
.B(n_530),
.Y(n_2109)
);

OAI21xp5_ASAP7_75t_SL g2110 ( 
.A1(n_1785),
.A2(n_533),
.B(n_534),
.Y(n_2110)
);

BUFx5_ASAP7_75t_L g2111 ( 
.A(n_1855),
.Y(n_2111)
);

OR2x6_ASAP7_75t_L g2112 ( 
.A(n_1965),
.B(n_535),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2000),
.B(n_1803),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_1846),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1962),
.B(n_536),
.Y(n_2115)
);

INVx5_ASAP7_75t_L g2116 ( 
.A(n_1855),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1967),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1801),
.Y(n_2118)
);

OAI21x1_ASAP7_75t_L g2119 ( 
.A1(n_1802),
.A2(n_537),
.B(n_538),
.Y(n_2119)
);

OAI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1948),
.A2(n_539),
.B(n_540),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_1944),
.A2(n_541),
.B(n_543),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_1857),
.B(n_545),
.Y(n_2122)
);

AOI221x1_ASAP7_75t_L g2123 ( 
.A1(n_1831),
.A2(n_547),
.B1(n_545),
.B2(n_546),
.C(n_548),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1900),
.Y(n_2124)
);

INVx5_ASAP7_75t_L g2125 ( 
.A(n_1957),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1921),
.A2(n_549),
.B(n_550),
.Y(n_2126)
);

AOI211x1_ASAP7_75t_L g2127 ( 
.A1(n_1896),
.A2(n_562),
.B(n_560),
.C(n_561),
.Y(n_2127)
);

OA21x2_ASAP7_75t_L g2128 ( 
.A1(n_1977),
.A2(n_560),
.B(n_561),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_L g2129 ( 
.A(n_1969),
.B(n_563),
.Y(n_2129)
);

AND2x6_ASAP7_75t_L g2130 ( 
.A(n_1955),
.B(n_564),
.Y(n_2130)
);

A2O1A1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_1877),
.A2(n_567),
.B(n_565),
.C(n_566),
.Y(n_2131)
);

OAI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1964),
.A2(n_565),
.B(n_566),
.Y(n_2132)
);

AOI21xp33_ASAP7_75t_L g2133 ( 
.A1(n_1918),
.A2(n_570),
.B(n_571),
.Y(n_2133)
);

AOI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_1945),
.A2(n_572),
.B(n_574),
.Y(n_2134)
);

OAI21x1_ASAP7_75t_L g2135 ( 
.A1(n_1983),
.A2(n_575),
.B(n_576),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1878),
.A2(n_580),
.B1(n_577),
.B2(n_579),
.Y(n_2136)
);

INVx1_ASAP7_75t_SL g2137 ( 
.A(n_2102),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_2035),
.A2(n_1920),
.B1(n_1815),
.B2(n_1884),
.Y(n_2138)
);

INVx2_ASAP7_75t_SL g2139 ( 
.A(n_2020),
.Y(n_2139)
);

BUFx2_ASAP7_75t_SL g2140 ( 
.A(n_2026),
.Y(n_2140)
);

OAI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_2026),
.A2(n_1849),
.B1(n_1903),
.B2(n_1994),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2030),
.Y(n_2142)
);

BUFx3_ASAP7_75t_L g2143 ( 
.A(n_2022),
.Y(n_2143)
);

CKINVDCx20_ASAP7_75t_R g2144 ( 
.A(n_2028),
.Y(n_2144)
);

INVx3_ASAP7_75t_SL g2145 ( 
.A(n_2012),
.Y(n_2145)
);

OAI22xp33_ASAP7_75t_SL g2146 ( 
.A1(n_2112),
.A2(n_1888),
.B1(n_1954),
.B2(n_1869),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2116),
.A2(n_1954),
.B1(n_1799),
.B2(n_1949),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2100),
.Y(n_2148)
);

BUFx8_ASAP7_75t_L g2149 ( 
.A(n_2054),
.Y(n_2149)
);

INVx5_ASAP7_75t_L g2150 ( 
.A(n_2125),
.Y(n_2150)
);

OAI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2056),
.A2(n_1864),
.B1(n_1906),
.B2(n_1958),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_2116),
.A2(n_1916),
.B1(n_1819),
.B2(n_1980),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_2069),
.Y(n_2153)
);

INVx4_ASAP7_75t_L g2154 ( 
.A(n_2012),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_2117),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_2009),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2124),
.Y(n_2157)
);

BUFx3_ASAP7_75t_L g2158 ( 
.A(n_2027),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2097),
.A2(n_1787),
.B1(n_1997),
.B2(n_1982),
.Y(n_2159)
);

CKINVDCx11_ASAP7_75t_R g2160 ( 
.A(n_2050),
.Y(n_2160)
);

INVx6_ASAP7_75t_L g2161 ( 
.A(n_2073),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2098),
.Y(n_2162)
);

INVx8_ASAP7_75t_L g2163 ( 
.A(n_2039),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_2110),
.A2(n_2004),
.B1(n_1996),
.B2(n_1963),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_SL g2165 ( 
.A1(n_2088),
.A2(n_1854),
.B1(n_1840),
.B2(n_2002),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2037),
.A2(n_1998),
.B1(n_1985),
.B2(n_1956),
.Y(n_2166)
);

BUFx3_ASAP7_75t_L g2167 ( 
.A(n_2085),
.Y(n_2167)
);

CKINVDCx11_ASAP7_75t_R g2168 ( 
.A(n_2065),
.Y(n_2168)
);

INVx6_ASAP7_75t_L g2169 ( 
.A(n_2103),
.Y(n_2169)
);

CKINVDCx11_ASAP7_75t_R g2170 ( 
.A(n_2025),
.Y(n_2170)
);

BUFx8_ASAP7_75t_SL g2171 ( 
.A(n_2019),
.Y(n_2171)
);

BUFx12f_ASAP7_75t_L g2172 ( 
.A(n_2068),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_2059),
.Y(n_2173)
);

BUFx12f_ASAP7_75t_L g2174 ( 
.A(n_2114),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_2066),
.Y(n_2175)
);

CKINVDCx11_ASAP7_75t_R g2176 ( 
.A(n_2038),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_2088),
.A2(n_1892),
.B1(n_1911),
.B2(n_1894),
.Y(n_2177)
);

INVx6_ASAP7_75t_L g2178 ( 
.A(n_2106),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_2106),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_SL g2180 ( 
.A1(n_2095),
.A2(n_1974),
.B1(n_1863),
.B2(n_1941),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_SL g2181 ( 
.A1(n_2130),
.A2(n_1922),
.B1(n_1943),
.B2(n_1986),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_SL g2182 ( 
.A1(n_2130),
.A2(n_1971),
.B1(n_1792),
.B2(n_1993),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2043),
.A2(n_1991),
.B1(n_1781),
.B2(n_1879),
.Y(n_2183)
);

OAI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2051),
.A2(n_1999),
.B1(n_1852),
.B2(n_1834),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2060),
.Y(n_2185)
);

OAI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2074),
.A2(n_1924),
.B1(n_1979),
.B2(n_1970),
.Y(n_2186)
);

NAND2x1p5_ASAP7_75t_L g2187 ( 
.A(n_2041),
.B(n_1874),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2060),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_2057),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_2032),
.Y(n_2190)
);

INVxp67_ASAP7_75t_L g2191 ( 
.A(n_2129),
.Y(n_2191)
);

OAI21xp5_ASAP7_75t_SL g2192 ( 
.A1(n_2046),
.A2(n_1908),
.B(n_1880),
.Y(n_2192)
);

NAND2x1p5_ASAP7_75t_L g2193 ( 
.A(n_2081),
.B(n_1874),
.Y(n_2193)
);

AOI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_2044),
.A2(n_1953),
.B1(n_1779),
.B2(n_1778),
.Y(n_2194)
);

OAI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2018),
.A2(n_1981),
.B1(n_1794),
.B2(n_1796),
.Y(n_2195)
);

INVx6_ASAP7_75t_L g2196 ( 
.A(n_2111),
.Y(n_2196)
);

CKINVDCx6p67_ASAP7_75t_R g2197 ( 
.A(n_2111),
.Y(n_2197)
);

CKINVDCx6p67_ASAP7_75t_R g2198 ( 
.A(n_2036),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2067),
.A2(n_1867),
.B1(n_1808),
.B2(n_1806),
.Y(n_2199)
);

AOI22xp33_ASAP7_75t_SL g2200 ( 
.A1(n_2052),
.A2(n_1971),
.B1(n_1919),
.B2(n_1973),
.Y(n_2200)
);

INVx6_ASAP7_75t_L g2201 ( 
.A(n_2010),
.Y(n_2201)
);

BUFx12f_ASAP7_75t_L g2202 ( 
.A(n_2010),
.Y(n_2202)
);

CKINVDCx11_ASAP7_75t_R g2203 ( 
.A(n_2089),
.Y(n_2203)
);

BUFx3_ASAP7_75t_L g2204 ( 
.A(n_2122),
.Y(n_2204)
);

BUFx8_ASAP7_75t_L g2205 ( 
.A(n_2047),
.Y(n_2205)
);

AOI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2014),
.A2(n_1860),
.B1(n_1866),
.B2(n_1865),
.Y(n_2206)
);

AOI22xp33_ASAP7_75t_SL g2207 ( 
.A1(n_2049),
.A2(n_1973),
.B1(n_1874),
.B2(n_1978),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_2031),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2061),
.A2(n_1804),
.B1(n_1830),
.B2(n_1828),
.Y(n_2209)
);

BUFx2_ASAP7_75t_L g2210 ( 
.A(n_2031),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_2013),
.A2(n_1870),
.B1(n_1885),
.B2(n_1875),
.Y(n_2211)
);

AOI22xp33_ASAP7_75t_L g2212 ( 
.A1(n_2011),
.A2(n_1890),
.B1(n_1897),
.B2(n_1893),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2118),
.A2(n_1959),
.B1(n_1807),
.B2(n_1845),
.Y(n_2213)
);

INVx1_ASAP7_75t_SL g2214 ( 
.A(n_2108),
.Y(n_2214)
);

OAI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_2084),
.A2(n_1800),
.B1(n_1805),
.B2(n_1793),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_SL g2216 ( 
.A(n_2023),
.Y(n_2216)
);

INVx6_ASAP7_75t_L g2217 ( 
.A(n_2015),
.Y(n_2217)
);

INVx4_ASAP7_75t_L g2218 ( 
.A(n_2128),
.Y(n_2218)
);

CKINVDCx6p67_ASAP7_75t_R g2219 ( 
.A(n_2091),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_2115),
.Y(n_2220)
);

INVx6_ASAP7_75t_L g2221 ( 
.A(n_2045),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2113),
.B(n_1812),
.Y(n_2222)
);

BUFx4f_ASAP7_75t_L g2223 ( 
.A(n_2017),
.Y(n_2223)
);

INVx4_ASAP7_75t_L g2224 ( 
.A(n_2048),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_2094),
.A2(n_1988),
.B1(n_1992),
.B2(n_1976),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2158),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_2197),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2185),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2181),
.B(n_2077),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2188),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_2196),
.Y(n_2231)
);

AOI21xp33_ASAP7_75t_SL g2232 ( 
.A1(n_2145),
.A2(n_2104),
.B(n_2120),
.Y(n_2232)
);

AOI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2223),
.A2(n_2105),
.B(n_2101),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2165),
.A2(n_2127),
.B1(n_2132),
.B2(n_2070),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2148),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2142),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2157),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2162),
.Y(n_2238)
);

BUFx3_ASAP7_75t_L g2239 ( 
.A(n_2156),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2196),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_2161),
.Y(n_2241)
);

OR2x6_ASAP7_75t_L g2242 ( 
.A(n_2154),
.B(n_2080),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_2153),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2217),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_2143),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2204),
.B(n_2047),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_2202),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_2208),
.B(n_2029),
.Y(n_2248)
);

CKINVDCx6p67_ASAP7_75t_R g2249 ( 
.A(n_2160),
.Y(n_2249)
);

OR2x6_ASAP7_75t_L g2250 ( 
.A(n_2140),
.B(n_2058),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_2201),
.Y(n_2251)
);

INVxp33_ASAP7_75t_L g2252 ( 
.A(n_2176),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2214),
.B(n_2033),
.Y(n_2253)
);

OAI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_2198),
.A2(n_2123),
.B1(n_2096),
.B2(n_2072),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2177),
.A2(n_2087),
.B(n_2083),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2175),
.B(n_2090),
.Y(n_2256)
);

HB1xp67_ASAP7_75t_SL g2257 ( 
.A(n_2149),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2155),
.B(n_2090),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2210),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2218),
.Y(n_2260)
);

INVx2_ASAP7_75t_SL g2261 ( 
.A(n_2150),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2224),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2179),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2221),
.Y(n_2264)
);

INVxp67_ASAP7_75t_L g2265 ( 
.A(n_2173),
.Y(n_2265)
);

AO21x2_ASAP7_75t_L g2266 ( 
.A1(n_2195),
.A2(n_2082),
.B(n_2079),
.Y(n_2266)
);

INVx1_ASAP7_75t_SL g2267 ( 
.A(n_2170),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2221),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2222),
.B(n_2063),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_2150),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2216),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2137),
.B(n_2064),
.Y(n_2272)
);

AO21x2_ASAP7_75t_L g2273 ( 
.A1(n_2215),
.A2(n_2092),
.B(n_2071),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2205),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_2187),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2190),
.Y(n_2276)
);

INVx4_ASAP7_75t_L g2277 ( 
.A(n_2241),
.Y(n_2277)
);

NAND3xp33_ASAP7_75t_L g2278 ( 
.A(n_2262),
.B(n_2191),
.C(n_2220),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2226),
.B(n_2167),
.Y(n_2279)
);

AOI221xp5_ASAP7_75t_L g2280 ( 
.A1(n_2234),
.A2(n_2138),
.B1(n_2141),
.B2(n_2151),
.C(n_2186),
.Y(n_2280)
);

INVx5_ASAP7_75t_L g2281 ( 
.A(n_2241),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2250),
.A2(n_2182),
.B1(n_2200),
.B2(n_2219),
.Y(n_2282)
);

INVx1_ASAP7_75t_SL g2283 ( 
.A(n_2239),
.Y(n_2283)
);

OA21x2_ASAP7_75t_L g2284 ( 
.A1(n_2260),
.A2(n_2099),
.B(n_2086),
.Y(n_2284)
);

CKINVDCx20_ASAP7_75t_R g2285 ( 
.A(n_2249),
.Y(n_2285)
);

OAI21xp5_ASAP7_75t_L g2286 ( 
.A1(n_2229),
.A2(n_2207),
.B(n_2180),
.Y(n_2286)
);

AOI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_2233),
.A2(n_2146),
.B(n_2147),
.Y(n_2287)
);

AND2x4_ASAP7_75t_SL g2288 ( 
.A(n_2243),
.B(n_2139),
.Y(n_2288)
);

BUFx8_ASAP7_75t_L g2289 ( 
.A(n_2257),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2254),
.A2(n_2109),
.B(n_2192),
.Y(n_2290)
);

AO32x2_ASAP7_75t_L g2291 ( 
.A1(n_2261),
.A2(n_2209),
.A3(n_2152),
.B1(n_2159),
.B2(n_2199),
.Y(n_2291)
);

OA21x2_ASAP7_75t_L g2292 ( 
.A1(n_2260),
.A2(n_2107),
.B(n_2135),
.Y(n_2292)
);

AOI221xp5_ASAP7_75t_L g2293 ( 
.A1(n_2232),
.A2(n_2184),
.B1(n_2183),
.B2(n_2164),
.C(n_2133),
.Y(n_2293)
);

BUFx4f_ASAP7_75t_SL g2294 ( 
.A(n_2245),
.Y(n_2294)
);

CKINVDCx11_ASAP7_75t_R g2295 ( 
.A(n_2267),
.Y(n_2295)
);

OAI22xp5_ASAP7_75t_SL g2296 ( 
.A1(n_2252),
.A2(n_2144),
.B1(n_2172),
.B2(n_2174),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2274),
.A2(n_2193),
.B1(n_2169),
.B2(n_2211),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2246),
.B(n_2055),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2269),
.A2(n_2203),
.B1(n_2166),
.B2(n_2093),
.Y(n_2299)
);

NOR2x1_ASAP7_75t_R g2300 ( 
.A(n_2247),
.B(n_2168),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2276),
.B(n_2178),
.Y(n_2301)
);

A2O1A1Ixp33_ASAP7_75t_L g2302 ( 
.A1(n_2227),
.A2(n_2042),
.B(n_2062),
.C(n_2163),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2266),
.A2(n_2136),
.B1(n_2212),
.B2(n_2213),
.Y(n_2303)
);

OR2x6_ASAP7_75t_L g2304 ( 
.A(n_2271),
.B(n_2016),
.Y(n_2304)
);

OAI21x1_ASAP7_75t_SL g2305 ( 
.A1(n_2271),
.A2(n_2053),
.B(n_2040),
.Y(n_2305)
);

AOI221xp5_ASAP7_75t_L g2306 ( 
.A1(n_2253),
.A2(n_2259),
.B1(n_2258),
.B2(n_2237),
.C(n_2238),
.Y(n_2306)
);

OAI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2255),
.A2(n_2034),
.B(n_2078),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2235),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2298),
.B(n_2306),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_2280),
.A2(n_2248),
.B1(n_2273),
.B2(n_2242),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2308),
.Y(n_2311)
);

AOI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_2293),
.A2(n_2242),
.B1(n_2256),
.B2(n_2264),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_2289),
.Y(n_2313)
);

INVx1_ASAP7_75t_SL g2314 ( 
.A(n_2283),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2282),
.A2(n_2299),
.B1(n_2287),
.B2(n_2304),
.Y(n_2315)
);

OAI221xp5_ASAP7_75t_SL g2316 ( 
.A1(n_2303),
.A2(n_2265),
.B1(n_2272),
.B2(n_2227),
.C(n_2270),
.Y(n_2316)
);

OAI21xp33_ASAP7_75t_L g2317 ( 
.A1(n_2290),
.A2(n_2268),
.B(n_2264),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2301),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2279),
.B(n_2251),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2278),
.Y(n_2320)
);

INVx11_ASAP7_75t_L g2321 ( 
.A(n_2294),
.Y(n_2321)
);

BUFx3_ASAP7_75t_L g2322 ( 
.A(n_2288),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_2277),
.Y(n_2323)
);

INVxp67_ASAP7_75t_SL g2324 ( 
.A(n_2284),
.Y(n_2324)
);

INVx1_ASAP7_75t_SL g2325 ( 
.A(n_2281),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2291),
.Y(n_2326)
);

OAI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_2315),
.A2(n_2286),
.B(n_2302),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2326),
.B(n_2236),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2316),
.A2(n_2297),
.B1(n_2285),
.B2(n_2244),
.Y(n_2329)
);

INVx4_ASAP7_75t_L g2330 ( 
.A(n_2321),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_R g2331 ( 
.A(n_2313),
.B(n_2295),
.Y(n_2331)
);

INVx4_ASAP7_75t_L g2332 ( 
.A(n_2322),
.Y(n_2332)
);

AOI221xp5_ASAP7_75t_L g2333 ( 
.A1(n_2315),
.A2(n_2307),
.B1(n_2305),
.B2(n_2296),
.C(n_2076),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2314),
.Y(n_2334)
);

OAI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2312),
.A2(n_2275),
.B1(n_2291),
.B2(n_2263),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_2323),
.Y(n_2336)
);

OAI221xp5_ASAP7_75t_L g2337 ( 
.A1(n_2310),
.A2(n_2206),
.B1(n_2225),
.B2(n_2189),
.C(n_2194),
.Y(n_2337)
);

OAI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_2316),
.A2(n_2240),
.B1(n_2231),
.B2(n_2292),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2320),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2309),
.B(n_2228),
.Y(n_2340)
);

INVx8_ASAP7_75t_L g2341 ( 
.A(n_2319),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2318),
.B(n_2230),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2311),
.Y(n_2343)
);

NOR3xp33_ASAP7_75t_L g2344 ( 
.A(n_2327),
.B(n_2333),
.C(n_2329),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2340),
.B(n_2309),
.Y(n_2345)
);

INVx1_ASAP7_75t_SL g2346 ( 
.A(n_2336),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2328),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2343),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2339),
.B(n_2317),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2334),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2350),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_2349),
.B(n_2332),
.Y(n_2352)
);

AOI222xp33_ASAP7_75t_L g2353 ( 
.A1(n_2345),
.A2(n_2300),
.B1(n_2335),
.B2(n_2330),
.C1(n_2317),
.C2(n_2338),
.Y(n_2353)
);

NOR2x1_ASAP7_75t_R g2354 ( 
.A(n_2344),
.B(n_2171),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2347),
.B(n_2342),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2348),
.Y(n_2356)
);

AOI211xp5_ASAP7_75t_L g2357 ( 
.A1(n_2344),
.A2(n_2337),
.B(n_2331),
.C(n_2325),
.Y(n_2357)
);

OAI31xp33_ASAP7_75t_SL g2358 ( 
.A1(n_2346),
.A2(n_2324),
.A3(n_2325),
.B(n_2341),
.Y(n_2358)
);

AND5x1_ASAP7_75t_L g2359 ( 
.A(n_2357),
.B(n_2358),
.C(n_2354),
.D(n_2353),
.E(n_2352),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2351),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2355),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2355),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2356),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2361),
.B(n_2075),
.Y(n_2364)
);

OAI221xp5_ASAP7_75t_L g2365 ( 
.A1(n_2359),
.A2(n_2131),
.B1(n_2006),
.B2(n_2021),
.C(n_1844),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2360),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2362),
.B(n_2126),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2363),
.B(n_2134),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2368),
.Y(n_2369)
);

OAI31xp33_ASAP7_75t_L g2370 ( 
.A1(n_2366),
.A2(n_2365),
.A3(n_2367),
.B(n_2364),
.Y(n_2370)
);

OAI322xp33_ASAP7_75t_L g2371 ( 
.A1(n_2369),
.A2(n_1950),
.A3(n_1951),
.B1(n_1902),
.B2(n_1818),
.C1(n_1816),
.C2(n_1813),
.Y(n_2371)
);

NAND4xp25_ASAP7_75t_L g2372 ( 
.A(n_2370),
.B(n_1780),
.C(n_2121),
.D(n_2024),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2372),
.Y(n_2373)
);

AOI211xp5_ASAP7_75t_L g2374 ( 
.A1(n_2373),
.A2(n_2371),
.B(n_2119),
.C(n_592),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2374),
.A2(n_1841),
.B1(n_1850),
.B2(n_1827),
.Y(n_2375)
);

NOR2x1_ASAP7_75t_L g2376 ( 
.A(n_2375),
.B(n_598),
.Y(n_2376)
);

OAI221xp5_ASAP7_75t_L g2377 ( 
.A1(n_2376),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.C(n_607),
.Y(n_2377)
);

O2A1O1Ixp33_ASAP7_75t_L g2378 ( 
.A1(n_2377),
.A2(n_611),
.B(n_609),
.C(n_610),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2378),
.Y(n_2379)
);

AOI22x1_ASAP7_75t_L g2380 ( 
.A1(n_2379),
.A2(n_613),
.B1(n_610),
.B2(n_612),
.Y(n_2380)
);

INVxp67_ASAP7_75t_SL g2381 ( 
.A(n_2380),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2381),
.B(n_615),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2382),
.B(n_616),
.Y(n_2383)
);

AO21x2_ASAP7_75t_L g2384 ( 
.A1(n_2383),
.A2(n_617),
.B(n_618),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2384),
.Y(n_2385)
);

OAI221xp5_ASAP7_75t_R g2386 ( 
.A1(n_2385),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.C(n_621),
.Y(n_2386)
);

AOI211xp5_ASAP7_75t_L g2387 ( 
.A1(n_2386),
.A2(n_621),
.B(n_619),
.C(n_620),
.Y(n_2387)
);


endmodule