module real_jpeg_16895_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

NAND2x1_ASAP7_75t_SL g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2x1_ASAP7_75t_SL g55 ( 
.A(n_2),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_71),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_2),
.B(n_74),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_2),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_2),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_5),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_6),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_6),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_6),
.B(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_7),
.Y(n_121)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_7),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_8),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_8),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_8),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_8),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_8),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_8),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_9),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_9),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_9),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_9),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_9),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_9),
.B(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_11),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_13),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_78),
.B(n_208),
.C(n_320),
.D(n_337),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_165),
.C(n_187),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_142),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_20),
.B(n_142),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_R g20 ( 
.A(n_21),
.B(n_66),
.C(n_107),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_21),
.B(n_66),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_42),
.C(n_53),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_23),
.A2(n_24),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_24),
.B(n_33),
.C(n_39),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_24),
.B(n_173),
.C(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_24),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_24),
.A2(n_223),
.B(n_224),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x4_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_36),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_25),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_30),
.Y(n_240)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_33),
.B(n_120),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_33),
.A2(n_115),
.B(n_122),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_33),
.A2(n_34),
.B1(n_50),
.B2(n_106),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_34),
.B(n_73),
.C(n_120),
.Y(n_235)
);

O2A1O1Ixp5_ASAP7_75t_L g260 ( 
.A1(n_34),
.A2(n_50),
.B(n_261),
.C(n_266),
.Y(n_260)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_36),
.Y(n_137)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_37),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_55),
.C(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_38),
.A2(n_39),
.B1(n_133),
.B2(n_221),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_39),
.A2(n_70),
.B(n_94),
.Y(n_93)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_70),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_45),
.C(n_50),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_43),
.B(n_235),
.C(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_43),
.A2(n_44),
.B1(n_236),
.B2(n_237),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_105),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_50),
.A2(n_106),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_50),
.B(n_73),
.C(n_150),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_51),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_55),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_54),
.B(n_59),
.C(n_63),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_54),
.A2(n_55),
.B1(n_75),
.B2(n_76),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_SL g337 ( 
.A(n_54),
.B(n_76),
.C(n_200),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_55),
.B(n_94),
.C(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_82),
.C(n_85),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_63),
.B(n_76),
.C(n_231),
.Y(n_311)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_91),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_68),
.B(n_79),
.C(n_91),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_73),
.C(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_98),
.B(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_98),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_73),
.A2(n_78),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_73),
.A2(n_78),
.B1(n_163),
.B2(n_164),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_80),
.C(n_88),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_75),
.A2(n_76),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

AOI22x1_ASAP7_75t_SL g244 ( 
.A1(n_75),
.A2(n_76),
.B1(n_136),
.B2(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_128),
.C(n_136),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_88),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_76),
.B(n_117),
.C(n_125),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_81),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_85),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_82),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_82),
.B(n_98),
.C(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_82),
.A2(n_98),
.B1(n_113),
.B2(n_126),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_115),
.B(n_122),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_85),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_85),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_85),
.B(n_116),
.Y(n_204)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_88),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_129),
.C(n_133),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_104),
.Y(n_91)
);

XOR2x1_ASAP7_75t_L g246 ( 
.A(n_92),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_96),
.B(n_104),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_97),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_98),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_100),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_100),
.A2(n_200),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_107),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_127),
.C(n_138),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_108),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.C(n_123),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_114),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_116),
.A2(n_117),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_120),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_119),
.A2(n_120),
.B1(n_204),
.B2(n_205),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_120),
.B(n_125),
.C(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_120),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_123),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_127),
.A2(n_138),
.B1(n_139),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_128),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_129),
.A2(n_133),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_133),
.Y(n_221)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_136),
.Y(n_245)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_145),
.C(n_156),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_156),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_154),
.C(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_161),
.C(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_166),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_186),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_167),
.B(n_186),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_185),
.C(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_179),
.B1(n_180),
.B2(n_184),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_207)
);

OAI211xp5_ASAP7_75t_L g320 ( 
.A1(n_187),
.A2(n_321),
.B(n_324),
.C(n_325),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_188),
.B(n_190),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_207),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_206),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_192),
.B(n_206),
.C(n_207),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_202),
.B2(n_203),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_195),
.Y(n_201)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_328)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_250),
.B(n_319),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_248),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_211),
.B(n_248),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.C(n_246),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_212),
.B(n_246),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_215),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_234),
.C(n_241),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_230),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_222),
.A2(n_223),
.B1(n_230),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_234),
.A2(n_242),
.B1(n_243),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI31xp33_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_296),
.A3(n_314),
.B(n_318),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_285),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_285),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_275),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_254),
.B(n_276),
.C(n_281),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_271),
.C(n_273),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.C(n_259),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_260),
.Y(n_313)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.C(n_292),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_295),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_312),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.C(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_317),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_317),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_336),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_334),
.Y(n_335)
);


endmodule