module fake_netlist_5_469_n_5363 (n_924, n_977, n_611, n_1126, n_1166, n_469, n_82, n_785, n_549, n_532, n_1161, n_1150, n_226, n_667, n_790, n_1055, n_111, n_880, n_544, n_1007, n_155, n_552, n_1198, n_1099, n_956, n_564, n_423, n_21, n_105, n_1021, n_4, n_551, n_688, n_800, n_671, n_819, n_1022, n_915, n_864, n_173, n_859, n_951, n_447, n_247, n_292, n_625, n_854, n_674, n_417, n_516, n_933, n_1152, n_497, n_606, n_275, n_26, n_877, n_2, n_755, n_1118, n_6, n_947, n_373, n_307, n_530, n_87, n_150, n_1107, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_191, n_1104, n_659, n_51, n_171, n_1182, n_579, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_709, n_317, n_1236, n_569, n_227, n_920, n_94, n_335, n_370, n_976, n_343, n_308, n_297, n_156, n_1078, n_775, n_219, n_157, n_600, n_223, n_264, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_436, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1030, n_72, n_415, n_1071, n_485, n_1165, n_496, n_958, n_1034, n_670, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_680, n_395, n_164, n_553, n_901, n_813, n_214, n_675, n_888, n_1167, n_637, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_468, n_213, n_129, n_342, n_464, n_363, n_197, n_1069, n_1075, n_460, n_889, n_973, n_477, n_571, n_461, n_1211, n_1197, n_907, n_190, n_989, n_1039, n_34, n_228, n_283, n_488, n_736, n_892, n_1000, n_1202, n_1002, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_440, n_793, n_478, n_476, n_534, n_884, n_345, n_944, n_91, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_596, n_558, n_702, n_822, n_728, n_266, n_1162, n_272, n_1199, n_352, n_53, n_1038, n_520, n_409, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_434, n_868, n_639, n_914, n_411, n_414, n_965, n_935, n_121, n_1175, n_817, n_360, n_36, n_64, n_759, n_28, n_806, n_324, n_187, n_1189, n_103, n_97, n_11, n_7, n_706, n_746, n_747, n_52, n_784, n_110, n_1244, n_431, n_1194, n_615, n_851, n_843, n_523, n_913, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_776, n_367, n_452, n_525, n_649, n_547, n_43, n_1191, n_116, n_284, n_1128, n_139, n_744, n_590, n_629, n_254, n_1233, n_23, n_526, n_293, n_372, n_677, n_244, n_47, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1008, n_946, n_1001, n_498, n_689, n_738, n_640, n_252, n_624, n_295, n_133, n_1010, n_1231, n_739, n_1195, n_610, n_936, n_568, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1158, n_563, n_1145, n_878, n_524, n_204, n_394, n_1049, n_1153, n_741, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_658, n_456, n_959, n_535, n_152, n_940, n_9, n_592, n_1169, n_45, n_1017, n_123, n_978, n_1054, n_1095, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_484, n_1033, n_442, n_131, n_636, n_660, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_374, n_185, n_396, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_723, n_1065, n_473, n_1043, n_355, n_486, n_614, n_337, n_88, n_1177, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_361, n_700, n_1237, n_573, n_69, n_1132, n_388, n_1127, n_761, n_1006, n_329, n_274, n_582, n_73, n_19, n_309, n_30, n_512, n_84, n_130, n_322, n_1249, n_652, n_1111, n_25, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_44, n_224, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_987, n_261, n_174, n_767, n_993, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_83, n_513, n_1094, n_560, n_340, n_1044, n_1205, n_346, n_1209, n_495, n_602, n_574, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_490, n_996, n_921, n_233, n_572, n_366, n_815, n_128, n_120, n_327, n_135, n_1037, n_1080, n_426, n_1082, n_589, n_716, n_562, n_62, n_952, n_1229, n_391, n_701, n_1023, n_645, n_539, n_803, n_1092, n_238, n_531, n_890, n_764, n_1056, n_162, n_960, n_222, n_1123, n_1047, n_634, n_199, n_32, n_348, n_1029, n_925, n_1206, n_424, n_256, n_950, n_380, n_419, n_444, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_376, n_967, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_483, n_683, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_983, n_38, n_280, n_873, n_378, n_1112, n_762, n_17, n_690, n_33, n_583, n_302, n_1203, n_821, n_321, n_1179, n_621, n_753, n_455, n_1048, n_212, n_385, n_507, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1185, n_991, n_828, n_779, n_576, n_1143, n_804, n_537, n_945, n_492, n_153, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_883, n_470, n_325, n_449, n_132, n_1214, n_900, n_856, n_918, n_942, n_189, n_1147, n_13, n_1077, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_831, n_964, n_1096, n_234, n_833, n_5, n_225, n_988, n_814, n_192, n_1201, n_1114, n_655, n_669, n_472, n_1176, n_387, n_1149, n_398, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_50, n_430, n_510, n_216, n_311, n_830, n_801, n_241, n_875, n_357, n_1110, n_445, n_749, n_1134, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_734, n_638, n_866, n_107, n_969, n_1019, n_1105, n_249, n_304, n_577, n_338, n_149, n_693, n_14, n_836, n_990, n_975, n_567, n_778, n_1122, n_151, n_306, n_458, n_770, n_1102, n_711, n_85, n_1187, n_1164, n_489, n_1174, n_617, n_876, n_1190, n_118, n_601, n_917, n_966, n_253, n_1116, n_1212, n_172, n_206, n_217, n_726, n_982, n_818, n_861, n_1183, n_899, n_210, n_774, n_1059, n_176, n_1133, n_557, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_393, n_108, n_487, n_665, n_66, n_177, n_421, n_910, n_768, n_205, n_1136, n_754, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_202, n_427, n_791, n_732, n_193, n_808, n_797, n_1025, n_500, n_1067, n_148, n_435, n_159, n_766, n_541, n_538, n_1117, n_799, n_687, n_715, n_1213, n_536, n_872, n_594, n_200, n_1155, n_89, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_626, n_1144, n_1137, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_194, n_855, n_1178, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_605, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_780, n_998, n_467, n_1227, n_840, n_501, n_823, n_245, n_725, n_672, n_581, n_382, n_554, n_898, n_1013, n_718, n_265, n_1120, n_719, n_443, n_198, n_714, n_909, n_997, n_932, n_612, n_788, n_119, n_559, n_825, n_508, n_506, n_737, n_986, n_509, n_147, n_67, n_1192, n_1024, n_1063, n_209, n_733, n_941, n_981, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_282, n_752, n_905, n_1108, n_782, n_1100, n_862, n_760, n_381, n_220, n_390, n_31, n_481, n_769, n_42, n_1046, n_271, n_934, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_570, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_138, n_961, n_771, n_276, n_95, n_1225, n_169, n_522, n_400, n_930, n_181, n_221, n_622, n_1087, n_386, n_994, n_848, n_1223, n_104, n_682, n_56, n_141, n_1247, n_922, n_816, n_591, n_145, n_313, n_631, n_479, n_1246, n_432, n_839, n_1210, n_328, n_140, n_369, n_871, n_598, n_685, n_928, n_608, n_78, n_772, n_499, n_517, n_98, n_402, n_413, n_1086, n_796, n_236, n_1012, n_1, n_903, n_740, n_203, n_384, n_80, n_35, n_277, n_1061, n_92, n_333, n_462, n_1193, n_258, n_1113, n_29, n_79, n_1226, n_722, n_188, n_844, n_201, n_471, n_852, n_40, n_1028, n_781, n_474, n_542, n_463, n_595, n_502, n_466, n_420, n_632, n_699, n_979, n_1245, n_846, n_465, n_76, n_362, n_170, n_27, n_161, n_273, n_585, n_270, n_616, n_81, n_745, n_1103, n_648, n_312, n_1076, n_1091, n_494, n_641, n_730, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1220, n_37, n_229, n_437, n_60, n_403, n_453, n_1130, n_720, n_0, n_863, n_805, n_113, n_712, n_246, n_1042, n_269, n_285, n_412, n_657, n_644, n_1160, n_491, n_1074, n_251, n_160, n_566, n_565, n_597, n_1181, n_1196, n_651, n_334, n_811, n_807, n_835, n_175, n_666, n_262, n_99, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1018, n_438, n_713, n_904, n_166, n_1180, n_533, n_278, n_5363);

input n_924;
input n_977;
input n_611;
input n_1126;
input n_1166;
input n_469;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1150;
input n_226;
input n_667;
input n_790;
input n_1055;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1198;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_688;
input n_800;
input n_671;
input n_819;
input n_1022;
input n_915;
input n_864;
input n_173;
input n_859;
input n_951;
input n_447;
input n_247;
input n_292;
input n_625;
input n_854;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_755;
input n_1118;
input n_6;
input n_947;
input n_373;
input n_307;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_191;
input n_1104;
input n_659;
input n_51;
input n_171;
input n_1182;
input n_579;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_709;
input n_317;
input n_1236;
input n_569;
input n_227;
input n_920;
input n_94;
input n_335;
input n_370;
input n_976;
input n_343;
input n_308;
input n_297;
input n_156;
input n_1078;
input n_775;
input n_219;
input n_157;
input n_600;
input n_223;
input n_264;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_436;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1030;
input n_72;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_496;
input n_958;
input n_1034;
input n_670;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_680;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_214;
input n_675;
input n_888;
input n_1167;
input n_637;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_197;
input n_1069;
input n_1075;
input n_460;
input n_889;
input n_973;
input n_477;
input n_571;
input n_461;
input n_1211;
input n_1197;
input n_907;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1002;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_440;
input n_793;
input n_478;
input n_476;
input n_534;
input n_884;
input n_345;
input n_944;
input n_91;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_596;
input n_558;
input n_702;
input n_822;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1199;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_409;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_434;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_965;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_64;
input n_759;
input n_28;
input n_806;
input n_324;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_706;
input n_746;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_843;
input n_523;
input n_913;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_776;
input n_367;
input n_452;
input n_525;
input n_649;
input n_547;
input n_43;
input n_1191;
input n_116;
input n_284;
input n_1128;
input n_139;
input n_744;
input n_590;
input n_629;
input n_254;
input n_1233;
input n_23;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1008;
input n_946;
input n_1001;
input n_498;
input n_689;
input n_738;
input n_640;
input n_252;
input n_624;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1195;
input n_610;
input n_936;
input n_568;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1158;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1049;
input n_1153;
input n_741;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_658;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_9;
input n_592;
input n_1169;
input n_45;
input n_1017;
input n_123;
input n_978;
input n_1054;
input n_1095;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_484;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_374;
input n_185;
input n_396;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_723;
input n_1065;
input n_473;
input n_1043;
input n_355;
input n_486;
input n_614;
input n_337;
input n_88;
input n_1177;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1132;
input n_388;
input n_1127;
input n_761;
input n_1006;
input n_329;
input n_274;
input n_582;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_84;
input n_130;
input n_322;
input n_1249;
input n_652;
input n_1111;
input n_25;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_44;
input n_224;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_987;
input n_261;
input n_174;
input n_767;
input n_993;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_83;
input n_513;
input n_1094;
input n_560;
input n_340;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_495;
input n_602;
input n_574;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_490;
input n_996;
input n_921;
input n_233;
input n_572;
input n_366;
input n_815;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1037;
input n_1080;
input n_426;
input n_1082;
input n_589;
input n_716;
input n_562;
input n_62;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_531;
input n_890;
input n_764;
input n_1056;
input n_162;
input n_960;
input n_222;
input n_1123;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_348;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_256;
input n_950;
input n_380;
input n_419;
input n_444;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_376;
input n_967;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_483;
input n_683;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_983;
input n_38;
input n_280;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1203;
input n_821;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_212;
input n_385;
input n_507;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_804;
input n_537;
input n_945;
input n_492;
input n_153;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_883;
input n_470;
input n_325;
input n_449;
input n_132;
input n_1214;
input n_900;
input n_856;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_13;
input n_1077;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_831;
input n_964;
input n_1096;
input n_234;
input n_833;
input n_5;
input n_225;
input n_988;
input n_814;
input n_192;
input n_1201;
input n_1114;
input n_655;
input n_669;
input n_472;
input n_1176;
input n_387;
input n_1149;
input n_398;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_445;
input n_749;
input n_1134;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_577;
input n_338;
input n_149;
input n_693;
input n_14;
input n_836;
input n_990;
input n_975;
input n_567;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1102;
input n_711;
input n_85;
input n_1187;
input n_1164;
input n_489;
input n_1174;
input n_617;
input n_876;
input n_1190;
input n_118;
input n_601;
input n_917;
input n_966;
input n_253;
input n_1116;
input n_1212;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_818;
input n_861;
input n_1183;
input n_899;
input n_210;
input n_774;
input n_1059;
input n_176;
input n_1133;
input n_557;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_393;
input n_108;
input n_487;
input n_665;
input n_66;
input n_177;
input n_421;
input n_910;
input n_768;
input n_205;
input n_1136;
input n_754;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_202;
input n_427;
input n_791;
input n_732;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_148;
input n_435;
input n_159;
input n_766;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1213;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1155;
input n_89;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_626;
input n_1144;
input n_1137;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_194;
input n_855;
input n_1178;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_605;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_780;
input n_998;
input n_467;
input n_1227;
input n_840;
input n_501;
input n_823;
input n_245;
input n_725;
input n_672;
input n_581;
input n_382;
input n_554;
input n_898;
input n_1013;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_198;
input n_714;
input n_909;
input n_997;
input n_932;
input n_612;
input n_788;
input n_119;
input n_559;
input n_825;
input n_508;
input n_506;
input n_737;
input n_986;
input n_509;
input n_147;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_733;
input n_941;
input n_981;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_282;
input n_752;
input n_905;
input n_1108;
input n_782;
input n_1100;
input n_862;
input n_760;
input n_381;
input n_220;
input n_390;
input n_31;
input n_481;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_570;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_138;
input n_961;
input n_771;
input n_276;
input n_95;
input n_1225;
input n_169;
input n_522;
input n_400;
input n_930;
input n_181;
input n_221;
input n_622;
input n_1087;
input n_386;
input n_994;
input n_848;
input n_1223;
input n_104;
input n_682;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_591;
input n_145;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_432;
input n_839;
input n_1210;
input n_328;
input n_140;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_78;
input n_772;
input n_499;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_236;
input n_1012;
input n_1;
input n_903;
input n_740;
input n_203;
input n_384;
input n_80;
input n_35;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_462;
input n_1193;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_40;
input n_1028;
input n_781;
input n_474;
input n_542;
input n_463;
input n_595;
input n_502;
input n_466;
input n_420;
input n_632;
input n_699;
input n_979;
input n_1245;
input n_846;
input n_465;
input n_76;
input n_362;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1103;
input n_648;
input n_312;
input n_1076;
input n_1091;
input n_494;
input n_641;
input n_730;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1220;
input n_37;
input n_229;
input n_437;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_863;
input n_805;
input n_113;
input n_712;
input n_246;
input n_1042;
input n_269;
input n_285;
input n_412;
input n_657;
input n_644;
input n_1160;
input n_491;
input n_1074;
input n_251;
input n_160;
input n_566;
input n_565;
input n_597;
input n_1181;
input n_1196;
input n_651;
input n_334;
input n_811;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_99;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1018;
input n_438;
input n_713;
input n_904;
input n_166;
input n_1180;
input n_533;
input n_278;

output n_5363;

wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_2487;
wire n_1695;
wire n_1466;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_1696;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_2091;
wire n_1517;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_4255;
wire n_1796;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_3983;
wire n_4405;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_1385;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_4786;
wire n_3257;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_3790;
wire n_3491;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_4391;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_4918;
wire n_3856;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4232;
wire n_4125;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_5210;
wire n_4967;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_3200;
wire n_1664;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_3468;
wire n_2910;
wire n_1893;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_4443;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_4452;
wire n_4348;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_3073;
wire n_4572;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_3040;
wire n_1938;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_5322;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_4761;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_2559;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_1657;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1491;
wire n_3639;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_2754;
wire n_1742;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1418;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_3628;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_2774;
wire n_1707;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_2476;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_3738;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_3521;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_2920;
wire n_4265;
wire n_5319;
wire n_2247;
wire n_1622;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_5088;
wire n_2302;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_5352;
wire n_4991;
wire n_1698;
wire n_2329;
wire n_2142;
wire n_3332;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_2985;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_3367;
wire n_4464;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_2356;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_4353;
wire n_2042;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_3667;
wire n_1987;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_1609;
wire n_5298;
wire n_1887;
wire n_4413;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_2255;
wire n_2272;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_2878;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_2656;
wire n_1274;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_1919;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_1283;
wire n_5325;
wire n_2637;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_3282;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_5173;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_4467;
wire n_2377;
wire n_2080;
wire n_2340;
wire n_3552;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1603;
wire n_1401;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_5243;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1318;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_2221;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_3862;
wire n_5214;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1772;
wire n_1476;
wire n_2818;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_3289;
wire n_1973;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_3497;
wire n_1601;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1505;
wire n_4012;
wire n_4636;
wire n_4584;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_2599;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1751;
wire n_1508;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_3766;
wire n_1353;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_1686;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_4144;
wire n_2165;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_5131;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_1294;
wire n_1257;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_5280;
wire n_1428;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_5206;
wire n_3222;
wire n_1267;
wire n_1801;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_2636;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_5139;
wire n_2319;
wire n_1393;
wire n_3481;
wire n_2808;
wire n_2676;
wire n_2679;
wire n_1709;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_4627;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_1639;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_2116;
wire n_1434;
wire n_1828;
wire n_2320;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5216;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_2595;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_3065;
wire n_4361;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_1630;
wire n_4891;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_3800;
wire n_2403;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2685;
wire n_2037;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_3078;
wire n_3253;
wire n_4027;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_5359;
wire n_2574;
wire n_5293;
wire n_1358;
wire n_4316;
wire n_3697;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5200;
wire n_1653;
wire n_1506;
wire n_2867;
wire n_1894;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_3902;
wire n_4730;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_2224;
wire n_1991;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_4853;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5077;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_5314;
wire n_1618;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_3512;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_2004;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_5217;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_2374;
wire n_1545;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_3186;
wire n_4955;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_2936;
wire n_1946;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_2249;
wire n_2180;
wire n_4135;
wire n_2632;
wire n_1547;
wire n_1755;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1986;
wire n_1471;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_5288;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_3296;
wire n_1775;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_2491;
wire n_1788;
wire n_5079;
wire n_3833;
wire n_1679;
wire n_4841;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_3471;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_3031;
wire n_3701;
wire n_3243;
wire n_1773;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1920;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_5054;
wire n_2467;
wire n_2288;
wire n_4063;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_4541;
wire n_3824;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_2534;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_1424;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1432;
wire n_3875;
wire n_4003;
wire n_5299;
wire n_2402;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1342;
wire n_1400;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_3342;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_3123;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_2217;
wire n_1453;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_2722;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_3432;
wire n_1628;
wire n_1514;
wire n_1771;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_1533;
wire n_5036;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_1782;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_2819;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_1641;
wire n_3184;
wire n_1361;
wire n_4828;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_3302;
wire n_5304;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_1627;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_5270;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4364;
wire n_4245;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_398),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_483),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_764),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1037),
.Y(n_1253)
);

BUFx10_ASAP7_75t_L g1254 ( 
.A(n_1035),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_21),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_868),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_463),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_317),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_433),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_869),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_38),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_99),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1031),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1238),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_412),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_854),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_1216),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1219),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1189),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_137),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_168),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_856),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_715),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_832),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_372),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_64),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_967),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_660),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1149),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1121),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_512),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1071),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_595),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1241),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_282),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1117),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_78),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_623),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1173),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_962),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_528),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_96),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_115),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_438),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_185),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1214),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_587),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_463),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1188),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_900),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_273),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1199),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_175),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_810),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_220),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_603),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_717),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_974),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_283),
.Y(n_1309)
);

INVxp33_ASAP7_75t_R g1310 ( 
.A(n_965),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_886),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_239),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1179),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_495),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_605),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1033),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1056),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_873),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1007),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_842),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_67),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1096),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_336),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_977),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_966),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1050),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1014),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_936),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_586),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_801),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_606),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1212),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_81),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_410),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_898),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1060),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1068),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_74),
.Y(n_1338)
);

CKINVDCx14_ASAP7_75t_R g1339 ( 
.A(n_1063),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_503),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1038),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_846),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_163),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_722),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1052),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_105),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1169),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_547),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1207),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1013),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1165),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_500),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_553),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_995),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_901),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1167),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_300),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_120),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_177),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1186),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_523),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_561),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1147),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_777),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_937),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_381),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_562),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_944),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_763),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_971),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1196),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_251),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_246),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_774),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_998),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1176),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_993),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_53),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_536),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_879),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_526),
.Y(n_1381)
);

BUFx5_ASAP7_75t_L g1382 ( 
.A(n_1204),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_275),
.Y(n_1383)
);

BUFx8_ASAP7_75t_SL g1384 ( 
.A(n_1203),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_606),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_981),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_763),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_281),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_685),
.Y(n_1389)
);

BUFx2_ASAP7_75t_SL g1390 ( 
.A(n_810),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1092),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_732),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_184),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_636),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_359),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_216),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_773),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_501),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1134),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1078),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1002),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_660),
.Y(n_1402)
);

BUFx10_ASAP7_75t_L g1403 ( 
.A(n_848),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1064),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_384),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1104),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1233),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_172),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_426),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_859),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_610),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_838),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_330),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_912),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1054),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1218),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_354),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_343),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1242),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1157),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_916),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_855),
.Y(n_1422)
);

CKINVDCx14_ASAP7_75t_R g1423 ( 
.A(n_994),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_473),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_157),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_841),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_843),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_194),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1069),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_371),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_985),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1243),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_372),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1089),
.Y(n_1434)
);

CKINVDCx14_ASAP7_75t_R g1435 ( 
.A(n_314),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1055),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1075),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_281),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_978),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_879),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1070),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_6),
.Y(n_1442)
);

CKINVDCx14_ASAP7_75t_R g1443 ( 
.A(n_395),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_742),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_637),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_301),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_702),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1059),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_989),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_206),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_663),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_818),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1142),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_14),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_976),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1213),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_1040),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_975),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1051),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1036),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1011),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_373),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1128),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_543),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_496),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_297),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1192),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_632),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1151),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_247),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_72),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_590),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1086),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_705),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1113),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1115),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_585),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1197),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_555),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1138),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_6),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_457),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_525),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1123),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_212),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_699),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_268),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_327),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1124),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_66),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_988),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_417),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1003),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_716),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_884),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_679),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1082),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_832),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_528),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_844),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_99),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1107),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_577),
.Y(n_1503)
);

INVxp33_ASAP7_75t_L g1504 ( 
.A(n_809),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1166),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_572),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_299),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_550),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1202),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1174),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_964),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1211),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_567),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_153),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1023),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_827),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_13),
.Y(n_1517)
);

BUFx10_ASAP7_75t_L g1518 ( 
.A(n_1109),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_592),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_717),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_373),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1032),
.Y(n_1522)
);

CKINVDCx16_ASAP7_75t_R g1523 ( 
.A(n_1131),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_152),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1125),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_231),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1232),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1222),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1248),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_336),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_744),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_100),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_778),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_66),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_254),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_52),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_394),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1146),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_94),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_972),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1249),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_248),
.Y(n_1542)
);

BUFx5_ASAP7_75t_L g1543 ( 
.A(n_1079),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_288),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_771),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1135),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1021),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_474),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_924),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_991),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_878),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1224),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1100),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_663),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_22),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_919),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1098),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_865),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_612),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1127),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_431),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1010),
.Y(n_1562)
);

BUFx10_ASAP7_75t_L g1563 ( 
.A(n_1163),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_711),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_850),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_270),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_440),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_283),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_842),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1229),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_42),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_376),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_601),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_316),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_857),
.Y(n_1575)
);

BUFx10_ASAP7_75t_L g1576 ( 
.A(n_1220),
.Y(n_1576)
);

BUFx8_ASAP7_75t_SL g1577 ( 
.A(n_1112),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1029),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_656),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1017),
.Y(n_1580)
);

BUFx2_ASAP7_75t_SL g1581 ( 
.A(n_19),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_982),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_706),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_106),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_757),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1244),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_134),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1234),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1225),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_997),
.Y(n_1590)
);

BUFx5_ASAP7_75t_L g1591 ( 
.A(n_1012),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_184),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_577),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_356),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_624),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_597),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_561),
.Y(n_1597)
);

BUFx10_ASAP7_75t_L g1598 ( 
.A(n_860),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1236),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1177),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1094),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_54),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_276),
.Y(n_1603)
);

BUFx5_ASAP7_75t_L g1604 ( 
.A(n_1015),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_345),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_2),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_468),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_305),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_270),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1108),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_23),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_191),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_775),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_347),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1006),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1136),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1097),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_636),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_156),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_366),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1140),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_550),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1155),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1226),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1119),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_272),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_354),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_885),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_858),
.Y(n_1629)
);

CKINVDCx20_ASAP7_75t_R g1630 ( 
.A(n_301),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1105),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_331),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_121),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1102),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_709),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1210),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_761),
.Y(n_1637)
);

CKINVDCx20_ASAP7_75t_R g1638 ( 
.A(n_443),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1145),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_395),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_167),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_40),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1178),
.Y(n_1643)
);

CKINVDCx16_ASAP7_75t_R g1644 ( 
.A(n_1084),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_958),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_353),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_881),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_806),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_62),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_882),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_877),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1215),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1076),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_488),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1182),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_130),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1065),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1041),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1072),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_874),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1201),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_148),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1053),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1066),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1058),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_286),
.Y(n_1666)
);

BUFx10_ASAP7_75t_L g1667 ( 
.A(n_665),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1221),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1194),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_358),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1008),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1049),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1150),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_189),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_399),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_620),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_198),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1237),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_267),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_125),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_757),
.Y(n_1681)
);

BUFx3_ASAP7_75t_L g1682 ( 
.A(n_1095),
.Y(n_1682)
);

BUFx2_ASAP7_75t_SL g1683 ( 
.A(n_317),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_635),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_980),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_24),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_249),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1085),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1239),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1016),
.Y(n_1690)
);

BUFx5_ASAP7_75t_L g1691 ( 
.A(n_1110),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1114),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_74),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1045),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_287),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_595),
.Y(n_1696)
);

CKINVDCx16_ASAP7_75t_R g1697 ( 
.A(n_837),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1130),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_461),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_492),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_947),
.Y(n_1701)
);

BUFx5_ASAP7_75t_L g1702 ( 
.A(n_210),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_863),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_585),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_862),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_159),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_983),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_527),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_335),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_81),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_546),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_953),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_807),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_712),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_968),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_552),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_458),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_455),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_152),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_197),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1081),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1062),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_445),
.Y(n_1723)
);

BUFx8_ASAP7_75t_SL g1724 ( 
.A(n_1180),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_48),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_754),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_206),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_458),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_394),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_176),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1004),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_938),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_287),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_536),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_452),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_10),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1022),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_870),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_588),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_228),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_883),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1172),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_751),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_630),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1209),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_428),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_769),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_266),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_75),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_867),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1245),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_973),
.Y(n_1752)
);

CKINVDCx20_ASAP7_75t_R g1753 ( 
.A(n_1067),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1025),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_728),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_47),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1120),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_665),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1206),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_791),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_387),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_880),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_63),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_591),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_740),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1183),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_166),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_652),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1090),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_514),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_436),
.Y(n_1771)
);

CKINVDCx20_ASAP7_75t_R g1772 ( 
.A(n_22),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_941),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1164),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_713),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1009),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_388),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1103),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1132),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_227),
.Y(n_1780)
);

CKINVDCx16_ASAP7_75t_R g1781 ( 
.A(n_451),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_278),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_494),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_845),
.Y(n_1784)
);

CKINVDCx16_ASAP7_75t_R g1785 ( 
.A(n_511),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1005),
.Y(n_1786)
);

BUFx5_ASAP7_75t_L g1787 ( 
.A(n_19),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_850),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1205),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_950),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_956),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_149),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1087),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1133),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_51),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_502),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_44),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1122),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_89),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_376),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_404),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1061),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_387),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_866),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_504),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1227),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_314),
.Y(n_1807)
);

CKINVDCx20_ASAP7_75t_R g1808 ( 
.A(n_1018),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_67),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_330),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1000),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1019),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1191),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_805),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_745),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_92),
.Y(n_1816)
);

CKINVDCx20_ASAP7_75t_R g1817 ( 
.A(n_860),
.Y(n_1817)
);

BUFx10_ASAP7_75t_L g1818 ( 
.A(n_1046),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1026),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1047),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_84),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_344),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1200),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_680),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_801),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_876),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_784),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1168),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_462),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_869),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_4),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_910),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1223),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_824),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_279),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_714),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1116),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1217),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1057),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_746),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_659),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_343),
.Y(n_1842)
);

CKINVDCx20_ASAP7_75t_R g1843 ( 
.A(n_535),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1137),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_260),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_230),
.Y(n_1846)
);

CKINVDCx20_ASAP7_75t_R g1847 ( 
.A(n_149),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_979),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1187),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_1158),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1093),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_792),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_872),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1106),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_35),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1048),
.Y(n_1856)
);

CKINVDCx16_ASAP7_75t_R g1857 ( 
.A(n_1083),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_875),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1143),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_72),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_843),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_491),
.Y(n_1862)
);

INVxp67_ASAP7_75t_L g1863 ( 
.A(n_1088),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_174),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_727),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_504),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_157),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_634),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_861),
.Y(n_1869)
);

CKINVDCx20_ASAP7_75t_R g1870 ( 
.A(n_526),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_83),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_486),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1141),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1193),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_388),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1034),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_586),
.Y(n_1877)
);

INVx2_ASAP7_75t_SL g1878 ( 
.A(n_1231),
.Y(n_1878)
);

CKINVDCx20_ASAP7_75t_R g1879 ( 
.A(n_720),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_24),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_246),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_304),
.Y(n_1882)
);

BUFx10_ASAP7_75t_L g1883 ( 
.A(n_309),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_854),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_138),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_568),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1181),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_426),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_686),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_195),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_419),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_476),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_538),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_542),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1171),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_811),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1126),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_654),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_624),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_396),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1118),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_587),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1099),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1091),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_864),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_852),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_970),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1161),
.Y(n_1908)
);

BUFx10_ASAP7_75t_L g1909 ( 
.A(n_516),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_562),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1039),
.Y(n_1911)
);

BUFx10_ASAP7_75t_L g1912 ( 
.A(n_547),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1240),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1160),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_28),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_450),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_999),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_73),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1162),
.Y(n_1919)
);

CKINVDCx16_ASAP7_75t_R g1920 ( 
.A(n_987),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1190),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_996),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_166),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_868),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1154),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_627),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_961),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1230),
.Y(n_1928)
);

BUFx10_ASAP7_75t_L g1929 ( 
.A(n_524),
.Y(n_1929)
);

CKINVDCx20_ASAP7_75t_R g1930 ( 
.A(n_599),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_344),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1077),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1208),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1246),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_323),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_887),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_847),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_849),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_545),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_473),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_396),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_744),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_516),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_113),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_796),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_969),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_851),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_497),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_44),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_990),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_39),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_136),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_79),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_805),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1073),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_69),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1156),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1027),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_713),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_838),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_743),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_714),
.Y(n_1962)
);

BUFx10_ASAP7_75t_L g1963 ( 
.A(n_521),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_434),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_818),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_227),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_33),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_899),
.Y(n_1968)
);

CKINVDCx14_ASAP7_75t_R g1969 ( 
.A(n_302),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_79),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_773),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_870),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_168),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_874),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_272),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_891),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_142),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_878),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_235),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1153),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_856),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_347),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_261),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_446),
.Y(n_1984)
);

CKINVDCx14_ASAP7_75t_R g1985 ( 
.A(n_1080),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1129),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_608),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_1228),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_613),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_467),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1148),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1074),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_62),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_907),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1170),
.Y(n_1995)
);

CKINVDCx20_ASAP7_75t_R g1996 ( 
.A(n_238),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_784),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1184),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_147),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_175),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_655),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_945),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1235),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_38),
.Y(n_2004)
);

CKINVDCx20_ASAP7_75t_R g2005 ( 
.A(n_871),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_192),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1001),
.Y(n_2007)
);

INVxp33_ASAP7_75t_R g2008 ( 
.A(n_1152),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1247),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1043),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1030),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1020),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_513),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_554),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_1139),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1159),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_539),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_418),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_366),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_180),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1024),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1198),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_691),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_709),
.Y(n_2024)
);

INVxp67_ASAP7_75t_SL g2025 ( 
.A(n_164),
.Y(n_2025)
);

INVx1_ASAP7_75t_SL g2026 ( 
.A(n_645),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_626),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_156),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_984),
.Y(n_2029)
);

CKINVDCx14_ASAP7_75t_R g2030 ( 
.A(n_411),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_839),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_221),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1111),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1195),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_40),
.Y(n_2035)
);

BUFx10_ASAP7_75t_L g2036 ( 
.A(n_882),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_257),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_915),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_789),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1185),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_986),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_992),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_251),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_117),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_765),
.Y(n_2045)
);

CKINVDCx14_ASAP7_75t_R g2046 ( 
.A(n_46),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_305),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_583),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_804),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1042),
.Y(n_2050)
);

INVxp67_ASAP7_75t_L g2051 ( 
.A(n_33),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_604),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_236),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_908),
.Y(n_2054)
);

CKINVDCx20_ASAP7_75t_R g2055 ( 
.A(n_241),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_599),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_674),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_558),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_412),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_273),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_91),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_830),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1044),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1028),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_592),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_433),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_0),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1101),
.Y(n_2068)
);

CKINVDCx20_ASAP7_75t_R g2069 ( 
.A(n_316),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_532),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_191),
.Y(n_2071)
);

CKINVDCx20_ASAP7_75t_R g2072 ( 
.A(n_1175),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_470),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_64),
.Y(n_2074)
);

CKINVDCx14_ASAP7_75t_R g2075 ( 
.A(n_306),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_639),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_527),
.Y(n_2077)
);

CKINVDCx5p33_ASAP7_75t_R g2078 ( 
.A(n_853),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_841),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_753),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1144),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_438),
.Y(n_2082)
);

CKINVDCx16_ASAP7_75t_R g2083 ( 
.A(n_481),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1702),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1702),
.Y(n_2085)
);

INVxp67_ASAP7_75t_L g2086 ( 
.A(n_1305),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1702),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1702),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1702),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1787),
.Y(n_2090)
);

INVxp67_ASAP7_75t_SL g2091 ( 
.A(n_1798),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1384),
.Y(n_2092)
);

INVxp67_ASAP7_75t_SL g2093 ( 
.A(n_1833),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1787),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1787),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1487),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1787),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1787),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1566),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1566),
.Y(n_2100)
);

INVxp67_ASAP7_75t_SL g2101 ( 
.A(n_1731),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1577),
.Y(n_2102)
);

CKINVDCx20_ASAP7_75t_R g2103 ( 
.A(n_2081),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1294),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1294),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1294),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1306),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1306),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1306),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1602),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2083),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1602),
.Y(n_2112)
);

INVxp67_ASAP7_75t_SL g2113 ( 
.A(n_1779),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1602),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1609),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1609),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_1250),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1735),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1609),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1739),
.Y(n_2120)
);

BUFx2_ASAP7_75t_L g2121 ( 
.A(n_1867),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1739),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1473),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1739),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1865),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1865),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1865),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_1301),
.B(n_0),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1902),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1902),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1902),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2076),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1954),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1954),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1954),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1960),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1960),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_1435),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1724),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1960),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2024),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2024),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_1697),
.Y(n_2143)
);

INVxp33_ASAP7_75t_SL g2144 ( 
.A(n_1372),
.Y(n_2144)
);

CKINVDCx14_ASAP7_75t_R g2145 ( 
.A(n_1443),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2024),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2076),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2076),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2082),
.Y(n_2149)
);

BUFx10_ASAP7_75t_L g2150 ( 
.A(n_1428),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2082),
.Y(n_2151)
);

INVxp33_ASAP7_75t_L g2152 ( 
.A(n_1485),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_1254),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1268),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_1781),
.Y(n_2155)
);

INVxp33_ASAP7_75t_L g2156 ( 
.A(n_1666),
.Y(n_2156)
);

INVxp67_ASAP7_75t_SL g2157 ( 
.A(n_1478),
.Y(n_2157)
);

CKINVDCx20_ASAP7_75t_R g2158 ( 
.A(n_2072),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2082),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1357),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1969),
.B(n_2),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1445),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1277),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1492),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1575),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1603),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1606),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1642),
.Y(n_2168)
);

BUFx10_ASAP7_75t_L g2169 ( 
.A(n_1251),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1679),
.Y(n_2170)
);

INVxp33_ASAP7_75t_L g2171 ( 
.A(n_1504),
.Y(n_2171)
);

INVxp33_ASAP7_75t_L g2172 ( 
.A(n_1257),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1728),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1862),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1885),
.Y(n_2175)
);

INVxp33_ASAP7_75t_SL g2176 ( 
.A(n_1252),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1916),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1254),
.Y(n_2178)
);

INVxp33_ASAP7_75t_SL g2179 ( 
.A(n_1255),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1956),
.Y(n_2180)
);

INVxp67_ASAP7_75t_L g2181 ( 
.A(n_1403),
.Y(n_2181)
);

INVxp33_ASAP7_75t_L g2182 ( 
.A(n_1260),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1974),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1999),
.Y(n_2184)
);

INVxp33_ASAP7_75t_L g2185 ( 
.A(n_1261),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1270),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1382),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1285),
.Y(n_2188)
);

INVxp67_ASAP7_75t_SL g2189 ( 
.A(n_1478),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2071),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2073),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2030),
.B(n_3),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1286),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2079),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1382),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_1403),
.Y(n_2196)
);

INVxp33_ASAP7_75t_SL g2197 ( 
.A(n_1256),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1288),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1297),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1309),
.Y(n_2200)
);

CKINVDCx14_ASAP7_75t_R g2201 ( 
.A(n_2046),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1329),
.Y(n_2202)
);

INVxp67_ASAP7_75t_L g2203 ( 
.A(n_1408),
.Y(n_2203)
);

INVxp67_ASAP7_75t_L g2204 ( 
.A(n_1408),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1333),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_1785),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1382),
.Y(n_2207)
);

INVxp67_ASAP7_75t_L g2208 ( 
.A(n_1442),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_1302),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2062),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1290),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1338),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_1411),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1342),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1348),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1359),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1364),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_SL g2218 ( 
.A(n_1442),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1382),
.Y(n_2219)
);

BUFx2_ASAP7_75t_SL g2220 ( 
.A(n_1264),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1373),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1378),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_1376),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1382),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1392),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2061),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2060),
.Y(n_2227)
);

INVxp67_ASAP7_75t_SL g2228 ( 
.A(n_1448),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1397),
.Y(n_2229)
);

INVxp33_ASAP7_75t_SL g2230 ( 
.A(n_1258),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1543),
.Y(n_2231)
);

INVxp67_ASAP7_75t_SL g2232 ( 
.A(n_1570),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1410),
.Y(n_2233)
);

CKINVDCx20_ASAP7_75t_R g2234 ( 
.A(n_1282),
.Y(n_2234)
);

BUFx2_ASAP7_75t_L g2235 ( 
.A(n_2075),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1412),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1413),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1422),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1543),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1424),
.Y(n_2240)
);

INVxp33_ASAP7_75t_SL g2241 ( 
.A(n_1262),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1426),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1438),
.Y(n_2243)
);

INVxp33_ASAP7_75t_SL g2244 ( 
.A(n_1265),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1444),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_1283),
.B(n_1),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1450),
.Y(n_2247)
);

CKINVDCx16_ASAP7_75t_R g2248 ( 
.A(n_1457),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1452),
.Y(n_2249)
);

INVxp67_ASAP7_75t_L g2250 ( 
.A(n_1598),
.Y(n_2250)
);

CKINVDCx16_ASAP7_75t_R g2251 ( 
.A(n_1523),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1454),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1462),
.Y(n_2253)
);

INVx5_ASAP7_75t_L g2254 ( 
.A(n_2169),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2145),
.Y(n_2255)
);

INVx5_ASAP7_75t_L g2256 ( 
.A(n_2169),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2132),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_2159),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_2123),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2104),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2123),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2123),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_2111),
.Y(n_2263)
);

INVx5_ASAP7_75t_L g2264 ( 
.A(n_2150),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2105),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2106),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2107),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_2201),
.Y(n_2268)
);

OAI22x1_ASAP7_75t_SL g2269 ( 
.A1(n_2144),
.A2(n_1275),
.B1(n_1311),
.B2(n_1273),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2108),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_2213),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_2109),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2161),
.A2(n_1339),
.B1(n_1985),
.B2(n_1423),
.Y(n_2273)
);

INVxp67_ASAP7_75t_L g2274 ( 
.A(n_2117),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2110),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2112),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2114),
.Y(n_2277)
);

OAI21x1_ASAP7_75t_L g2278 ( 
.A1(n_2097),
.A2(n_1280),
.B(n_1279),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2115),
.Y(n_2279)
);

INVx3_ASAP7_75t_L g2280 ( 
.A(n_2213),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2153),
.Y(n_2281)
);

AOI22x1_ASAP7_75t_SL g2282 ( 
.A1(n_2103),
.A2(n_1366),
.B1(n_1446),
.B2(n_1344),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_2116),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2119),
.Y(n_2284)
);

INVx4_ASAP7_75t_L g2285 ( 
.A(n_2154),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2120),
.Y(n_2286)
);

INVxp33_ASAP7_75t_SL g2287 ( 
.A(n_2092),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_2122),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2124),
.Y(n_2289)
);

INVx6_ASAP7_75t_L g2290 ( 
.A(n_2150),
.Y(n_2290)
);

BUFx12f_ASAP7_75t_L g2291 ( 
.A(n_2102),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2138),
.B(n_1644),
.Y(n_2292)
);

AOI22xp5_ASAP7_75t_SL g2293 ( 
.A1(n_2171),
.A2(n_1500),
.B1(n_1514),
.B2(n_1496),
.Y(n_2293)
);

BUFx12f_ASAP7_75t_L g2294 ( 
.A(n_2139),
.Y(n_2294)
);

HB1xp67_ASAP7_75t_L g2295 ( 
.A(n_2143),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2125),
.Y(n_2296)
);

HB1xp67_ASAP7_75t_L g2297 ( 
.A(n_2155),
.Y(n_2297)
);

OAI21x1_ASAP7_75t_L g2298 ( 
.A1(n_2187),
.A2(n_1335),
.B(n_1317),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2126),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_2127),
.Y(n_2300)
);

BUFx6f_ASAP7_75t_L g2301 ( 
.A(n_2129),
.Y(n_2301)
);

INVx5_ASAP7_75t_L g2302 ( 
.A(n_2235),
.Y(n_2302)
);

CKINVDCx20_ASAP7_75t_R g2303 ( 
.A(n_2158),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2178),
.B(n_2101),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_2160),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2163),
.B(n_1322),
.Y(n_2306)
);

BUFx12f_ASAP7_75t_L g2307 ( 
.A(n_2193),
.Y(n_2307)
);

INVx6_ASAP7_75t_L g2308 ( 
.A(n_2248),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2130),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2209),
.B(n_1857),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_2206),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2226),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_2162),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2131),
.Y(n_2314)
);

INVxp33_ASAP7_75t_SL g2315 ( 
.A(n_2211),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_2133),
.Y(n_2316)
);

INVx2_ASAP7_75t_SL g2317 ( 
.A(n_2096),
.Y(n_2317)
);

BUFx12f_ASAP7_75t_L g2318 ( 
.A(n_2121),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_2134),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_2135),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2136),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2137),
.Y(n_2322)
);

BUFx12f_ASAP7_75t_L g2323 ( 
.A(n_2128),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2223),
.B(n_1920),
.Y(n_2324)
);

AND2x6_ASAP7_75t_L g2325 ( 
.A(n_2192),
.B(n_1259),
.Y(n_2325)
);

OA21x2_ASAP7_75t_L g2326 ( 
.A1(n_2084),
.A2(n_1863),
.B(n_1416),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2140),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2141),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2142),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2146),
.Y(n_2330)
);

INVx5_ASAP7_75t_L g2331 ( 
.A(n_2251),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2147),
.Y(n_2332)
);

BUFx12f_ASAP7_75t_L g2333 ( 
.A(n_2246),
.Y(n_2333)
);

AND2x4_ASAP7_75t_L g2334 ( 
.A(n_2113),
.B(n_1639),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2148),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2149),
.Y(n_2336)
);

INVx5_ASAP7_75t_L g2337 ( 
.A(n_2195),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2151),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2085),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2186),
.Y(n_2340)
);

AOI22x1_ASAP7_75t_SL g2341 ( 
.A1(n_2234),
.A2(n_1571),
.B1(n_1592),
.B2(n_1537),
.Y(n_2341)
);

INVx5_ASAP7_75t_L g2342 ( 
.A(n_2207),
.Y(n_2342)
);

BUFx6f_ASAP7_75t_L g2343 ( 
.A(n_2188),
.Y(n_2343)
);

AND2x4_ASAP7_75t_L g2344 ( 
.A(n_2228),
.B(n_1682),
.Y(n_2344)
);

INVxp67_ASAP7_75t_SL g2345 ( 
.A(n_2232),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2091),
.B(n_1820),
.Y(n_2346)
);

BUFx6f_ASAP7_75t_L g2347 ( 
.A(n_2190),
.Y(n_2347)
);

BUFx3_ASAP7_75t_L g2348 ( 
.A(n_2164),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2093),
.A2(n_1341),
.B1(n_1365),
.B2(n_1308),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2087),
.Y(n_2350)
);

INVx5_ASAP7_75t_L g2351 ( 
.A(n_2219),
.Y(n_2351)
);

OAI22x1_ASAP7_75t_R g2352 ( 
.A1(n_2191),
.A2(n_1630),
.B1(n_1638),
.B2(n_1608),
.Y(n_2352)
);

INVx4_ASAP7_75t_L g2353 ( 
.A(n_2218),
.Y(n_2353)
);

BUFx8_ASAP7_75t_L g2354 ( 
.A(n_2218),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2088),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2089),
.Y(n_2356)
);

INVx3_ASAP7_75t_L g2357 ( 
.A(n_2165),
.Y(n_2357)
);

BUFx8_ASAP7_75t_L g2358 ( 
.A(n_2166),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_2167),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2194),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2090),
.Y(n_2361)
);

INVx5_ASAP7_75t_L g2362 ( 
.A(n_2224),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2152),
.B(n_1267),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2181),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_2196),
.Y(n_2365)
);

CKINVDCx16_ASAP7_75t_R g2366 ( 
.A(n_2220),
.Y(n_2366)
);

BUFx6f_ASAP7_75t_L g2367 ( 
.A(n_2198),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2157),
.B(n_1625),
.Y(n_2368)
);

OA21x2_ASAP7_75t_L g2369 ( 
.A1(n_2094),
.A2(n_1269),
.B(n_1253),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2095),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2098),
.Y(n_2371)
);

BUFx8_ASAP7_75t_SL g2372 ( 
.A(n_2168),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_2199),
.Y(n_2373)
);

BUFx2_ASAP7_75t_L g2374 ( 
.A(n_2203),
.Y(n_2374)
);

BUFx3_ASAP7_75t_L g2375 ( 
.A(n_2170),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2086),
.B(n_1336),
.Y(n_2376)
);

BUFx6f_ASAP7_75t_L g2377 ( 
.A(n_2200),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2118),
.B(n_1407),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_2173),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2176),
.A2(n_1460),
.B1(n_1546),
.B2(n_1368),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_2189),
.B(n_1420),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_2179),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2202),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_2205),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_2156),
.B(n_2172),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_2204),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2099),
.Y(n_2387)
);

OAI22xp5_ASAP7_75t_SL g2388 ( 
.A1(n_2208),
.A2(n_1699),
.B1(n_1705),
.B2(n_1641),
.Y(n_2388)
);

INVx5_ASAP7_75t_L g2389 ( 
.A(n_2231),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2174),
.B(n_1790),
.Y(n_2390)
);

BUFx2_ASAP7_75t_L g2391 ( 
.A(n_2250),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2175),
.B(n_1793),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2197),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2230),
.Y(n_2394)
);

INVx5_ASAP7_75t_L g2395 ( 
.A(n_2239),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2100),
.Y(n_2396)
);

BUFx12f_ASAP7_75t_L g2397 ( 
.A(n_2241),
.Y(n_2397)
);

BUFx12f_ASAP7_75t_L g2398 ( 
.A(n_2244),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_2210),
.Y(n_2399)
);

INVx6_ASAP7_75t_L g2400 ( 
.A(n_2182),
.Y(n_2400)
);

HB1xp67_ASAP7_75t_L g2401 ( 
.A(n_2177),
.Y(n_2401)
);

INVx5_ASAP7_75t_L g2402 ( 
.A(n_2185),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2212),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2180),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2214),
.Y(n_2405)
);

CKINVDCx16_ASAP7_75t_R g2406 ( 
.A(n_2183),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2215),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2184),
.Y(n_2408)
);

INVx4_ASAP7_75t_L g2409 ( 
.A(n_2216),
.Y(n_2409)
);

INVx4_ASAP7_75t_L g2410 ( 
.A(n_2217),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2221),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_2222),
.Y(n_2412)
);

BUFx12f_ASAP7_75t_L g2413 ( 
.A(n_2225),
.Y(n_2413)
);

INVx2_ASAP7_75t_SL g2414 ( 
.A(n_2227),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2229),
.Y(n_2415)
);

OAI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2233),
.A2(n_1398),
.B1(n_2051),
.B2(n_1358),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2236),
.B(n_1267),
.Y(n_2417)
);

INVx3_ASAP7_75t_L g2418 ( 
.A(n_2237),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2238),
.Y(n_2419)
);

BUFx6f_ASAP7_75t_L g2420 ( 
.A(n_2240),
.Y(n_2420)
);

BUFx2_ASAP7_75t_L g2421 ( 
.A(n_2242),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_2243),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2245),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2247),
.B(n_1562),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2249),
.Y(n_2425)
);

BUFx12f_ASAP7_75t_L g2426 ( 
.A(n_2252),
.Y(n_2426)
);

BUFx2_ASAP7_75t_L g2427 ( 
.A(n_2253),
.Y(n_2427)
);

CKINVDCx16_ASAP7_75t_R g2428 ( 
.A(n_2145),
.Y(n_2428)
);

INVx4_ASAP7_75t_L g2429 ( 
.A(n_2154),
.Y(n_2429)
);

BUFx8_ASAP7_75t_SL g2430 ( 
.A(n_2218),
.Y(n_2430)
);

AOI22xp5_ASAP7_75t_L g2431 ( 
.A1(n_2144),
.A2(n_1636),
.B1(n_1659),
.B2(n_1586),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2132),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_2132),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2160),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2132),
.Y(n_2435)
);

BUFx2_ASAP7_75t_L g2436 ( 
.A(n_2145),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2111),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2132),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2132),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2132),
.Y(n_2440)
);

BUFx6f_ASAP7_75t_L g2441 ( 
.A(n_2132),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2132),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2132),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2132),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2132),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2132),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2145),
.B(n_1377),
.Y(n_2447)
);

INVx2_ASAP7_75t_SL g2448 ( 
.A(n_2169),
.Y(n_2448)
);

INVx2_ASAP7_75t_SL g2449 ( 
.A(n_2169),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2132),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2132),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2132),
.Y(n_2452)
);

INVx3_ASAP7_75t_L g2453 ( 
.A(n_2132),
.Y(n_2453)
);

AND2x4_ASAP7_75t_L g2454 ( 
.A(n_2138),
.B(n_1811),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2154),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2132),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2132),
.Y(n_2457)
);

BUFx6f_ASAP7_75t_L g2458 ( 
.A(n_2132),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2138),
.B(n_1823),
.Y(n_2459)
);

BUFx3_ASAP7_75t_L g2460 ( 
.A(n_2160),
.Y(n_2460)
);

INVx5_ASAP7_75t_L g2461 ( 
.A(n_2169),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2132),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2132),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2132),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2132),
.Y(n_2465)
);

CKINVDCx20_ASAP7_75t_R g2466 ( 
.A(n_2103),
.Y(n_2466)
);

CKINVDCx20_ASAP7_75t_R g2467 ( 
.A(n_2103),
.Y(n_2467)
);

HB1xp67_ASAP7_75t_L g2468 ( 
.A(n_2111),
.Y(n_2468)
);

AND2x4_ASAP7_75t_L g2469 ( 
.A(n_2138),
.B(n_1901),
.Y(n_2469)
);

BUFx6f_ASAP7_75t_L g2470 ( 
.A(n_2132),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2160),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2154),
.Y(n_2472)
);

BUFx12f_ASAP7_75t_L g2473 ( 
.A(n_2092),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2132),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2160),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2154),
.B(n_1878),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2154),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2132),
.Y(n_2478)
);

BUFx12f_ASAP7_75t_L g2479 ( 
.A(n_2092),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2132),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2132),
.Y(n_2481)
);

BUFx6f_ASAP7_75t_L g2482 ( 
.A(n_2132),
.Y(n_2482)
);

INVx5_ASAP7_75t_L g2483 ( 
.A(n_2169),
.Y(n_2483)
);

INVx5_ASAP7_75t_L g2484 ( 
.A(n_2169),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2132),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2132),
.Y(n_2486)
);

INVx5_ASAP7_75t_L g2487 ( 
.A(n_2169),
.Y(n_2487)
);

BUFx12f_ASAP7_75t_L g2488 ( 
.A(n_2092),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2132),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2132),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2138),
.B(n_1917),
.Y(n_2491)
);

HB1xp67_ASAP7_75t_L g2492 ( 
.A(n_2111),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_2132),
.Y(n_2493)
);

BUFx3_ASAP7_75t_L g2494 ( 
.A(n_2160),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_2132),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2160),
.Y(n_2496)
);

BUFx12f_ASAP7_75t_L g2497 ( 
.A(n_2092),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2132),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2132),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2132),
.Y(n_2500)
);

BUFx8_ASAP7_75t_SL g2501 ( 
.A(n_2218),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2132),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2132),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2132),
.Y(n_2504)
);

INVx2_ASAP7_75t_SL g2505 ( 
.A(n_2169),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2132),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2132),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_2132),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_2154),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2132),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2132),
.Y(n_2511)
);

BUFx3_ASAP7_75t_L g2512 ( 
.A(n_2160),
.Y(n_2512)
);

BUFx2_ASAP7_75t_L g2513 ( 
.A(n_2145),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2132),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2132),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2132),
.Y(n_2516)
);

AND2x4_ASAP7_75t_L g2517 ( 
.A(n_2138),
.B(n_1991),
.Y(n_2517)
);

OAI21xp33_ASAP7_75t_L g2518 ( 
.A1(n_2152),
.A2(n_1481),
.B(n_1477),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2154),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2132),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2138),
.B(n_1263),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2132),
.Y(n_2522)
);

BUFx8_ASAP7_75t_SL g2523 ( 
.A(n_2218),
.Y(n_2523)
);

AOI22x1_ASAP7_75t_SL g2524 ( 
.A1(n_2103),
.A2(n_1771),
.B1(n_1772),
.B2(n_1716),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_2132),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2132),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2132),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2132),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2132),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2145),
.B(n_1377),
.Y(n_2530)
);

BUFx3_ASAP7_75t_L g2531 ( 
.A(n_2160),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2154),
.Y(n_2532)
);

INVxp67_ASAP7_75t_L g2533 ( 
.A(n_2111),
.Y(n_2533)
);

OAI22x1_ASAP7_75t_SL g2534 ( 
.A1(n_2144),
.A2(n_1836),
.B1(n_1843),
.B2(n_1817),
.Y(n_2534)
);

BUFx8_ASAP7_75t_SL g2535 ( 
.A(n_2218),
.Y(n_2535)
);

NOR2xp67_ASAP7_75t_L g2536 ( 
.A(n_2154),
.B(n_1955),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2111),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2138),
.B(n_1986),
.Y(n_2538)
);

AOI22x1_ASAP7_75t_SL g2539 ( 
.A1(n_2103),
.A2(n_1869),
.B1(n_1870),
.B2(n_1847),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2132),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_2132),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2132),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2132),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2132),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2132),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_SL g2546 ( 
.A(n_2248),
.B(n_1391),
.Y(n_2546)
);

INVx4_ASAP7_75t_L g2547 ( 
.A(n_2154),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2154),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_2132),
.Y(n_2549)
);

OAI21x1_ASAP7_75t_L g2550 ( 
.A1(n_2097),
.A2(n_1347),
.B(n_1345),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2132),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2132),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2132),
.Y(n_2553)
);

HB1xp67_ASAP7_75t_L g2554 ( 
.A(n_2111),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2138),
.B(n_1284),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2144),
.A2(n_1753),
.B1(n_1769),
.B2(n_1678),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2132),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2132),
.Y(n_2558)
);

AND2x4_ASAP7_75t_L g2559 ( 
.A(n_2138),
.B(n_1289),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2132),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2132),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2132),
.Y(n_2562)
);

BUFx6f_ASAP7_75t_L g2563 ( 
.A(n_2132),
.Y(n_2563)
);

OA21x2_ASAP7_75t_L g2564 ( 
.A1(n_2084),
.A2(n_1299),
.B(n_1296),
.Y(n_2564)
);

BUFx8_ASAP7_75t_SL g2565 ( 
.A(n_2218),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_SL g2566 ( 
.A1(n_2144),
.A2(n_1879),
.B1(n_1896),
.B2(n_1872),
.Y(n_2566)
);

INVxp67_ASAP7_75t_L g2567 ( 
.A(n_2111),
.Y(n_2567)
);

INVx5_ASAP7_75t_L g2568 ( 
.A(n_2169),
.Y(n_2568)
);

AND2x6_ASAP7_75t_L g2569 ( 
.A(n_2161),
.B(n_1303),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2132),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2132),
.Y(n_2571)
);

BUFx8_ASAP7_75t_SL g2572 ( 
.A(n_2218),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2176),
.B(n_1313),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2132),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2132),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2138),
.B(n_1327),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2132),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2154),
.B(n_1351),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2154),
.B(n_1355),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2132),
.Y(n_2580)
);

OAI22xp5_ASAP7_75t_L g2581 ( 
.A1(n_2144),
.A2(n_1271),
.B1(n_1272),
.B2(n_1266),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2171),
.B(n_1391),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2154),
.B(n_1509),
.Y(n_2583)
);

CKINVDCx20_ASAP7_75t_R g2584 ( 
.A(n_2303),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2345),
.B(n_1300),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2405),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2344),
.B(n_1794),
.Y(n_2587)
);

CKINVDCx20_ASAP7_75t_R g2588 ( 
.A(n_2466),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2261),
.Y(n_2589)
);

BUFx8_ASAP7_75t_L g2590 ( 
.A(n_2291),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2407),
.Y(n_2591)
);

BUFx6f_ASAP7_75t_L g2592 ( 
.A(n_2259),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2455),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2472),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2419),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2310),
.B(n_1316),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2477),
.Y(n_2597)
);

CKINVDCx20_ASAP7_75t_R g2598 ( 
.A(n_2467),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2324),
.B(n_1319),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2340),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2343),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2262),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2385),
.B(n_2400),
.Y(n_2603)
);

INVxp67_ASAP7_75t_L g2604 ( 
.A(n_2363),
.Y(n_2604)
);

BUFx3_ASAP7_75t_L g2605 ( 
.A(n_2305),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2402),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2258),
.Y(n_2607)
);

NAND2x1_ASAP7_75t_L g2608 ( 
.A(n_2369),
.B(n_1473),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2433),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2263),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2509),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2578),
.B(n_1324),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2519),
.Y(n_2613)
);

CKINVDCx20_ASAP7_75t_R g2614 ( 
.A(n_2366),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2347),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2532),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2548),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2579),
.B(n_1325),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2315),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2360),
.Y(n_2620)
);

BUFx6f_ASAP7_75t_L g2621 ( 
.A(n_2438),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2441),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2367),
.Y(n_2623)
);

CKINVDCx20_ASAP7_75t_R g2624 ( 
.A(n_2428),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2373),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2281),
.B(n_1808),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_2307),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2377),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2287),
.Y(n_2629)
);

CKINVDCx20_ASAP7_75t_R g2630 ( 
.A(n_2308),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_2294),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2334),
.B(n_1850),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2384),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2304),
.B(n_1859),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2399),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_2473),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2411),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2457),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2479),
.Y(n_2639)
);

NAND2xp33_ASAP7_75t_R g2640 ( 
.A(n_2365),
.B(n_2374),
.Y(n_2640)
);

CKINVDCx5p33_ASAP7_75t_R g2641 ( 
.A(n_2488),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2412),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2420),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2350),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2356),
.Y(n_2645)
);

OAI21x1_ASAP7_75t_L g2646 ( 
.A1(n_2278),
.A2(n_1541),
.B(n_1510),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2370),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2497),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_2382),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2339),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2355),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2295),
.Y(n_2652)
);

AND2x2_ASAP7_75t_SL g2653 ( 
.A(n_2546),
.B(n_1310),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2361),
.Y(n_2654)
);

NAND2xp33_ASAP7_75t_SL g2655 ( 
.A(n_2292),
.B(n_1930),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2458),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2371),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2393),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2313),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2348),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2583),
.B(n_1326),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2394),
.Y(n_2662)
);

INVx3_ASAP7_75t_L g2663 ( 
.A(n_2462),
.Y(n_2663)
);

BUFx6f_ASAP7_75t_L g2664 ( 
.A(n_2470),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2381),
.B(n_1598),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_2397),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2536),
.B(n_2573),
.Y(n_2667)
);

INVxp67_ASAP7_75t_L g2668 ( 
.A(n_2364),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2375),
.Y(n_2669)
);

CKINVDCx20_ASAP7_75t_R g2670 ( 
.A(n_2331),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2434),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_2555),
.B(n_2015),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2317),
.B(n_1447),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_2398),
.Y(n_2674)
);

BUFx6f_ASAP7_75t_L g2675 ( 
.A(n_2474),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2297),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_2285),
.Y(n_2677)
);

CKINVDCx5p33_ASAP7_75t_R g2678 ( 
.A(n_2429),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_R g2679 ( 
.A(n_2255),
.B(n_1332),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2482),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2486),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2460),
.Y(n_2682)
);

CKINVDCx5p33_ASAP7_75t_R g2683 ( 
.A(n_2547),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2471),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2475),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2376),
.B(n_1667),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2368),
.B(n_1349),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2430),
.Y(n_2688)
);

CKINVDCx20_ASAP7_75t_R g2689 ( 
.A(n_2268),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2501),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2494),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2496),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2493),
.Y(n_2693)
);

AND2x4_ASAP7_75t_L g2694 ( 
.A(n_2559),
.B(n_1726),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2523),
.Y(n_2695)
);

BUFx6f_ASAP7_75t_L g2696 ( 
.A(n_2495),
.Y(n_2696)
);

CKINVDCx20_ASAP7_75t_R g2697 ( 
.A(n_2436),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2535),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2325),
.A2(n_2025),
.B1(n_1499),
.B2(n_1559),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_L g2700 ( 
.A(n_2346),
.B(n_1276),
.C(n_1274),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2512),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2498),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2500),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2531),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2387),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2504),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2396),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2525),
.Y(n_2708)
);

CKINVDCx20_ASAP7_75t_R g2709 ( 
.A(n_2513),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2565),
.Y(n_2710)
);

BUFx6f_ASAP7_75t_L g2711 ( 
.A(n_2526),
.Y(n_2711)
);

BUFx2_ASAP7_75t_L g2712 ( 
.A(n_2318),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2572),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2576),
.B(n_1810),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2527),
.Y(n_2715)
);

CKINVDCx5p33_ASAP7_75t_R g2716 ( 
.A(n_2254),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2454),
.B(n_1518),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2383),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_2541),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2403),
.Y(n_2720)
);

NOR2xp67_ASAP7_75t_L g2721 ( 
.A(n_2256),
.B(n_1350),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2415),
.Y(n_2722)
);

CKINVDCx20_ASAP7_75t_R g2723 ( 
.A(n_2380),
.Y(n_2723)
);

CKINVDCx20_ASAP7_75t_R g2724 ( 
.A(n_2406),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_2545),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2461),
.Y(n_2726)
);

NAND3xp33_ASAP7_75t_L g2727 ( 
.A(n_2421),
.B(n_1281),
.C(n_1278),
.Y(n_2727)
);

HB1xp67_ASAP7_75t_L g2728 ( 
.A(n_2437),
.Y(n_2728)
);

CKINVDCx20_ASAP7_75t_R g2729 ( 
.A(n_2431),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2483),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2425),
.Y(n_2731)
);

HB1xp67_ASAP7_75t_L g2732 ( 
.A(n_2468),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2459),
.B(n_1518),
.Y(n_2733)
);

AND2x2_ASAP7_75t_L g2734 ( 
.A(n_2378),
.B(n_1667),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2414),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2549),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2551),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2484),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2401),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2408),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2427),
.B(n_2070),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2487),
.Y(n_2742)
);

AND2x4_ASAP7_75t_L g2743 ( 
.A(n_2302),
.B(n_1464),
.Y(n_2743)
);

CKINVDCx20_ASAP7_75t_R g2744 ( 
.A(n_2556),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2418),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2422),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2260),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2568),
.Y(n_2748)
);

BUFx6f_ASAP7_75t_L g2749 ( 
.A(n_2557),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2306),
.B(n_1354),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2349),
.Y(n_2751)
);

INVxp67_ASAP7_75t_L g2752 ( 
.A(n_2386),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2469),
.B(n_1883),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2563),
.Y(n_2754)
);

BUFx6f_ASAP7_75t_L g2755 ( 
.A(n_2570),
.Y(n_2755)
);

CKINVDCx20_ASAP7_75t_R g2756 ( 
.A(n_2492),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2354),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2333),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2265),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2266),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2323),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2267),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_2448),
.Y(n_2763)
);

NOR2xp67_ASAP7_75t_L g2764 ( 
.A(n_2449),
.B(n_1356),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2476),
.B(n_1360),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2577),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2491),
.B(n_1883),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2505),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2302),
.B(n_1483),
.Y(n_2769)
);

BUFx10_ASAP7_75t_L g2770 ( 
.A(n_2290),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2372),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2270),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2435),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2279),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2326),
.B(n_1370),
.Y(n_2775)
);

CKINVDCx16_ASAP7_75t_R g2776 ( 
.A(n_2352),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2440),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2296),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_SL g2779 ( 
.A(n_2517),
.B(n_1563),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2442),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2443),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2273),
.B(n_1399),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_2391),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_2413),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2521),
.B(n_1494),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2426),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2299),
.Y(n_2787)
);

XOR2xp5_ASAP7_75t_L g2788 ( 
.A(n_2282),
.B(n_1400),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2272),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_L g2790 ( 
.A(n_2283),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2452),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2463),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2309),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_L g2794 ( 
.A(n_2284),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2464),
.Y(n_2795)
);

CKINVDCx5p33_ASAP7_75t_R g2796 ( 
.A(n_2341),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2314),
.Y(n_2797)
);

CKINVDCx20_ASAP7_75t_R g2798 ( 
.A(n_2537),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2337),
.B(n_1401),
.Y(n_2799)
);

AND2x6_ASAP7_75t_L g2800 ( 
.A(n_2447),
.B(n_1473),
.Y(n_2800)
);

CKINVDCx5p33_ASAP7_75t_R g2801 ( 
.A(n_2524),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2329),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2478),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_R g2804 ( 
.A(n_2530),
.B(n_1404),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2330),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_2539),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_2325),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2338),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2480),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2424),
.B(n_1563),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2481),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2312),
.B(n_2274),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2502),
.Y(n_2813)
);

CKINVDCx20_ASAP7_75t_R g2814 ( 
.A(n_2554),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2300),
.Y(n_2815)
);

AND2x4_ASAP7_75t_L g2816 ( 
.A(n_2538),
.B(n_2423),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2503),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2311),
.B(n_1909),
.Y(n_2818)
);

BUFx6f_ASAP7_75t_L g2819 ( 
.A(n_2301),
.Y(n_2819)
);

INVxp67_ASAP7_75t_L g2820 ( 
.A(n_2582),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2533),
.B(n_1909),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2510),
.Y(n_2822)
);

OAI21x1_ASAP7_75t_L g2823 ( 
.A1(n_2550),
.A2(n_1560),
.B(n_1550),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2567),
.B(n_2008),
.Y(n_2824)
);

CKINVDCx20_ASAP7_75t_R g2825 ( 
.A(n_2293),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2516),
.Y(n_2826)
);

CKINVDCx20_ASAP7_75t_R g2827 ( 
.A(n_2566),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_R g2828 ( 
.A(n_2353),
.B(n_1406),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_2569),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2522),
.Y(n_2830)
);

CKINVDCx5p33_ASAP7_75t_R g2831 ( 
.A(n_2569),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2581),
.Y(n_2832)
);

CKINVDCx5p33_ASAP7_75t_R g2833 ( 
.A(n_2264),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2540),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2316),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2417),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2543),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2544),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2388),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2558),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2560),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2404),
.A2(n_1291),
.B1(n_1292),
.B2(n_1287),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2561),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_2269),
.Y(n_2844)
);

BUFx8_ASAP7_75t_L g2845 ( 
.A(n_2534),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_2358),
.Y(n_2846)
);

AND2x6_ASAP7_75t_L g2847 ( 
.A(n_2357),
.B(n_1497),
.Y(n_2847)
);

INVxp67_ASAP7_75t_L g2848 ( 
.A(n_2390),
.Y(n_2848)
);

AND2x4_ASAP7_75t_L g2849 ( 
.A(n_2359),
.B(n_1503),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2562),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2409),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2571),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2319),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2416),
.Y(n_2854)
);

OA21x2_ASAP7_75t_L g2855 ( 
.A1(n_2298),
.A2(n_1694),
.B(n_1600),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2379),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2275),
.Y(n_2857)
);

CKINVDCx20_ASAP7_75t_R g2858 ( 
.A(n_2392),
.Y(n_2858)
);

CKINVDCx20_ASAP7_75t_R g2859 ( 
.A(n_2518),
.Y(n_2859)
);

HB1xp67_ASAP7_75t_L g2860 ( 
.A(n_2320),
.Y(n_2860)
);

BUFx3_ASAP7_75t_L g2861 ( 
.A(n_2342),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2288),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2276),
.Y(n_2863)
);

AND2x4_ASAP7_75t_L g2864 ( 
.A(n_2271),
.B(n_1507),
.Y(n_2864)
);

NAND2xp33_ASAP7_75t_L g2865 ( 
.A(n_2321),
.B(n_1497),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2277),
.Y(n_2866)
);

OAI22xp5_ASAP7_75t_SL g2867 ( 
.A1(n_2280),
.A2(n_1996),
.B1(n_2005),
.B2(n_1965),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2286),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2289),
.Y(n_2869)
);

NAND2xp33_ASAP7_75t_L g2870 ( 
.A(n_2332),
.B(n_1497),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2453),
.Y(n_2871)
);

INVxp67_ASAP7_75t_L g2872 ( 
.A(n_2508),
.Y(n_2872)
);

INVx1_ASAP7_75t_SL g2873 ( 
.A(n_2514),
.Y(n_2873)
);

INVx3_ASAP7_75t_L g2874 ( 
.A(n_2410),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2322),
.Y(n_2875)
);

BUFx6f_ASAP7_75t_L g2876 ( 
.A(n_2327),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_2328),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2335),
.Y(n_2878)
);

CKINVDCx20_ASAP7_75t_R g2879 ( 
.A(n_2564),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2336),
.Y(n_2880)
);

CKINVDCx20_ASAP7_75t_R g2881 ( 
.A(n_2351),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2362),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2389),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2257),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2432),
.Y(n_2885)
);

OA21x2_ASAP7_75t_L g2886 ( 
.A1(n_2439),
.A2(n_1922),
.B(n_1838),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_2444),
.Y(n_2887)
);

CKINVDCx5p33_ASAP7_75t_R g2888 ( 
.A(n_2445),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2395),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2446),
.Y(n_2890)
);

CKINVDCx20_ASAP7_75t_R g2891 ( 
.A(n_2450),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_2451),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2456),
.B(n_1293),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_2465),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2485),
.B(n_1414),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2489),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2586),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2848),
.B(n_1328),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2591),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2773),
.Y(n_2900)
);

OAI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_2879),
.A2(n_1968),
.B1(n_2038),
.B2(n_1957),
.Y(n_2901)
);

NOR2x1p5_ASAP7_75t_L g2902 ( 
.A(n_2786),
.B(n_1295),
.Y(n_2902)
);

BUFx10_ASAP7_75t_L g2903 ( 
.A(n_2688),
.Y(n_2903)
);

BUFx4f_ASAP7_75t_L g2904 ( 
.A(n_2653),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2595),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2777),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_2593),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2667),
.B(n_1421),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2780),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2603),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2781),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2604),
.B(n_1432),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2791),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2644),
.A2(n_1581),
.B1(n_1683),
.B2(n_1390),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_2792),
.Y(n_2915)
);

INVxp67_ASAP7_75t_L g2916 ( 
.A(n_2673),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2816),
.B(n_1434),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2795),
.Y(n_2918)
);

OAI22xp33_ASAP7_75t_L g2919 ( 
.A1(n_2699),
.A2(n_1565),
.B1(n_1710),
.B2(n_1468),
.Y(n_2919)
);

BUFx2_ASAP7_75t_L g2920 ( 
.A(n_2756),
.Y(n_2920)
);

AND2x6_ASAP7_75t_L g2921 ( 
.A(n_2665),
.B(n_1337),
.Y(n_2921)
);

INVx3_ASAP7_75t_L g2922 ( 
.A(n_2592),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2789),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2705),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2803),
.Y(n_2925)
);

NAND2xp33_ASAP7_75t_SL g2926 ( 
.A(n_2859),
.B(n_2049),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_L g2927 ( 
.A(n_2820),
.B(n_1729),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2596),
.B(n_1437),
.Y(n_2928)
);

INVx3_ASAP7_75t_L g2929 ( 
.A(n_2592),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2822),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2834),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2707),
.Y(n_2932)
);

BUFx10_ASAP7_75t_L g2933 ( 
.A(n_2690),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2852),
.Y(n_2934)
);

INVx1_ASAP7_75t_SL g2935 ( 
.A(n_2798),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2857),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_2594),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2609),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2866),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2612),
.B(n_1363),
.Y(n_2940)
);

CKINVDCx5p33_ASAP7_75t_R g2941 ( 
.A(n_2597),
.Y(n_2941)
);

INVx3_ASAP7_75t_L g2942 ( 
.A(n_2609),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2747),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2759),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2868),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2869),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2875),
.Y(n_2947)
);

INVxp67_ASAP7_75t_SL g2948 ( 
.A(n_2872),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2686),
.B(n_2490),
.Y(n_2949)
);

NAND2xp33_ASAP7_75t_SL g2950 ( 
.A(n_2807),
.B(n_2055),
.Y(n_2950)
);

INVx2_ASAP7_75t_SL g2951 ( 
.A(n_2610),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2618),
.B(n_1371),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2650),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2651),
.Y(n_2954)
);

NOR2xp33_ASAP7_75t_L g2955 ( 
.A(n_2668),
.B(n_1733),
.Y(n_2955)
);

INVx2_ASAP7_75t_SL g2956 ( 
.A(n_2652),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2752),
.B(n_1866),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2585),
.B(n_1890),
.Y(n_2958)
);

INVx3_ASAP7_75t_L g2959 ( 
.A(n_2621),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2654),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2760),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2657),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2762),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2809),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2811),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2813),
.Y(n_2966)
);

NOR2x1p5_ASAP7_75t_L g2967 ( 
.A(n_2784),
.B(n_2846),
.Y(n_2967)
);

NAND3xp33_ASAP7_75t_L g2968 ( 
.A(n_2700),
.B(n_1304),
.C(n_1298),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2772),
.Y(n_2969)
);

CKINVDCx5p33_ASAP7_75t_R g2970 ( 
.A(n_2611),
.Y(n_2970)
);

BUFx10_ASAP7_75t_L g2971 ( 
.A(n_2695),
.Y(n_2971)
);

BUFx6f_ASAP7_75t_L g2972 ( 
.A(n_2621),
.Y(n_2972)
);

AND2x6_ASAP7_75t_L g2973 ( 
.A(n_2753),
.B(n_1375),
.Y(n_2973)
);

INVx2_ASAP7_75t_SL g2974 ( 
.A(n_2676),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2817),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2728),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2599),
.B(n_1900),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2826),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2661),
.B(n_1386),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2830),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2664),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_2677),
.B(n_1441),
.Y(n_2982)
);

BUFx3_ASAP7_75t_L g2983 ( 
.A(n_2630),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2837),
.Y(n_2984)
);

INVx4_ASAP7_75t_L g2985 ( 
.A(n_2789),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2838),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2840),
.Y(n_2987)
);

BUFx2_ASAP7_75t_L g2988 ( 
.A(n_2814),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2774),
.Y(n_2989)
);

INVx3_ASAP7_75t_L g2990 ( 
.A(n_2664),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2841),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2778),
.Y(n_2992)
);

BUFx6f_ASAP7_75t_L g2993 ( 
.A(n_2675),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2787),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2843),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2850),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2793),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2718),
.Y(n_2998)
);

BUFx2_ASAP7_75t_L g2999 ( 
.A(n_2724),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_2678),
.B(n_1449),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_2734),
.B(n_2499),
.Y(n_3001)
);

BUFx2_ASAP7_75t_L g3002 ( 
.A(n_2732),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2675),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2720),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2797),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2683),
.B(n_1455),
.Y(n_3006)
);

BUFx2_ASAP7_75t_L g3007 ( 
.A(n_2783),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2696),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2645),
.B(n_1415),
.Y(n_3009)
);

AOI22xp5_ASAP7_75t_L g3010 ( 
.A1(n_2832),
.A2(n_1459),
.B1(n_1461),
.B2(n_1458),
.Y(n_3010)
);

BUFx2_ASAP7_75t_L g3011 ( 
.A(n_2626),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2836),
.B(n_1467),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2722),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2731),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_L g3015 ( 
.A(n_2696),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2885),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2802),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_2711),
.Y(n_3018)
);

BUFx6f_ASAP7_75t_SL g3019 ( 
.A(n_2770),
.Y(n_3019)
);

OR2x6_ASAP7_75t_L g3020 ( 
.A(n_2712),
.B(n_1520),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2750),
.B(n_1948),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2805),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2647),
.B(n_1419),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2808),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2812),
.B(n_2767),
.Y(n_3025)
);

INVx5_ASAP7_75t_L g3026 ( 
.A(n_2790),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2896),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2863),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_L g3029 ( 
.A(n_2711),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2878),
.Y(n_3030)
);

INVx2_ASAP7_75t_SL g3031 ( 
.A(n_2743),
.Y(n_3031)
);

INVx3_ASAP7_75t_L g3032 ( 
.A(n_2719),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2890),
.Y(n_3033)
);

OR2x6_ASAP7_75t_L g3034 ( 
.A(n_2606),
.B(n_1526),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2880),
.Y(n_3035)
);

INVx4_ASAP7_75t_L g3036 ( 
.A(n_2790),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2589),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2602),
.Y(n_3038)
);

INVx5_ASAP7_75t_L g3039 ( 
.A(n_2794),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2745),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2894),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2894),
.Y(n_3042)
);

INVx4_ASAP7_75t_L g3043 ( 
.A(n_2794),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_2782),
.B(n_1475),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2775),
.A2(n_1431),
.B1(n_1436),
.B2(n_1429),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2746),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2862),
.Y(n_3047)
);

OR2x6_ASAP7_75t_L g3048 ( 
.A(n_2672),
.B(n_1530),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2856),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2864),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2860),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2818),
.B(n_2506),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2687),
.B(n_1439),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2871),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2821),
.B(n_2507),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2804),
.B(n_1484),
.Y(n_3056)
);

AOI21x1_ASAP7_75t_L g3057 ( 
.A1(n_2608),
.A2(n_2515),
.B(n_2511),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2876),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2876),
.Y(n_3059)
);

INVx3_ASAP7_75t_L g3060 ( 
.A(n_2719),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2871),
.Y(n_3061)
);

OAI22x1_ASAP7_75t_L g3062 ( 
.A1(n_2839),
.A2(n_2026),
.B1(n_2028),
.B2(n_1951),
.Y(n_3062)
);

INVx2_ASAP7_75t_SL g3063 ( 
.A(n_2769),
.Y(n_3063)
);

AND3x2_ASAP7_75t_L g3064 ( 
.A(n_2824),
.B(n_1471),
.C(n_1470),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2607),
.Y(n_3065)
);

INVx3_ASAP7_75t_L g3066 ( 
.A(n_2725),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2622),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2763),
.B(n_1489),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2659),
.Y(n_3069)
);

INVx2_ASAP7_75t_SL g3070 ( 
.A(n_2884),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2660),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2669),
.Y(n_3072)
);

OAI22xp5_ASAP7_75t_L g3073 ( 
.A1(n_2765),
.A2(n_1456),
.B1(n_1463),
.B2(n_1453),
.Y(n_3073)
);

CKINVDCx5p33_ASAP7_75t_R g3074 ( 
.A(n_2613),
.Y(n_3074)
);

AOI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2785),
.A2(n_1476),
.B1(n_1480),
.B2(n_1469),
.Y(n_3075)
);

BUFx3_ASAP7_75t_L g3076 ( 
.A(n_2605),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2671),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_SL g3078 ( 
.A1(n_2751),
.A2(n_2069),
.B1(n_1576),
.B2(n_1818),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2682),
.Y(n_3079)
);

INVx1_ASAP7_75t_SL g3080 ( 
.A(n_2881),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2717),
.B(n_1307),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2638),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2874),
.B(n_1512),
.Y(n_3083)
);

BUFx10_ASAP7_75t_L g3084 ( 
.A(n_2698),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2656),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2800),
.B(n_1525),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_SL g3087 ( 
.A(n_2768),
.B(n_1491),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2800),
.B(n_2895),
.Y(n_3088)
);

OAI22xp33_ASAP7_75t_L g3089 ( 
.A1(n_2854),
.A2(n_1528),
.B1(n_1538),
.B2(n_1527),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2680),
.Y(n_3090)
);

OAI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2829),
.A2(n_2831),
.B1(n_2640),
.B2(n_2727),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2684),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2685),
.Y(n_3093)
);

NAND3xp33_ASAP7_75t_L g3094 ( 
.A(n_2842),
.B(n_1314),
.C(n_1312),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2691),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2725),
.Y(n_3096)
);

INVx3_ASAP7_75t_L g3097 ( 
.A(n_2737),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2681),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2800),
.B(n_1578),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2692),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_SL g3101 ( 
.A(n_2587),
.B(n_1493),
.Y(n_3101)
);

BUFx6f_ASAP7_75t_SL g3102 ( 
.A(n_2634),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2693),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_SL g3104 ( 
.A(n_2877),
.B(n_1502),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2701),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2702),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2704),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2873),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2694),
.A2(n_1590),
.B1(n_1621),
.B2(n_1601),
.Y(n_3109)
);

INVx8_ASAP7_75t_L g3110 ( 
.A(n_2584),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2849),
.Y(n_3111)
);

INVx8_ASAP7_75t_L g3112 ( 
.A(n_2588),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2887),
.B(n_1505),
.Y(n_3113)
);

INVx3_ASAP7_75t_L g3114 ( 
.A(n_2737),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_2616),
.Y(n_3115)
);

BUFx10_ASAP7_75t_L g3116 ( 
.A(n_2710),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2600),
.Y(n_3117)
);

NOR2xp33_ASAP7_75t_SL g3118 ( 
.A(n_2619),
.B(n_1576),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2601),
.Y(n_3119)
);

BUFx3_ASAP7_75t_L g3120 ( 
.A(n_2598),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2615),
.Y(n_3121)
);

NAND2xp33_ASAP7_75t_SL g3122 ( 
.A(n_2733),
.B(n_1315),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_2617),
.Y(n_3123)
);

CKINVDCx5p33_ASAP7_75t_R g3124 ( 
.A(n_2649),
.Y(n_3124)
);

BUFx3_ASAP7_75t_L g3125 ( 
.A(n_2815),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2735),
.B(n_1631),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2893),
.B(n_1643),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2703),
.Y(n_3128)
);

INVx3_ASAP7_75t_L g3129 ( 
.A(n_2749),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2620),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2749),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2623),
.Y(n_3132)
);

CKINVDCx5p33_ASAP7_75t_R g3133 ( 
.A(n_2658),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2764),
.B(n_1653),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2625),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2628),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2741),
.B(n_2632),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2633),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2916),
.B(n_2662),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_3025),
.B(n_2739),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2958),
.B(n_2629),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2897),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2899),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2900),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2927),
.B(n_2729),
.Y(n_3145)
);

AOI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_3021),
.A2(n_2655),
.B1(n_2723),
.B2(n_2744),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_3070),
.B(n_2888),
.Y(n_3147)
);

BUFx3_ASAP7_75t_L g3148 ( 
.A(n_2972),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2905),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2906),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2977),
.B(n_2851),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2957),
.B(n_2955),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2910),
.B(n_2892),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_3127),
.B(n_2740),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2951),
.B(n_2956),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_3108),
.B(n_2858),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2924),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_2974),
.B(n_2779),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2909),
.Y(n_3159)
);

BUFx2_ASAP7_75t_R g3160 ( 
.A(n_3124),
.Y(n_3160)
);

NOR2xp33_ASAP7_75t_L g3161 ( 
.A(n_2976),
.B(n_2810),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2911),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2932),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2943),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2913),
.Y(n_3165)
);

INVx2_ASAP7_75t_SL g3166 ( 
.A(n_3026),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_3002),
.Y(n_3167)
);

INVx1_ASAP7_75t_SL g3168 ( 
.A(n_3007),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2915),
.Y(n_3169)
);

NOR2xp67_ASAP7_75t_L g3170 ( 
.A(n_3133),
.B(n_2627),
.Y(n_3170)
);

OR2x2_ASAP7_75t_L g3171 ( 
.A(n_2935),
.B(n_2867),
.Y(n_3171)
);

NAND2xp33_ASAP7_75t_L g3172 ( 
.A(n_3088),
.B(n_2716),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_3010),
.B(n_2614),
.Y(n_3173)
);

A2O1A1Ixp33_ASAP7_75t_L g3174 ( 
.A1(n_2940),
.A2(n_2714),
.B(n_2823),
.C(n_2646),
.Y(n_3174)
);

BUFx5_ASAP7_75t_L g3175 ( 
.A(n_2944),
.Y(n_3175)
);

NAND3xp33_ASAP7_75t_L g3176 ( 
.A(n_3078),
.B(n_3094),
.C(n_2914),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2904),
.B(n_2721),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_3091),
.B(n_2679),
.Y(n_3178)
);

INVxp67_ASAP7_75t_L g3179 ( 
.A(n_2920),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2952),
.B(n_2799),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2961),
.Y(n_3181)
);

XOR2x2_ASAP7_75t_L g3182 ( 
.A(n_3081),
.B(n_2788),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2963),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_3113),
.B(n_3104),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2982),
.B(n_3000),
.Y(n_3185)
);

BUFx3_ASAP7_75t_L g3186 ( 
.A(n_2972),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2979),
.B(n_1657),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_3006),
.B(n_2689),
.Y(n_3188)
);

AOI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_2969),
.A2(n_2825),
.B1(n_2891),
.B2(n_2827),
.Y(n_3189)
);

NOR3xp33_ASAP7_75t_L g3190 ( 
.A(n_2950),
.B(n_2776),
.C(n_2758),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_3053),
.B(n_2989),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2948),
.B(n_2697),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_3052),
.B(n_2706),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2918),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2992),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_2898),
.B(n_2815),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2994),
.B(n_1658),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2997),
.B(n_1671),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_SL g3199 ( 
.A(n_3005),
.B(n_2819),
.Y(n_3199)
);

INVx2_ASAP7_75t_SL g3200 ( 
.A(n_3026),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3017),
.B(n_1672),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3022),
.B(n_1688),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_3024),
.B(n_1692),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2925),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3055),
.B(n_1701),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_3027),
.B(n_1707),
.Y(n_3206)
);

INVx1_ASAP7_75t_SL g3207 ( 
.A(n_2988),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3028),
.Y(n_3208)
);

NAND3xp33_ASAP7_75t_L g3209 ( 
.A(n_3118),
.B(n_2730),
.C(n_2726),
.Y(n_3209)
);

BUFx3_ASAP7_75t_L g3210 ( 
.A(n_2993),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3030),
.Y(n_3211)
);

INVxp67_ASAP7_75t_L g3212 ( 
.A(n_2949),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_3033),
.B(n_2819),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2930),
.B(n_1742),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2931),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2934),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2936),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2901),
.B(n_1757),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2939),
.Y(n_3219)
);

OAI22xp33_ASAP7_75t_L g3220 ( 
.A1(n_3016),
.A2(n_2761),
.B1(n_2674),
.B2(n_2666),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_3083),
.A2(n_2855),
.B(n_2886),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3001),
.B(n_2708),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2907),
.B(n_2709),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_3069),
.B(n_2853),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2945),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_2993),
.Y(n_3226)
);

XNOR2xp5_ASAP7_75t_L g3227 ( 
.A(n_2937),
.B(n_2624),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2946),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_2947),
.B(n_1766),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3045),
.B(n_1778),
.Y(n_3230)
);

NOR3xp33_ASAP7_75t_L g3231 ( 
.A(n_2926),
.B(n_2637),
.C(n_2635),
.Y(n_3231)
);

NOR2xp33_ASAP7_75t_L g3232 ( 
.A(n_2941),
.B(n_2670),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2964),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2965),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_3039),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2966),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2975),
.B(n_1791),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2978),
.B(n_1806),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2980),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_3071),
.B(n_2853),
.Y(n_3240)
);

NAND2xp33_ASAP7_75t_SL g3241 ( 
.A(n_2970),
.B(n_2828),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2984),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_3072),
.B(n_2631),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2986),
.B(n_1832),
.Y(n_3244)
);

NAND3xp33_ASAP7_75t_L g3245 ( 
.A(n_2968),
.B(n_2742),
.C(n_2738),
.Y(n_3245)
);

AOI22xp5_ASAP7_75t_L g3246 ( 
.A1(n_3077),
.A2(n_1895),
.B1(n_1897),
.B2(n_1849),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2987),
.B(n_1904),
.Y(n_3247)
);

NOR3xp33_ASAP7_75t_L g3248 ( 
.A(n_2919),
.B(n_2643),
.C(n_2642),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2991),
.B(n_2995),
.Y(n_3249)
);

NOR2xp33_ASAP7_75t_L g3250 ( 
.A(n_3074),
.B(n_2748),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2996),
.B(n_1914),
.Y(n_3251)
);

AO221x1_ASAP7_75t_L g3252 ( 
.A1(n_3089),
.A2(n_2755),
.B1(n_2663),
.B2(n_1551),
.C(n_1561),
.Y(n_3252)
);

NAND2x1_ASAP7_75t_L g3253 ( 
.A(n_3037),
.B(n_2835),
.Y(n_3253)
);

BUFx5_ASAP7_75t_L g3254 ( 
.A(n_3040),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3009),
.B(n_1921),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_3115),
.B(n_3123),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3038),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_2953),
.Y(n_3258)
);

INVxp67_ASAP7_75t_L g3259 ( 
.A(n_3015),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_3068),
.B(n_2755),
.Y(n_3260)
);

XOR2xp5_ASAP7_75t_L g3261 ( 
.A(n_2999),
.B(n_2636),
.Y(n_3261)
);

OR2x2_ASAP7_75t_L g3262 ( 
.A(n_3080),
.B(n_2715),
.Y(n_3262)
);

AO221x1_ASAP7_75t_L g3263 ( 
.A1(n_3062),
.A2(n_1569),
.B1(n_1579),
.B2(n_1542),
.C(n_1534),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_3023),
.B(n_1958),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2954),
.B(n_2960),
.Y(n_3265)
);

NOR3xp33_ASAP7_75t_L g3266 ( 
.A(n_3087),
.B(n_2844),
.C(n_2801),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2962),
.B(n_2011),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2998),
.B(n_2022),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3004),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3137),
.B(n_2736),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3013),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_2908),
.B(n_2754),
.Y(n_3272)
);

AO221x1_ASAP7_75t_L g3273 ( 
.A1(n_3011),
.A2(n_1607),
.B1(n_1614),
.B2(n_1597),
.C(n_1585),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_2928),
.A2(n_2766),
.B(n_2865),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3014),
.B(n_3035),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_3079),
.B(n_2639),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_3046),
.B(n_3047),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_3049),
.B(n_2029),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3134),
.B(n_2040),
.Y(n_3279)
);

NOR2xp33_ASAP7_75t_L g3280 ( 
.A(n_3092),
.B(n_2833),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3093),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3095),
.B(n_3100),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_SL g3283 ( 
.A(n_3105),
.B(n_2641),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3107),
.B(n_2042),
.Y(n_3284)
);

NOR2xp33_ASAP7_75t_L g3285 ( 
.A(n_2912),
.B(n_2648),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_3051),
.B(n_2771),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3109),
.B(n_2050),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3041),
.B(n_2883),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_3042),
.B(n_1511),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_3044),
.B(n_2796),
.Y(n_3290)
);

BUFx5_ASAP7_75t_L g3291 ( 
.A(n_3054),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2921),
.B(n_2064),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_3058),
.B(n_1515),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2921),
.B(n_1522),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2921),
.B(n_1529),
.Y(n_3295)
);

INVxp33_ASAP7_75t_L g3296 ( 
.A(n_3015),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3117),
.Y(n_3297)
);

AO22x2_ASAP7_75t_L g3298 ( 
.A1(n_3176),
.A2(n_3120),
.B1(n_1626),
.B2(n_1656),
.Y(n_3298)
);

NAND2xp33_ASAP7_75t_L g3299 ( 
.A(n_3175),
.B(n_2973),
.Y(n_3299)
);

INVx3_ASAP7_75t_R g3300 ( 
.A(n_3262),
.Y(n_3300)
);

CKINVDCx11_ASAP7_75t_R g3301 ( 
.A(n_3207),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3142),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_3226),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3144),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3143),
.Y(n_3305)
);

INVxp67_ASAP7_75t_SL g3306 ( 
.A(n_3167),
.Y(n_3306)
);

HB1xp67_ASAP7_75t_L g3307 ( 
.A(n_3226),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3149),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_3152),
.B(n_3076),
.Y(n_3309)
);

OAI21xp33_ASAP7_75t_L g3310 ( 
.A1(n_3145),
.A2(n_3126),
.B(n_3075),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3150),
.Y(n_3311)
);

NAND2x1p5_ASAP7_75t_L g3312 ( 
.A(n_3148),
.B(n_3039),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3159),
.Y(n_3313)
);

AO22x2_ASAP7_75t_L g3314 ( 
.A1(n_3178),
.A2(n_1670),
.B1(n_1674),
.B2(n_1620),
.Y(n_3314)
);

CKINVDCx5p33_ASAP7_75t_R g3315 ( 
.A(n_3160),
.Y(n_3315)
);

CKINVDCx20_ASAP7_75t_R g3316 ( 
.A(n_3227),
.Y(n_3316)
);

AOI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3151),
.A2(n_2973),
.B1(n_3056),
.B2(n_3012),
.Y(n_3317)
);

INVxp67_ASAP7_75t_L g3318 ( 
.A(n_3155),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3157),
.Y(n_3319)
);

OAI221xp5_ASAP7_75t_L g3320 ( 
.A1(n_3146),
.A2(n_3122),
.B1(n_3048),
.B2(n_3111),
.C(n_3050),
.Y(n_3320)
);

HB1xp67_ASAP7_75t_L g3321 ( 
.A(n_3186),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3163),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3191),
.B(n_2973),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3164),
.Y(n_3324)
);

NAND2x1p5_ASAP7_75t_L g3325 ( 
.A(n_3210),
.B(n_2923),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3154),
.B(n_3059),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3181),
.Y(n_3327)
);

OAI221xp5_ASAP7_75t_L g3328 ( 
.A1(n_3212),
.A2(n_3048),
.B1(n_3063),
.B2(n_3031),
.C(n_3101),
.Y(n_3328)
);

AO22x2_ASAP7_75t_L g3329 ( 
.A1(n_3171),
.A2(n_1695),
.B1(n_1696),
.B2(n_1693),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_SL g3330 ( 
.A1(n_3173),
.A2(n_3110),
.B1(n_3112),
.B2(n_3102),
.Y(n_3330)
);

AND2x4_ASAP7_75t_L g3331 ( 
.A(n_3270),
.B(n_2983),
.Y(n_3331)
);

AND2x4_ASAP7_75t_L g3332 ( 
.A(n_3288),
.B(n_3125),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3162),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3183),
.Y(n_3334)
);

AO22x2_ASAP7_75t_L g3335 ( 
.A1(n_3141),
.A2(n_1703),
.B1(n_1706),
.B2(n_1700),
.Y(n_3335)
);

AO22x2_ASAP7_75t_L g3336 ( 
.A1(n_3195),
.A2(n_1711),
.B1(n_1714),
.B2(n_1708),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3208),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3211),
.Y(n_3338)
);

AOI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3184),
.A2(n_2917),
.B1(n_3067),
.B2(n_3065),
.Y(n_3339)
);

AO22x2_ASAP7_75t_L g3340 ( 
.A1(n_3168),
.A2(n_3297),
.B1(n_3248),
.B2(n_3156),
.Y(n_3340)
);

CKINVDCx5p33_ASAP7_75t_R g3341 ( 
.A(n_3256),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3281),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3249),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3265),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3140),
.B(n_3061),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3275),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3233),
.Y(n_3347)
);

INVxp67_ASAP7_75t_L g3348 ( 
.A(n_3158),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3242),
.Y(n_3349)
);

BUFx3_ASAP7_75t_L g3350 ( 
.A(n_3166),
.Y(n_3350)
);

BUFx8_ASAP7_75t_L g3351 ( 
.A(n_3200),
.Y(n_3351)
);

BUFx6f_ASAP7_75t_L g3352 ( 
.A(n_3235),
.Y(n_3352)
);

NOR2xp67_ASAP7_75t_L g3353 ( 
.A(n_3209),
.B(n_2985),
.Y(n_3353)
);

AO22x2_ASAP7_75t_L g3354 ( 
.A1(n_3190),
.A2(n_3266),
.B1(n_3179),
.B2(n_3245),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3269),
.Y(n_3355)
);

NAND2x1p5_ASAP7_75t_L g3356 ( 
.A(n_3170),
.B(n_3036),
.Y(n_3356)
);

NAND2xp33_ASAP7_75t_L g3357 ( 
.A(n_3175),
.B(n_3018),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3271),
.Y(n_3358)
);

AOI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3185),
.A2(n_3085),
.B1(n_3090),
.B2(n_3082),
.Y(n_3359)
);

AND2x4_ASAP7_75t_L g3360 ( 
.A(n_3222),
.B(n_3043),
.Y(n_3360)
);

BUFx8_ASAP7_75t_L g3361 ( 
.A(n_3193),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3215),
.Y(n_3362)
);

AO22x2_ASAP7_75t_L g3363 ( 
.A1(n_3147),
.A2(n_1730),
.B1(n_1738),
.B2(n_1725),
.Y(n_3363)
);

AO22x2_ASAP7_75t_L g3364 ( 
.A1(n_3292),
.A2(n_1747),
.B1(n_1748),
.B2(n_1746),
.Y(n_3364)
);

AO22x2_ASAP7_75t_L g3365 ( 
.A1(n_3218),
.A2(n_1755),
.B1(n_1758),
.B2(n_1750),
.Y(n_3365)
);

CKINVDCx5p33_ASAP7_75t_R g3366 ( 
.A(n_3250),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3139),
.B(n_3034),
.Y(n_3367)
);

NAND2x1p5_ASAP7_75t_L g3368 ( 
.A(n_3153),
.B(n_3018),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3225),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_3192),
.B(n_3110),
.Y(n_3370)
);

AOI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_3290),
.A2(n_3103),
.B1(n_3106),
.B2(n_3098),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3165),
.Y(n_3372)
);

OR2x2_ASAP7_75t_L g3373 ( 
.A(n_3205),
.B(n_3112),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3169),
.Y(n_3374)
);

CKINVDCx5p33_ASAP7_75t_R g3375 ( 
.A(n_3223),
.Y(n_3375)
);

CKINVDCx5p33_ASAP7_75t_R g3376 ( 
.A(n_3232),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_3259),
.B(n_2938),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3194),
.Y(n_3378)
);

AO22x2_ASAP7_75t_L g3379 ( 
.A1(n_3231),
.A2(n_1762),
.B1(n_1764),
.B2(n_1761),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3204),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3216),
.Y(n_3381)
);

AND2x4_ASAP7_75t_L g3382 ( 
.A(n_3213),
.B(n_2942),
.Y(n_3382)
);

NOR2xp67_ASAP7_75t_L g3383 ( 
.A(n_3285),
.B(n_3286),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3217),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_3175),
.B(n_3029),
.Y(n_3385)
);

AOI22xp5_ASAP7_75t_L g3386 ( 
.A1(n_3180),
.A2(n_3128),
.B1(n_3121),
.B2(n_3119),
.Y(n_3386)
);

A2O1A1Ixp33_ASAP7_75t_L g3387 ( 
.A1(n_3161),
.A2(n_3073),
.B(n_3099),
.C(n_3086),
.Y(n_3387)
);

AO22x2_ASAP7_75t_L g3388 ( 
.A1(n_3252),
.A2(n_3282),
.B1(n_3243),
.B2(n_3276),
.Y(n_3388)
);

AO22x2_ASAP7_75t_L g3389 ( 
.A1(n_3283),
.A2(n_1782),
.B1(n_1797),
.B2(n_1780),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3219),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3228),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3257),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3277),
.Y(n_3393)
);

NAND2x1p5_ASAP7_75t_L g3394 ( 
.A(n_3177),
.B(n_3029),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3175),
.B(n_3064),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3254),
.B(n_3130),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3254),
.B(n_3132),
.Y(n_3397)
);

OR2x6_ASAP7_75t_L g3398 ( 
.A(n_3253),
.B(n_3096),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3234),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3236),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3230),
.A2(n_3136),
.B1(n_3138),
.B2(n_3135),
.Y(n_3401)
);

CKINVDCx20_ASAP7_75t_R g3402 ( 
.A(n_3241),
.Y(n_3402)
);

AO22x2_ASAP7_75t_L g3403 ( 
.A1(n_3261),
.A2(n_1807),
.B1(n_1816),
.B2(n_1803),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3239),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3258),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3254),
.B(n_2959),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_3188),
.B(n_3034),
.Y(n_3407)
);

AO22x2_ASAP7_75t_L g3408 ( 
.A1(n_3182),
.A2(n_1841),
.B1(n_1860),
.B2(n_1831),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3254),
.B(n_2981),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3291),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3291),
.B(n_2990),
.Y(n_3411)
);

AND2x4_ASAP7_75t_L g3412 ( 
.A(n_3224),
.B(n_3003),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3291),
.B(n_3008),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3214),
.Y(n_3414)
);

CKINVDCx16_ASAP7_75t_R g3415 ( 
.A(n_3189),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3229),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3197),
.Y(n_3417)
);

NOR2xp33_ASAP7_75t_L g3418 ( 
.A(n_3296),
.B(n_3096),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3291),
.Y(n_3419)
);

AO22x2_ASAP7_75t_L g3420 ( 
.A1(n_3199),
.A2(n_1880),
.B1(n_1881),
.B2(n_1875),
.Y(n_3420)
);

INVx4_ASAP7_75t_L g3421 ( 
.A(n_3220),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3198),
.Y(n_3422)
);

AO22x2_ASAP7_75t_L g3423 ( 
.A1(n_3240),
.A2(n_3196),
.B1(n_3263),
.B2(n_1892),
.Y(n_3423)
);

AND2x2_ASAP7_75t_SL g3424 ( 
.A(n_3172),
.B(n_3131),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3280),
.B(n_2902),
.Y(n_3425)
);

AO22x2_ASAP7_75t_L g3426 ( 
.A1(n_3273),
.A2(n_1894),
.B1(n_1905),
.B2(n_1886),
.Y(n_3426)
);

INVx3_ASAP7_75t_L g3427 ( 
.A(n_3294),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3201),
.Y(n_3428)
);

BUFx2_ASAP7_75t_L g3429 ( 
.A(n_3202),
.Y(n_3429)
);

AND2x4_ASAP7_75t_L g3430 ( 
.A(n_3260),
.B(n_3032),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3393),
.B(n_3203),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_3348),
.B(n_3272),
.Y(n_3432)
);

OAI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3417),
.A2(n_3428),
.B(n_3422),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3299),
.A2(n_3174),
.B(n_3221),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3302),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3309),
.B(n_2903),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_3318),
.B(n_3341),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_R g3438 ( 
.A(n_3366),
.B(n_2713),
.Y(n_3438)
);

AOI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3357),
.A2(n_3187),
.B(n_3279),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_3301),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3343),
.B(n_3206),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3344),
.B(n_3284),
.Y(n_3442)
);

OAI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3387),
.A2(n_3264),
.B(n_3255),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3346),
.B(n_3278),
.Y(n_3444)
);

A2O1A1Ixp33_ASAP7_75t_L g3445 ( 
.A1(n_3310),
.A2(n_3287),
.B(n_3274),
.C(n_3295),
.Y(n_3445)
);

AND2x2_ASAP7_75t_L g3446 ( 
.A(n_3345),
.B(n_3060),
.Y(n_3446)
);

INVx1_ASAP7_75t_SL g3447 ( 
.A(n_3331),
.Y(n_3447)
);

INVx8_ASAP7_75t_L g3448 ( 
.A(n_3332),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_3305),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3323),
.A2(n_3289),
.B(n_3238),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3308),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_3383),
.B(n_3375),
.Y(n_3452)
);

CKINVDCx5p33_ASAP7_75t_R g3453 ( 
.A(n_3376),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3414),
.A2(n_3244),
.B(n_3237),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3326),
.B(n_3247),
.Y(n_3455)
);

A2O1A1Ixp33_ASAP7_75t_L g3456 ( 
.A1(n_3317),
.A2(n_3251),
.B(n_3268),
.C(n_3267),
.Y(n_3456)
);

AOI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3416),
.A2(n_3293),
.B(n_2870),
.Y(n_3457)
);

O2A1O1Ixp5_ASAP7_75t_L g3458 ( 
.A1(n_3385),
.A2(n_3057),
.B(n_3097),
.C(n_3066),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_L g3459 ( 
.A(n_3421),
.B(n_2933),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3396),
.A2(n_3246),
.B(n_1715),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3360),
.B(n_3114),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3319),
.Y(n_3462)
);

AOI21x1_ASAP7_75t_L g3463 ( 
.A1(n_3397),
.A2(n_2528),
.B(n_2520),
.Y(n_3463)
);

INVx2_ASAP7_75t_SL g3464 ( 
.A(n_3361),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3406),
.A2(n_1715),
.B(n_1616),
.Y(n_3465)
);

AOI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_3407),
.A2(n_2806),
.B1(n_3020),
.B2(n_2967),
.Y(n_3466)
);

INVx3_ASAP7_75t_L g3467 ( 
.A(n_3352),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3322),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3429),
.B(n_2971),
.Y(n_3469)
);

OAI321xp33_ASAP7_75t_L g3470 ( 
.A1(n_3320),
.A2(n_1940),
.A3(n_1926),
.B1(n_1945),
.B2(n_1938),
.C(n_1915),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3409),
.A2(n_1715),
.B(n_1616),
.Y(n_3471)
);

OAI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3386),
.A2(n_1547),
.B(n_1540),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3314),
.B(n_3129),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3427),
.A2(n_1759),
.B(n_1616),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3411),
.A2(n_1844),
.B(n_1759),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3324),
.Y(n_3476)
);

NAND2x1p5_ASAP7_75t_L g3477 ( 
.A(n_3303),
.B(n_3131),
.Y(n_3477)
);

INVx1_ASAP7_75t_SL g3478 ( 
.A(n_3321),
.Y(n_3478)
);

BUFx6f_ASAP7_75t_L g3479 ( 
.A(n_3352),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3327),
.B(n_2529),
.Y(n_3480)
);

INVx3_ASAP7_75t_L g3481 ( 
.A(n_3350),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3334),
.B(n_3337),
.Y(n_3482)
);

NAND2x1p5_ASAP7_75t_L g3483 ( 
.A(n_3430),
.B(n_2922),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3338),
.Y(n_3484)
);

OAI21xp33_ASAP7_75t_L g3485 ( 
.A1(n_3329),
.A2(n_3020),
.B(n_2757),
.Y(n_3485)
);

INVxp67_ASAP7_75t_L g3486 ( 
.A(n_3306),
.Y(n_3486)
);

BUFx3_ASAP7_75t_L g3487 ( 
.A(n_3351),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3347),
.Y(n_3488)
);

OAI21xp33_ASAP7_75t_L g3489 ( 
.A1(n_3363),
.A2(n_1320),
.B(n_1318),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3413),
.A2(n_1844),
.B(n_1759),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3298),
.A2(n_1818),
.B1(n_1591),
.B2(n_1604),
.Y(n_3491)
);

O2A1O1Ixp33_ASAP7_75t_L g3492 ( 
.A1(n_3328),
.A2(n_1966),
.B(n_1981),
.C(n_1961),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3342),
.B(n_2542),
.Y(n_3493)
);

INVx1_ASAP7_75t_SL g3494 ( 
.A(n_3307),
.Y(n_3494)
);

CKINVDCx5p33_ASAP7_75t_R g3495 ( 
.A(n_3315),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3349),
.B(n_2552),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3410),
.A2(n_1980),
.B(n_1844),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3419),
.A2(n_1980),
.B(n_1552),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3355),
.Y(n_3499)
);

NAND3xp33_ASAP7_75t_L g3500 ( 
.A(n_3425),
.B(n_2845),
.C(n_2590),
.Y(n_3500)
);

INVx3_ASAP7_75t_L g3501 ( 
.A(n_3312),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3358),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3373),
.A2(n_1980),
.B(n_1553),
.Y(n_3503)
);

HB1xp67_ASAP7_75t_L g3504 ( 
.A(n_3300),
.Y(n_3504)
);

INVx3_ASAP7_75t_L g3505 ( 
.A(n_3325),
.Y(n_3505)
);

OAI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3399),
.A2(n_3405),
.B(n_3404),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3362),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3340),
.A2(n_1591),
.B1(n_1604),
.B2(n_1543),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3339),
.A2(n_1556),
.B(n_1549),
.Y(n_3509)
);

BUFx4f_ASAP7_75t_L g3510 ( 
.A(n_3356),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3388),
.B(n_2553),
.Y(n_3511)
);

BUFx8_ASAP7_75t_L g3512 ( 
.A(n_3367),
.Y(n_3512)
);

AOI22xp5_ASAP7_75t_L g3513 ( 
.A1(n_3370),
.A2(n_3116),
.B1(n_3084),
.B2(n_3019),
.Y(n_3513)
);

O2A1O1Ixp33_ASAP7_75t_L g3514 ( 
.A1(n_3395),
.A2(n_1990),
.B(n_1997),
.C(n_1989),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_3424),
.A2(n_3401),
.B(n_3369),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3400),
.A2(n_1580),
.B(n_1557),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3304),
.A2(n_1588),
.B(n_1582),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3372),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3311),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3374),
.B(n_2574),
.Y(n_3520)
);

BUFx6f_ASAP7_75t_L g3521 ( 
.A(n_3377),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3378),
.B(n_2575),
.Y(n_3522)
);

AOI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_3313),
.A2(n_1599),
.B(n_1589),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3333),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3380),
.B(n_2580),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3391),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3381),
.A2(n_1615),
.B(n_1610),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3384),
.B(n_2929),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_L g3529 ( 
.A(n_3415),
.B(n_2882),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3390),
.B(n_1617),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3392),
.A2(n_1624),
.B(n_1623),
.Y(n_3531)
);

BUFx6f_ASAP7_75t_L g3532 ( 
.A(n_3418),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3359),
.A2(n_1645),
.B(n_1634),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3335),
.B(n_1652),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3371),
.A2(n_1661),
.B(n_1655),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3420),
.B(n_1663),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_3330),
.B(n_1912),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3364),
.B(n_1912),
.Y(n_3538)
);

AO21x2_ASAP7_75t_L g3539 ( 
.A1(n_3434),
.A2(n_3353),
.B(n_3412),
.Y(n_3539)
);

CKINVDCx5p33_ASAP7_75t_R g3540 ( 
.A(n_3453),
.Y(n_3540)
);

OAI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3432),
.A2(n_3368),
.B1(n_3394),
.B2(n_3402),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3435),
.Y(n_3542)
);

A2O1A1Ixp33_ASAP7_75t_L g3543 ( 
.A1(n_3470),
.A2(n_3382),
.B(n_3379),
.C(n_3389),
.Y(n_3543)
);

BUFx3_ASAP7_75t_L g3544 ( 
.A(n_3479),
.Y(n_3544)
);

HB1xp67_ASAP7_75t_L g3545 ( 
.A(n_3478),
.Y(n_3545)
);

OR2x2_ASAP7_75t_L g3546 ( 
.A(n_3433),
.B(n_3398),
.Y(n_3546)
);

O2A1O1Ixp33_ASAP7_75t_L g3547 ( 
.A1(n_3492),
.A2(n_2014),
.B(n_2017),
.C(n_2004),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3449),
.Y(n_3548)
);

O2A1O1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_3537),
.A2(n_2023),
.B(n_2037),
.C(n_2020),
.Y(n_3549)
);

OAI21xp33_ASAP7_75t_L g3550 ( 
.A1(n_3489),
.A2(n_3365),
.B(n_3408),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3482),
.Y(n_3551)
);

INVx4_ASAP7_75t_L g3552 ( 
.A(n_3479),
.Y(n_3552)
);

O2A1O1Ixp33_ASAP7_75t_L g3553 ( 
.A1(n_3534),
.A2(n_2048),
.B(n_2053),
.C(n_2047),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3437),
.B(n_3452),
.Y(n_3554)
);

AND2x4_ASAP7_75t_L g3555 ( 
.A(n_3467),
.B(n_3316),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3443),
.A2(n_3456),
.B(n_3445),
.Y(n_3556)
);

AOI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_3439),
.A2(n_3354),
.B(n_3423),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3451),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_R g3559 ( 
.A(n_3495),
.B(n_2861),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3446),
.B(n_3426),
.Y(n_3560)
);

OAI21xp33_ASAP7_75t_SL g3561 ( 
.A1(n_3455),
.A2(n_2056),
.B(n_1594),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3462),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3519),
.B(n_3336),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3431),
.B(n_3403),
.Y(n_3564)
);

OAI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3466),
.A2(n_1323),
.B1(n_1330),
.B2(n_1321),
.Y(n_3565)
);

AOI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3463),
.A2(n_1619),
.B(n_1573),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_3532),
.B(n_2889),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_3459),
.B(n_1664),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3454),
.A2(n_1668),
.B(n_1665),
.Y(n_3569)
);

NAND2x1p5_ASAP7_75t_L g3570 ( 
.A(n_3510),
.B(n_1633),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3441),
.B(n_1331),
.Y(n_3571)
);

O2A1O1Ixp33_ASAP7_75t_L g3572 ( 
.A1(n_3514),
.A2(n_1756),
.B(n_1765),
.C(n_1650),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3442),
.B(n_1334),
.Y(n_3573)
);

BUFx2_ASAP7_75t_L g3574 ( 
.A(n_3532),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3488),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3444),
.B(n_1340),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3468),
.Y(n_3577)
);

AOI21xp5_ASAP7_75t_L g3578 ( 
.A1(n_3450),
.A2(n_1673),
.B(n_1669),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3436),
.B(n_1343),
.Y(n_3579)
);

NOR3xp33_ASAP7_75t_SL g3580 ( 
.A(n_3500),
.B(n_1352),
.C(n_1346),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3499),
.Y(n_3581)
);

A2O1A1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_3515),
.A2(n_1825),
.B(n_1877),
.C(n_1821),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_SL g3583 ( 
.A(n_3485),
.B(n_3469),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_3472),
.A2(n_1963),
.B1(n_2036),
.B2(n_1929),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3447),
.B(n_1353),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3486),
.B(n_1361),
.Y(n_3586)
);

O2A1O1Ixp33_ASAP7_75t_L g3587 ( 
.A1(n_3536),
.A2(n_1941),
.B(n_1971),
.C(n_1949),
.Y(n_3587)
);

OAI21xp33_ASAP7_75t_L g3588 ( 
.A1(n_3491),
.A2(n_1367),
.B(n_1362),
.Y(n_3588)
);

AOI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_3529),
.A2(n_1689),
.B1(n_1690),
.B2(n_1685),
.Y(n_3589)
);

NOR2xp33_ASAP7_75t_L g3590 ( 
.A(n_3494),
.B(n_1698),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3524),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3526),
.B(n_3506),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3448),
.B(n_1369),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_SL g3594 ( 
.A(n_3513),
.B(n_3473),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3460),
.A2(n_1721),
.B(n_1712),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3521),
.Y(n_3596)
);

NAND2x1p5_ASAP7_75t_L g3597 ( 
.A(n_3481),
.B(n_2067),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_3457),
.A2(n_1732),
.B(n_1722),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3476),
.Y(n_3599)
);

O2A1O1Ixp33_ASAP7_75t_L g3600 ( 
.A1(n_3511),
.A2(n_3538),
.B(n_3504),
.C(n_3503),
.Y(n_3600)
);

INVx1_ASAP7_75t_SL g3601 ( 
.A(n_3448),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3484),
.B(n_1374),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3461),
.B(n_1379),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3502),
.Y(n_3604)
);

INVx3_ASAP7_75t_L g3605 ( 
.A(n_3521),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3507),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_3498),
.A2(n_1745),
.B(n_1737),
.Y(n_3607)
);

A2O1A1Ixp33_ASAP7_75t_L g3608 ( 
.A1(n_3509),
.A2(n_1752),
.B(n_1754),
.C(n_1751),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3518),
.B(n_1380),
.Y(n_3609)
);

CKINVDCx5p33_ASAP7_75t_R g3610 ( 
.A(n_3438),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3528),
.Y(n_3611)
);

BUFx8_ASAP7_75t_L g3612 ( 
.A(n_3487),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3474),
.A2(n_1774),
.B(n_1773),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_3477),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_SL g3615 ( 
.A(n_3530),
.B(n_1776),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3480),
.Y(n_3616)
);

INVxp33_ASAP7_75t_L g3617 ( 
.A(n_3483),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3512),
.B(n_3501),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_3505),
.B(n_1786),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3496),
.B(n_1381),
.Y(n_3620)
);

INVx4_ASAP7_75t_L g3621 ( 
.A(n_3464),
.Y(n_3621)
);

A2O1A1Ixp33_ASAP7_75t_L g3622 ( 
.A1(n_3535),
.A2(n_3533),
.B(n_3531),
.C(n_3527),
.Y(n_3622)
);

A2O1A1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_3516),
.A2(n_1802),
.B(n_1812),
.C(n_1789),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3440),
.B(n_3493),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3520),
.B(n_1813),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3522),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3525),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_SL g3628 ( 
.A(n_3517),
.B(n_1929),
.Y(n_3628)
);

INVx4_ASAP7_75t_L g3629 ( 
.A(n_3458),
.Y(n_3629)
);

OAI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_3508),
.A2(n_1385),
.B1(n_1387),
.B2(n_1383),
.Y(n_3630)
);

OAI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3523),
.A2(n_1389),
.B1(n_1393),
.B2(n_1388),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3465),
.A2(n_1828),
.B(n_1819),
.Y(n_3632)
);

O2A1O1Ixp5_ASAP7_75t_L g3633 ( 
.A1(n_3471),
.A2(n_1591),
.B(n_1604),
.C(n_1543),
.Y(n_3633)
);

INVx1_ASAP7_75t_SL g3634 ( 
.A(n_3475),
.Y(n_3634)
);

O2A1O1Ixp33_ASAP7_75t_L g3635 ( 
.A1(n_3490),
.A2(n_2036),
.B(n_1963),
.C(n_1395),
.Y(n_3635)
);

BUFx6f_ASAP7_75t_L g3636 ( 
.A(n_3497),
.Y(n_3636)
);

AND2x4_ASAP7_75t_L g3637 ( 
.A(n_3467),
.B(n_888),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3443),
.A2(n_1839),
.B(n_1837),
.Y(n_3638)
);

BUFx6f_ASAP7_75t_L g3639 ( 
.A(n_3479),
.Y(n_3639)
);

O2A1O1Ixp33_ASAP7_75t_L g3640 ( 
.A1(n_3470),
.A2(n_1396),
.B(n_1402),
.C(n_1394),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_3437),
.B(n_1848),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3431),
.B(n_1405),
.Y(n_3642)
);

INVxp67_ASAP7_75t_L g3643 ( 
.A(n_3437),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3443),
.A2(n_1854),
.B(n_1851),
.Y(n_3644)
);

A2O1A1Ixp33_ASAP7_75t_L g3645 ( 
.A1(n_3470),
.A2(n_1873),
.B(n_1874),
.C(n_1856),
.Y(n_3645)
);

CKINVDCx5p33_ASAP7_75t_R g3646 ( 
.A(n_3453),
.Y(n_3646)
);

AOI21x1_ASAP7_75t_L g3647 ( 
.A1(n_3566),
.A2(n_3557),
.B(n_3638),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_3643),
.B(n_3554),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3616),
.B(n_1409),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3556),
.A2(n_3633),
.B(n_3600),
.Y(n_3650)
);

AOI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_3622),
.A2(n_1887),
.B(n_1876),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3584),
.A2(n_1418),
.B1(n_1425),
.B2(n_1417),
.Y(n_3652)
);

AOI211x1_ASAP7_75t_L g3653 ( 
.A1(n_3550),
.A2(n_1430),
.B(n_1433),
.C(n_1427),
.Y(n_3653)
);

OAI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3578),
.A2(n_1591),
.B(n_1543),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3577),
.Y(n_3655)
);

OAI21x1_ASAP7_75t_L g3656 ( 
.A1(n_3599),
.A2(n_1604),
.B(n_1591),
.Y(n_3656)
);

INVx5_ASAP7_75t_L g3657 ( 
.A(n_3639),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3626),
.B(n_1440),
.Y(n_3658)
);

NOR4xp25_ASAP7_75t_L g3659 ( 
.A(n_3553),
.B(n_4),
.C(n_1),
.D(n_3),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3604),
.Y(n_3660)
);

NAND2x1p5_ASAP7_75t_L g3661 ( 
.A(n_3574),
.B(n_889),
.Y(n_3661)
);

OAI21x1_ASAP7_75t_L g3662 ( 
.A1(n_3606),
.A2(n_1691),
.B(n_1604),
.Y(n_3662)
);

OAI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_3644),
.A2(n_3561),
.B(n_3569),
.Y(n_3663)
);

AO21x1_ASAP7_75t_L g3664 ( 
.A1(n_3594),
.A2(n_1691),
.B(n_5),
.Y(n_3664)
);

AOI22xp5_ASAP7_75t_L g3665 ( 
.A1(n_3583),
.A2(n_1465),
.B1(n_1466),
.B2(n_1451),
.Y(n_3665)
);

NAND2x1_ASAP7_75t_L g3666 ( 
.A(n_3636),
.B(n_2847),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3539),
.A2(n_1907),
.B(n_1903),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3634),
.A2(n_1911),
.B(n_1908),
.Y(n_3668)
);

BUFx2_ASAP7_75t_L g3669 ( 
.A(n_3545),
.Y(n_3669)
);

OAI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3641),
.A2(n_2847),
.B(n_1919),
.Y(n_3670)
);

BUFx6f_ASAP7_75t_L g3671 ( 
.A(n_3639),
.Y(n_3671)
);

OR2x2_ASAP7_75t_L g3672 ( 
.A(n_3564),
.B(n_1913),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3629),
.A2(n_1927),
.B(n_1925),
.Y(n_3673)
);

AND2x6_ASAP7_75t_L g3674 ( 
.A(n_3560),
.B(n_3563),
.Y(n_3674)
);

OAI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3635),
.A2(n_2847),
.B(n_1932),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_3544),
.B(n_3605),
.Y(n_3676)
);

OAI21x1_ASAP7_75t_L g3677 ( 
.A1(n_3598),
.A2(n_1691),
.B(n_892),
.Y(n_3677)
);

OAI21xp5_ASAP7_75t_SL g3678 ( 
.A1(n_3565),
.A2(n_1474),
.B(n_1472),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3627),
.B(n_1479),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3542),
.Y(n_3680)
);

NAND3xp33_ASAP7_75t_L g3681 ( 
.A(n_3587),
.B(n_1486),
.C(n_1482),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3615),
.A2(n_1933),
.B(n_1928),
.Y(n_3682)
);

NOR2xp33_ASAP7_75t_L g3683 ( 
.A(n_3624),
.B(n_1934),
.Y(n_3683)
);

AO31x2_ASAP7_75t_L g3684 ( 
.A1(n_3582),
.A2(n_1691),
.A3(n_8),
.B(n_5),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3579),
.B(n_3540),
.Y(n_3685)
);

OAI21xp33_ASAP7_75t_L g3686 ( 
.A1(n_3628),
.A2(n_1490),
.B(n_1488),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3558),
.Y(n_3687)
);

AOI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3625),
.A2(n_1946),
.B(n_1936),
.Y(n_3688)
);

BUFx4_ASAP7_75t_SL g3689 ( 
.A(n_3646),
.Y(n_3689)
);

AO31x2_ASAP7_75t_L g3690 ( 
.A1(n_3543),
.A2(n_1691),
.A3(n_9),
.B(n_7),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_L g3691 ( 
.A(n_3610),
.B(n_1495),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3548),
.Y(n_3692)
);

NOR2xp33_ASAP7_75t_L g3693 ( 
.A(n_3541),
.B(n_1950),
.Y(n_3693)
);

AO32x2_ASAP7_75t_L g3694 ( 
.A1(n_3630),
.A2(n_1506),
.A3(n_1508),
.B1(n_1501),
.B2(n_1498),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3551),
.B(n_1513),
.Y(n_3695)
);

INVx1_ASAP7_75t_SL g3696 ( 
.A(n_3555),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3562),
.Y(n_3697)
);

NAND2xp33_ASAP7_75t_R g3698 ( 
.A(n_3559),
.B(n_3580),
.Y(n_3698)
);

AOI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_3592),
.A2(n_3636),
.B(n_3608),
.Y(n_3699)
);

AOI221x1_ASAP7_75t_L g3700 ( 
.A1(n_3588),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3546),
.A2(n_1988),
.B(n_1976),
.Y(n_3701)
);

AOI22x1_ASAP7_75t_SL g3702 ( 
.A1(n_3621),
.A2(n_1517),
.B1(n_1519),
.B2(n_1516),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3611),
.B(n_1521),
.Y(n_3703)
);

BUFx3_ASAP7_75t_L g3704 ( 
.A(n_3596),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3575),
.Y(n_3705)
);

NOR2xp67_ASAP7_75t_L g3706 ( 
.A(n_3586),
.B(n_890),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3581),
.B(n_1524),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3568),
.A2(n_1994),
.B(n_1992),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3591),
.B(n_1995),
.Y(n_3709)
);

AOI21x1_ASAP7_75t_L g3710 ( 
.A1(n_3595),
.A2(n_2002),
.B(n_1998),
.Y(n_3710)
);

OAI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3632),
.A2(n_894),
.B(n_893),
.Y(n_3711)
);

OAI21x1_ASAP7_75t_L g3712 ( 
.A1(n_3572),
.A2(n_896),
.B(n_895),
.Y(n_3712)
);

OAI21x1_ASAP7_75t_L g3713 ( 
.A1(n_3613),
.A2(n_902),
.B(n_897),
.Y(n_3713)
);

OAI21x1_ASAP7_75t_L g3714 ( 
.A1(n_3607),
.A2(n_904),
.B(n_903),
.Y(n_3714)
);

AO22x1_ASAP7_75t_L g3715 ( 
.A1(n_3612),
.A2(n_1532),
.B1(n_1533),
.B2(n_1531),
.Y(n_3715)
);

INVx5_ASAP7_75t_L g3716 ( 
.A(n_3596),
.Y(n_3716)
);

INVxp67_ASAP7_75t_SL g3717 ( 
.A(n_3614),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3602),
.Y(n_3718)
);

OAI21x1_ASAP7_75t_L g3719 ( 
.A1(n_3547),
.A2(n_906),
.B(n_905),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3623),
.A2(n_3573),
.B(n_3571),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3576),
.B(n_3642),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3552),
.B(n_909),
.Y(n_3722)
);

NAND3x1_ASAP7_75t_L g3723 ( 
.A(n_3618),
.B(n_11),
.C(n_12),
.Y(n_3723)
);

AND2x4_ASAP7_75t_L g3724 ( 
.A(n_3601),
.B(n_911),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_SL g3725 ( 
.A(n_3597),
.B(n_2054),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3620),
.A2(n_2007),
.B(n_2003),
.Y(n_3726)
);

O2A1O1Ixp5_ASAP7_75t_SL g3727 ( 
.A1(n_3631),
.A2(n_1536),
.B(n_1539),
.C(n_1535),
.Y(n_3727)
);

INVxp33_ASAP7_75t_SL g3728 ( 
.A(n_3567),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3619),
.A2(n_2010),
.B(n_2009),
.Y(n_3729)
);

OAI21xp5_ASAP7_75t_SL g3730 ( 
.A1(n_3640),
.A2(n_1545),
.B(n_1544),
.Y(n_3730)
);

AOI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3590),
.A2(n_1554),
.B1(n_1555),
.B2(n_1548),
.Y(n_3731)
);

OAI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3645),
.A2(n_2016),
.B(n_2012),
.Y(n_3732)
);

OAI22xp5_ASAP7_75t_SL g3733 ( 
.A1(n_3570),
.A2(n_1564),
.B1(n_1567),
.B2(n_1558),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3609),
.B(n_2045),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3549),
.A2(n_914),
.B(n_913),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3589),
.B(n_2058),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3585),
.B(n_2059),
.Y(n_3737)
);

INVx3_ASAP7_75t_L g3738 ( 
.A(n_3637),
.Y(n_3738)
);

A2O1A1Ixp33_ASAP7_75t_L g3739 ( 
.A1(n_3593),
.A2(n_1572),
.B(n_1629),
.C(n_1605),
.Y(n_3739)
);

OAI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3720),
.A2(n_3693),
.B(n_3727),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3650),
.A2(n_3603),
.B(n_918),
.Y(n_3741)
);

A2O1A1Ixp33_ASAP7_75t_L g3742 ( 
.A1(n_3686),
.A2(n_3617),
.B(n_1574),
.C(n_1583),
.Y(n_3742)
);

AOI22xp33_ASAP7_75t_SL g3743 ( 
.A1(n_3663),
.A2(n_1584),
.B1(n_1587),
.B2(n_1568),
.Y(n_3743)
);

OAI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3683),
.A2(n_1595),
.B1(n_1596),
.B2(n_1593),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3687),
.Y(n_3745)
);

OAI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3662),
.A2(n_920),
.B(n_917),
.Y(n_3746)
);

OR2x2_ASAP7_75t_L g3747 ( 
.A(n_3669),
.B(n_11),
.Y(n_3747)
);

OAI21x1_ASAP7_75t_L g3748 ( 
.A1(n_3647),
.A2(n_922),
.B(n_921),
.Y(n_3748)
);

AOI22xp5_ASAP7_75t_L g3749 ( 
.A1(n_3730),
.A2(n_1612),
.B1(n_1613),
.B2(n_1611),
.Y(n_3749)
);

OAI21x1_ASAP7_75t_L g3750 ( 
.A1(n_3656),
.A2(n_925),
.B(n_923),
.Y(n_3750)
);

OAI21x1_ASAP7_75t_L g3751 ( 
.A1(n_3654),
.A2(n_927),
.B(n_926),
.Y(n_3751)
);

OAI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3678),
.A2(n_1622),
.B1(n_1627),
.B2(n_1618),
.Y(n_3752)
);

NOR2x1_ASAP7_75t_R g3753 ( 
.A(n_3716),
.B(n_1628),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3677),
.A2(n_929),
.B(n_928),
.Y(n_3754)
);

AND2x4_ASAP7_75t_L g3755 ( 
.A(n_3717),
.B(n_930),
.Y(n_3755)
);

OAI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3651),
.A2(n_2033),
.B(n_2021),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3655),
.Y(n_3757)
);

INVx6_ASAP7_75t_L g3758 ( 
.A(n_3657),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3699),
.A2(n_2041),
.B(n_2034),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3660),
.Y(n_3760)
);

OAI21x1_ASAP7_75t_L g3761 ( 
.A1(n_3712),
.A2(n_932),
.B(n_931),
.Y(n_3761)
);

OAI21x1_ASAP7_75t_L g3762 ( 
.A1(n_3714),
.A2(n_934),
.B(n_933),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3711),
.A2(n_939),
.B(n_935),
.Y(n_3763)
);

BUFx2_ASAP7_75t_SL g3764 ( 
.A(n_3657),
.Y(n_3764)
);

AOI22xp33_ASAP7_75t_L g3765 ( 
.A1(n_3681),
.A2(n_1635),
.B1(n_1637),
.B2(n_1632),
.Y(n_3765)
);

O2A1O1Ixp33_ASAP7_75t_SL g3766 ( 
.A1(n_3725),
.A2(n_21),
.B(n_31),
.C(n_12),
.Y(n_3766)
);

OAI21x1_ASAP7_75t_L g3767 ( 
.A1(n_3713),
.A2(n_942),
.B(n_940),
.Y(n_3767)
);

AOI22xp33_ASAP7_75t_L g3768 ( 
.A1(n_3674),
.A2(n_1646),
.B1(n_1647),
.B2(n_1640),
.Y(n_3768)
);

OA21x2_ASAP7_75t_L g3769 ( 
.A1(n_3667),
.A2(n_3664),
.B(n_3700),
.Y(n_3769)
);

OAI21x1_ASAP7_75t_L g3770 ( 
.A1(n_3719),
.A2(n_946),
.B(n_943),
.Y(n_3770)
);

OA21x2_ASAP7_75t_L g3771 ( 
.A1(n_3673),
.A2(n_2068),
.B(n_2063),
.Y(n_3771)
);

INVx2_ASAP7_75t_L g3772 ( 
.A(n_3705),
.Y(n_3772)
);

HB1xp67_ASAP7_75t_L g3773 ( 
.A(n_3680),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3692),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3697),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3735),
.A2(n_949),
.B(n_948),
.Y(n_3776)
);

OA21x2_ASAP7_75t_L g3777 ( 
.A1(n_3701),
.A2(n_1649),
.B(n_1648),
.Y(n_3777)
);

OR2x6_ASAP7_75t_L g3778 ( 
.A(n_3661),
.B(n_951),
.Y(n_3778)
);

O2A1O1Ixp5_ASAP7_75t_SL g3779 ( 
.A1(n_3718),
.A2(n_1654),
.B(n_1660),
.C(n_1651),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3721),
.B(n_1662),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3684),
.Y(n_3781)
);

CKINVDCx20_ASAP7_75t_R g3782 ( 
.A(n_3696),
.Y(n_3782)
);

INVx3_ASAP7_75t_L g3783 ( 
.A(n_3671),
.Y(n_3783)
);

OAI21x1_ASAP7_75t_L g3784 ( 
.A1(n_3710),
.A2(n_954),
.B(n_952),
.Y(n_3784)
);

BUFx6f_ASAP7_75t_L g3785 ( 
.A(n_3671),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3690),
.Y(n_3786)
);

NOR2xp33_ASAP7_75t_L g3787 ( 
.A(n_3648),
.B(n_3728),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_SL g3788 ( 
.A1(n_3670),
.A2(n_1676),
.B(n_1675),
.Y(n_3788)
);

O2A1O1Ixp33_ASAP7_75t_SL g3789 ( 
.A1(n_3736),
.A2(n_25),
.B(n_34),
.C(n_13),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3674),
.B(n_14),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3690),
.Y(n_3791)
);

OA21x2_ASAP7_75t_L g3792 ( 
.A1(n_3668),
.A2(n_1680),
.B(n_1677),
.Y(n_3792)
);

AOI22xp33_ASAP7_75t_L g3793 ( 
.A1(n_3674),
.A2(n_1684),
.B1(n_1686),
.B2(n_1681),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3684),
.Y(n_3794)
);

OAI22xp5_ASAP7_75t_L g3795 ( 
.A1(n_3653),
.A2(n_1704),
.B1(n_1709),
.B2(n_1687),
.Y(n_3795)
);

CKINVDCx20_ASAP7_75t_R g3796 ( 
.A(n_3704),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3709),
.Y(n_3797)
);

INVx3_ASAP7_75t_L g3798 ( 
.A(n_3676),
.Y(n_3798)
);

BUFx12f_ASAP7_75t_L g3799 ( 
.A(n_3716),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3707),
.Y(n_3800)
);

OAI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3723),
.A2(n_1717),
.B1(n_1718),
.B2(n_1713),
.Y(n_3801)
);

BUFx3_ASAP7_75t_L g3802 ( 
.A(n_3738),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3679),
.Y(n_3803)
);

NAND3xp33_ASAP7_75t_L g3804 ( 
.A(n_3659),
.B(n_1720),
.C(n_1719),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3703),
.Y(n_3805)
);

AO21x2_ASAP7_75t_L g3806 ( 
.A1(n_3732),
.A2(n_1727),
.B(n_1723),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3666),
.A2(n_957),
.B(n_955),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3695),
.B(n_1734),
.Y(n_3808)
);

AOI21x1_ASAP7_75t_L g3809 ( 
.A1(n_3726),
.A2(n_1740),
.B(n_1736),
.Y(n_3809)
);

INVx1_ASAP7_75t_SL g3810 ( 
.A(n_3689),
.Y(n_3810)
);

BUFx3_ASAP7_75t_L g3811 ( 
.A(n_3685),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3672),
.B(n_15),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3722),
.Y(n_3813)
);

NOR2xp67_ASAP7_75t_L g3814 ( 
.A(n_3649),
.B(n_15),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3675),
.A2(n_3706),
.B1(n_3724),
.B2(n_3652),
.Y(n_3815)
);

INVx2_ASAP7_75t_SL g3816 ( 
.A(n_3758),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3745),
.Y(n_3817)
);

BUFx2_ASAP7_75t_R g3818 ( 
.A(n_3764),
.Y(n_3818)
);

CKINVDCx20_ASAP7_75t_R g3819 ( 
.A(n_3796),
.Y(n_3819)
);

CKINVDCx5p33_ASAP7_75t_R g3820 ( 
.A(n_3799),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3773),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_L g3822 ( 
.A1(n_3741),
.A2(n_3729),
.B(n_3682),
.Y(n_3822)
);

OAI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3740),
.A2(n_3708),
.B(n_3665),
.Y(n_3823)
);

CKINVDCx20_ASAP7_75t_R g3824 ( 
.A(n_3782),
.Y(n_3824)
);

HB1xp67_ASAP7_75t_L g3825 ( 
.A(n_3757),
.Y(n_3825)
);

AOI22xp33_ASAP7_75t_L g3826 ( 
.A1(n_3804),
.A2(n_3734),
.B1(n_3658),
.B2(n_3733),
.Y(n_3826)
);

BUFx2_ASAP7_75t_L g3827 ( 
.A(n_3802),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3760),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3772),
.Y(n_3829)
);

AO21x2_ASAP7_75t_L g3830 ( 
.A1(n_3786),
.A2(n_3688),
.B(n_3739),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3743),
.A2(n_3737),
.B1(n_3691),
.B2(n_1743),
.Y(n_3831)
);

INVx2_ASAP7_75t_SL g3832 ( 
.A(n_3798),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3811),
.B(n_3715),
.Y(n_3833)
);

INVxp33_ASAP7_75t_L g3834 ( 
.A(n_3787),
.Y(n_3834)
);

CKINVDCx20_ASAP7_75t_R g3835 ( 
.A(n_3810),
.Y(n_3835)
);

INVx6_ASAP7_75t_L g3836 ( 
.A(n_3785),
.Y(n_3836)
);

AND2x4_ASAP7_75t_L g3837 ( 
.A(n_3774),
.B(n_959),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3775),
.Y(n_3838)
);

BUFx4f_ASAP7_75t_SL g3839 ( 
.A(n_3785),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3781),
.Y(n_3840)
);

INVx3_ASAP7_75t_L g3841 ( 
.A(n_3783),
.Y(n_3841)
);

BUFx10_ASAP7_75t_L g3842 ( 
.A(n_3803),
.Y(n_3842)
);

OR2x6_ASAP7_75t_L g3843 ( 
.A(n_3778),
.B(n_3698),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3791),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3794),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3797),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3806),
.A2(n_1744),
.B1(n_1749),
.B2(n_1741),
.Y(n_3847)
);

AND2x4_ASAP7_75t_L g3848 ( 
.A(n_3813),
.B(n_960),
.Y(n_3848)
);

NAND2x1p5_ASAP7_75t_L g3849 ( 
.A(n_3755),
.B(n_3731),
.Y(n_3849)
);

AOI22xp33_ASAP7_75t_SL g3850 ( 
.A1(n_3769),
.A2(n_3790),
.B1(n_3777),
.B2(n_3801),
.Y(n_3850)
);

OA21x2_ASAP7_75t_L g3851 ( 
.A1(n_3748),
.A2(n_1763),
.B(n_1760),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_3792),
.A2(n_1768),
.B1(n_1770),
.B2(n_1767),
.Y(n_3852)
);

OR2x6_ASAP7_75t_L g3853 ( 
.A(n_3778),
.B(n_3702),
.Y(n_3853)
);

CKINVDCx6p67_ASAP7_75t_R g3854 ( 
.A(n_3747),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3800),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3805),
.B(n_1775),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3812),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3754),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3750),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3746),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3762),
.Y(n_3861)
);

AOI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3759),
.A2(n_1783),
.B1(n_1784),
.B2(n_1777),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3763),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3751),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_SL g3865 ( 
.A1(n_3771),
.A2(n_3756),
.B1(n_3770),
.B2(n_3776),
.Y(n_3865)
);

INVx3_ASAP7_75t_L g3866 ( 
.A(n_3807),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3767),
.Y(n_3867)
);

INVx2_ASAP7_75t_SL g3868 ( 
.A(n_3780),
.Y(n_3868)
);

INVx3_ASAP7_75t_L g3869 ( 
.A(n_3784),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3814),
.B(n_1788),
.Y(n_3870)
);

INVx3_ASAP7_75t_SL g3871 ( 
.A(n_3753),
.Y(n_3871)
);

BUFx2_ASAP7_75t_SL g3872 ( 
.A(n_3749),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3761),
.Y(n_3873)
);

BUFx2_ASAP7_75t_R g3874 ( 
.A(n_3808),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3789),
.Y(n_3875)
);

AOI22xp5_ASAP7_75t_L g3876 ( 
.A1(n_3815),
.A2(n_1795),
.B1(n_1796),
.B2(n_1792),
.Y(n_3876)
);

INVx3_ASAP7_75t_L g3877 ( 
.A(n_3809),
.Y(n_3877)
);

NAND2x1p5_ASAP7_75t_L g3878 ( 
.A(n_3788),
.B(n_3694),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3766),
.Y(n_3879)
);

OA21x2_ASAP7_75t_L g3880 ( 
.A1(n_3768),
.A2(n_1800),
.B(n_1799),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3795),
.Y(n_3881)
);

INVx2_ASAP7_75t_SL g3882 ( 
.A(n_3744),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3793),
.Y(n_3883)
);

INVx2_ASAP7_75t_SL g3884 ( 
.A(n_3752),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3742),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3765),
.Y(n_3886)
);

OAI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3779),
.A2(n_3694),
.B(n_1804),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3773),
.B(n_16),
.Y(n_3888)
);

INVx1_ASAP7_75t_SL g3889 ( 
.A(n_3811),
.Y(n_3889)
);

BUFx2_ASAP7_75t_L g3890 ( 
.A(n_3773),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3757),
.Y(n_3891)
);

BUFx3_ASAP7_75t_L g3892 ( 
.A(n_3796),
.Y(n_3892)
);

BUFx2_ASAP7_75t_L g3893 ( 
.A(n_3890),
.Y(n_3893)
);

CKINVDCx20_ASAP7_75t_R g3894 ( 
.A(n_3819),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3855),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3828),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3825),
.Y(n_3897)
);

AOI22xp33_ASAP7_75t_SL g3898 ( 
.A1(n_3872),
.A2(n_1805),
.B1(n_1809),
.B2(n_1801),
.Y(n_3898)
);

OAI22xp5_ASAP7_75t_L g3899 ( 
.A1(n_3878),
.A2(n_1815),
.B1(n_1822),
.B2(n_1814),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3891),
.Y(n_3900)
);

OAI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_3843),
.A2(n_1826),
.B1(n_1827),
.B2(n_1824),
.Y(n_3901)
);

AOI22xp33_ASAP7_75t_L g3902 ( 
.A1(n_3823),
.A2(n_2032),
.B1(n_2035),
.B2(n_2031),
.Y(n_3902)
);

OAI21xp33_ASAP7_75t_L g3903 ( 
.A1(n_3850),
.A2(n_1830),
.B(n_1829),
.Y(n_3903)
);

INVx2_ASAP7_75t_SL g3904 ( 
.A(n_3827),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_SL g3905 ( 
.A1(n_3881),
.A2(n_1835),
.B1(n_1840),
.B2(n_1834),
.Y(n_3905)
);

OAI21xp5_ASAP7_75t_SL g3906 ( 
.A1(n_3876),
.A2(n_16),
.B(n_17),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3884),
.A2(n_2074),
.B1(n_2077),
.B2(n_2066),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3817),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3883),
.A2(n_2080),
.B1(n_2078),
.B2(n_1845),
.Y(n_3909)
);

AOI222xp33_ASAP7_75t_L g3910 ( 
.A1(n_3886),
.A2(n_1853),
.B1(n_1846),
.B2(n_1855),
.C1(n_1852),
.C2(n_1842),
.Y(n_3910)
);

HB1xp67_ASAP7_75t_L g3911 ( 
.A(n_3821),
.Y(n_3911)
);

AND2x4_ASAP7_75t_SL g3912 ( 
.A(n_3824),
.B(n_963),
.Y(n_3912)
);

BUFx6f_ASAP7_75t_L g3913 ( 
.A(n_3836),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3843),
.A2(n_1861),
.B1(n_1864),
.B2(n_1858),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3829),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3844),
.Y(n_3916)
);

INVx4_ASAP7_75t_R g3917 ( 
.A(n_3889),
.Y(n_3917)
);

CKINVDCx11_ASAP7_75t_R g3918 ( 
.A(n_3835),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3885),
.A2(n_3830),
.B1(n_3882),
.B2(n_3880),
.Y(n_3919)
);

AOI22xp33_ASAP7_75t_SL g3920 ( 
.A1(n_3875),
.A2(n_1871),
.B1(n_1882),
.B2(n_1868),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3832),
.B(n_17),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3857),
.B(n_18),
.Y(n_3922)
);

INVx4_ASAP7_75t_L g3923 ( 
.A(n_3820),
.Y(n_3923)
);

AOI22xp33_ASAP7_75t_SL g3924 ( 
.A1(n_3851),
.A2(n_1888),
.B1(n_1889),
.B2(n_1884),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3877),
.A2(n_1993),
.B1(n_2000),
.B2(n_1987),
.Y(n_3925)
);

OAI21xp5_ASAP7_75t_SL g3926 ( 
.A1(n_3826),
.A2(n_18),
.B(n_20),
.Y(n_3926)
);

INVx1_ASAP7_75t_SL g3927 ( 
.A(n_3818),
.Y(n_3927)
);

NOR2x1_ASAP7_75t_L g3928 ( 
.A(n_3838),
.B(n_20),
.Y(n_3928)
);

AOI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3868),
.A2(n_2018),
.B1(n_2019),
.B2(n_2013),
.Y(n_3929)
);

BUFx2_ASAP7_75t_L g3930 ( 
.A(n_3841),
.Y(n_3930)
);

INVx4_ASAP7_75t_L g3931 ( 
.A(n_3839),
.Y(n_3931)
);

OAI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3879),
.A2(n_1893),
.B1(n_1898),
.B2(n_1891),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3842),
.Y(n_3933)
);

AOI22xp33_ASAP7_75t_L g3934 ( 
.A1(n_3887),
.A2(n_2052),
.B1(n_2057),
.B2(n_2044),
.Y(n_3934)
);

INVxp67_ASAP7_75t_L g3935 ( 
.A(n_3846),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3888),
.B(n_1899),
.Y(n_3936)
);

AOI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3865),
.A2(n_1910),
.B1(n_1918),
.B2(n_1906),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3892),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3854),
.A2(n_3862),
.B1(n_3847),
.B2(n_3833),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3840),
.Y(n_3940)
);

OAI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3834),
.A2(n_1924),
.B1(n_1931),
.B2(n_1923),
.Y(n_3941)
);

BUFx4f_ASAP7_75t_SL g3942 ( 
.A(n_3871),
.Y(n_3942)
);

BUFx6f_ASAP7_75t_L g3943 ( 
.A(n_3816),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3845),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3853),
.A2(n_1982),
.B1(n_1983),
.B2(n_1979),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3858),
.B(n_1935),
.Y(n_3946)
);

INVx2_ASAP7_75t_SL g3947 ( 
.A(n_3837),
.Y(n_3947)
);

NOR2x1_ASAP7_75t_R g3948 ( 
.A(n_3874),
.B(n_1937),
.Y(n_3948)
);

OAI22xp5_ASAP7_75t_L g3949 ( 
.A1(n_3849),
.A2(n_1942),
.B1(n_1943),
.B2(n_1939),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3867),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3861),
.Y(n_3951)
);

OAI22xp5_ASAP7_75t_L g3952 ( 
.A1(n_3853),
.A2(n_1947),
.B1(n_1952),
.B2(n_1944),
.Y(n_3952)
);

AOI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3852),
.A2(n_1967),
.B1(n_1970),
.B2(n_1964),
.Y(n_3953)
);

BUFx2_ASAP7_75t_L g3954 ( 
.A(n_3866),
.Y(n_3954)
);

OAI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3831),
.A2(n_1959),
.B1(n_1962),
.B2(n_1953),
.Y(n_3955)
);

AOI22xp33_ASAP7_75t_L g3956 ( 
.A1(n_3863),
.A2(n_1978),
.B1(n_1984),
.B2(n_1977),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3856),
.A2(n_1973),
.B1(n_1975),
.B2(n_1972),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3859),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3848),
.A2(n_2043),
.B1(n_2065),
.B2(n_2039),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_R g3960 ( 
.A(n_3918),
.B(n_3942),
.Y(n_3960)
);

INVxp67_ASAP7_75t_L g3961 ( 
.A(n_3893),
.Y(n_3961)
);

NAND2xp33_ASAP7_75t_R g3962 ( 
.A(n_3930),
.B(n_3870),
.Y(n_3962)
);

INVxp67_ASAP7_75t_L g3963 ( 
.A(n_3911),
.Y(n_3963)
);

AND2x4_ASAP7_75t_L g3964 ( 
.A(n_3933),
.B(n_3873),
.Y(n_3964)
);

OR2x6_ASAP7_75t_L g3965 ( 
.A(n_3904),
.B(n_3928),
.Y(n_3965)
);

NAND2xp33_ASAP7_75t_R g3966 ( 
.A(n_3938),
.B(n_3869),
.Y(n_3966)
);

AND2x4_ASAP7_75t_L g3967 ( 
.A(n_3897),
.B(n_3860),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3935),
.B(n_3864),
.Y(n_3968)
);

NAND2xp33_ASAP7_75t_R g3969 ( 
.A(n_3948),
.B(n_23),
.Y(n_3969)
);

INVxp67_ASAP7_75t_L g3970 ( 
.A(n_3936),
.Y(n_3970)
);

AND2x4_ASAP7_75t_L g3971 ( 
.A(n_3947),
.B(n_3822),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3895),
.B(n_2001),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3896),
.B(n_2006),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3900),
.B(n_2027),
.Y(n_3974)
);

OR2x2_ASAP7_75t_L g3975 ( 
.A(n_3951),
.B(n_25),
.Y(n_3975)
);

NOR2xp33_ASAP7_75t_R g3976 ( 
.A(n_3894),
.B(n_26),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3916),
.Y(n_3977)
);

NAND2xp33_ASAP7_75t_R g3978 ( 
.A(n_3921),
.B(n_26),
.Y(n_3978)
);

AND2x2_ASAP7_75t_SL g3979 ( 
.A(n_3919),
.B(n_27),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_R g3980 ( 
.A(n_3927),
.B(n_27),
.Y(n_3980)
);

CKINVDCx5p33_ASAP7_75t_R g3981 ( 
.A(n_3923),
.Y(n_3981)
);

OR2x6_ASAP7_75t_L g3982 ( 
.A(n_3943),
.B(n_3931),
.Y(n_3982)
);

NAND2xp33_ASAP7_75t_R g3983 ( 
.A(n_3922),
.B(n_28),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_R g3984 ( 
.A(n_3943),
.B(n_29),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3908),
.B(n_29),
.Y(n_3985)
);

INVx2_ASAP7_75t_L g3986 ( 
.A(n_3940),
.Y(n_3986)
);

OR2x6_ASAP7_75t_L g3987 ( 
.A(n_3913),
.B(n_30),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3958),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_3915),
.B(n_30),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3944),
.Y(n_3990)
);

OR2x6_ASAP7_75t_L g3991 ( 
.A(n_3913),
.B(n_31),
.Y(n_3991)
);

INVxp67_ASAP7_75t_L g3992 ( 
.A(n_3946),
.Y(n_3992)
);

INVxp67_ASAP7_75t_L g3993 ( 
.A(n_3949),
.Y(n_3993)
);

NOR2xp33_ASAP7_75t_R g3994 ( 
.A(n_3945),
.B(n_3939),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_SL g3995 ( 
.A(n_3899),
.B(n_3898),
.Y(n_3995)
);

BUFx3_ASAP7_75t_L g3996 ( 
.A(n_3912),
.Y(n_3996)
);

NOR2xp33_ASAP7_75t_R g3997 ( 
.A(n_3917),
.B(n_32),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3950),
.B(n_3954),
.Y(n_3998)
);

BUFx3_ASAP7_75t_L g3999 ( 
.A(n_3952),
.Y(n_3999)
);

OR2x4_ASAP7_75t_L g4000 ( 
.A(n_3926),
.B(n_32),
.Y(n_4000)
);

NOR2xp33_ASAP7_75t_R g4001 ( 
.A(n_3907),
.B(n_34),
.Y(n_4001)
);

CKINVDCx16_ASAP7_75t_R g4002 ( 
.A(n_3901),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_L g4003 ( 
.A(n_3914),
.B(n_35),
.Y(n_4003)
);

OR2x6_ASAP7_75t_L g4004 ( 
.A(n_3906),
.B(n_36),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3902),
.B(n_36),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3937),
.B(n_3905),
.Y(n_4006)
);

BUFx10_ASAP7_75t_L g4007 ( 
.A(n_3941),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3903),
.Y(n_4008)
);

BUFx3_ASAP7_75t_L g4009 ( 
.A(n_3932),
.Y(n_4009)
);

INVxp67_ASAP7_75t_L g4010 ( 
.A(n_3910),
.Y(n_4010)
);

NOR2xp33_ASAP7_75t_R g4011 ( 
.A(n_3959),
.B(n_37),
.Y(n_4011)
);

NAND2xp33_ASAP7_75t_R g4012 ( 
.A(n_3920),
.B(n_37),
.Y(n_4012)
);

NOR2xp33_ASAP7_75t_R g4013 ( 
.A(n_3929),
.B(n_39),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3924),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_L g4015 ( 
.A(n_3957),
.B(n_41),
.Y(n_4015)
);

NAND2xp33_ASAP7_75t_R g4016 ( 
.A(n_3909),
.B(n_41),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3956),
.B(n_42),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3934),
.B(n_43),
.Y(n_4018)
);

NOR2xp33_ASAP7_75t_R g4019 ( 
.A(n_3953),
.B(n_43),
.Y(n_4019)
);

XNOR2xp5_ASAP7_75t_L g4020 ( 
.A(n_3955),
.B(n_45),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3925),
.B(n_45),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3916),
.Y(n_4022)
);

INVxp67_ASAP7_75t_L g4023 ( 
.A(n_3893),
.Y(n_4023)
);

NOR2xp33_ASAP7_75t_L g4024 ( 
.A(n_3923),
.B(n_46),
.Y(n_4024)
);

AND2x4_ASAP7_75t_L g4025 ( 
.A(n_3933),
.B(n_47),
.Y(n_4025)
);

AND2x4_ASAP7_75t_L g4026 ( 
.A(n_3933),
.B(n_48),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3893),
.B(n_49),
.Y(n_4027)
);

INVxp67_ASAP7_75t_L g4028 ( 
.A(n_3893),
.Y(n_4028)
);

INVxp67_ASAP7_75t_L g4029 ( 
.A(n_3893),
.Y(n_4029)
);

NAND2xp33_ASAP7_75t_R g4030 ( 
.A(n_3893),
.B(n_49),
.Y(n_4030)
);

NAND2xp33_ASAP7_75t_R g4031 ( 
.A(n_3893),
.B(n_50),
.Y(n_4031)
);

BUFx3_ASAP7_75t_L g4032 ( 
.A(n_3918),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_R g4033 ( 
.A(n_3918),
.B(n_50),
.Y(n_4033)
);

INVx2_ASAP7_75t_SL g4034 ( 
.A(n_3917),
.Y(n_4034)
);

INVxp67_ASAP7_75t_L g4035 ( 
.A(n_3893),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3916),
.Y(n_4036)
);

BUFx3_ASAP7_75t_L g4037 ( 
.A(n_3918),
.Y(n_4037)
);

NAND2xp33_ASAP7_75t_R g4038 ( 
.A(n_3893),
.B(n_51),
.Y(n_4038)
);

NAND2xp33_ASAP7_75t_R g4039 ( 
.A(n_3893),
.B(n_52),
.Y(n_4039)
);

NAND2xp33_ASAP7_75t_R g4040 ( 
.A(n_3893),
.B(n_53),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3893),
.B(n_54),
.Y(n_4041)
);

NAND2xp33_ASAP7_75t_R g4042 ( 
.A(n_3893),
.B(n_55),
.Y(n_4042)
);

NOR2xp33_ASAP7_75t_R g4043 ( 
.A(n_3918),
.B(n_55),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_R g4044 ( 
.A(n_3918),
.B(n_56),
.Y(n_4044)
);

AND2x4_ASAP7_75t_L g4045 ( 
.A(n_3933),
.B(n_56),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3916),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3911),
.B(n_57),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3916),
.Y(n_4048)
);

XNOR2xp5_ASAP7_75t_L g4049 ( 
.A(n_3894),
.B(n_57),
.Y(n_4049)
);

INVxp67_ASAP7_75t_L g4050 ( 
.A(n_3893),
.Y(n_4050)
);

NAND2xp33_ASAP7_75t_R g4051 ( 
.A(n_3893),
.B(n_58),
.Y(n_4051)
);

AND2x4_ASAP7_75t_L g4052 ( 
.A(n_3933),
.B(n_58),
.Y(n_4052)
);

NAND2xp33_ASAP7_75t_R g4053 ( 
.A(n_3893),
.B(n_59),
.Y(n_4053)
);

INVxp67_ASAP7_75t_L g4054 ( 
.A(n_3893),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3916),
.Y(n_4055)
);

NAND2xp33_ASAP7_75t_R g4056 ( 
.A(n_3893),
.B(n_59),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3911),
.B(n_60),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_R g4058 ( 
.A(n_3918),
.B(n_60),
.Y(n_4058)
);

AND2x4_ASAP7_75t_L g4059 ( 
.A(n_3933),
.B(n_61),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_R g4060 ( 
.A(n_3918),
.B(n_61),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_R g4061 ( 
.A(n_3918),
.B(n_63),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3893),
.B(n_65),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_3893),
.B(n_65),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3893),
.B(n_68),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3916),
.Y(n_4065)
);

AND2x4_ASAP7_75t_L g4066 ( 
.A(n_3933),
.B(n_68),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3911),
.B(n_69),
.Y(n_4067)
);

AND2x4_ASAP7_75t_L g4068 ( 
.A(n_3933),
.B(n_70),
.Y(n_4068)
);

NAND2xp33_ASAP7_75t_R g4069 ( 
.A(n_3893),
.B(n_70),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_R g4070 ( 
.A(n_3918),
.B(n_71),
.Y(n_4070)
);

AND2x4_ASAP7_75t_L g4071 ( 
.A(n_3933),
.B(n_71),
.Y(n_4071)
);

INVxp67_ASAP7_75t_L g4072 ( 
.A(n_3893),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3893),
.B(n_73),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3916),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_3919),
.B(n_75),
.Y(n_4075)
);

XNOR2xp5_ASAP7_75t_L g4076 ( 
.A(n_3894),
.B(n_76),
.Y(n_4076)
);

BUFx3_ASAP7_75t_L g4077 ( 
.A(n_3918),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3964),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3961),
.B(n_4023),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_4028),
.B(n_76),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3992),
.B(n_77),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_4029),
.B(n_77),
.Y(n_4082)
);

OR2x2_ASAP7_75t_L g4083 ( 
.A(n_3963),
.B(n_78),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3977),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3967),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4035),
.B(n_80),
.Y(n_4086)
);

INVx3_ASAP7_75t_L g4087 ( 
.A(n_3982),
.Y(n_4087)
);

BUFx2_ASAP7_75t_SL g4088 ( 
.A(n_4034),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3986),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_4022),
.Y(n_4090)
);

BUFx2_ASAP7_75t_L g4091 ( 
.A(n_3965),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_4050),
.B(n_80),
.Y(n_4092)
);

INVxp67_ASAP7_75t_SL g4093 ( 
.A(n_4030),
.Y(n_4093)
);

INVxp67_ASAP7_75t_SL g4094 ( 
.A(n_4031),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_4054),
.B(n_82),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_4036),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_4072),
.B(n_82),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4046),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_4010),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_3965),
.B(n_85),
.Y(n_4100)
);

HB1xp67_ASAP7_75t_L g4101 ( 
.A(n_3990),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3968),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3971),
.B(n_86),
.Y(n_4103)
);

BUFx6f_ASAP7_75t_L g4104 ( 
.A(n_4032),
.Y(n_4104)
);

INVxp67_ASAP7_75t_L g4105 ( 
.A(n_4038),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_4048),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4055),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_4065),
.Y(n_4108)
);

OR2x2_ASAP7_75t_L g4109 ( 
.A(n_4074),
.B(n_86),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_3982),
.B(n_87),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3988),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3985),
.Y(n_4112)
);

BUFx2_ASAP7_75t_L g4113 ( 
.A(n_3997),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3975),
.Y(n_4114)
);

HB1xp67_ASAP7_75t_L g4115 ( 
.A(n_4027),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3998),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_3989),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3973),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3974),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_4041),
.B(n_87),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3972),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_4004),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_4047),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4062),
.B(n_88),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_4025),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4057),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4026),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4063),
.B(n_90),
.Y(n_4128)
);

BUFx2_ASAP7_75t_L g4129 ( 
.A(n_3960),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_4067),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_4064),
.B(n_91),
.Y(n_4131)
);

BUFx2_ASAP7_75t_L g4132 ( 
.A(n_4037),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4073),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_4045),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_4052),
.Y(n_4135)
);

OR2x2_ASAP7_75t_L g4136 ( 
.A(n_3970),
.B(n_92),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4075),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4059),
.Y(n_4138)
);

BUFx2_ASAP7_75t_L g4139 ( 
.A(n_4077),
.Y(n_4139)
);

AND2x2_ASAP7_75t_L g4140 ( 
.A(n_3996),
.B(n_93),
.Y(n_4140)
);

INVx4_ASAP7_75t_R g4141 ( 
.A(n_4039),
.Y(n_4141)
);

AND2x2_ASAP7_75t_L g4142 ( 
.A(n_4066),
.B(n_93),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4068),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4071),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4008),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_3981),
.B(n_94),
.Y(n_4146)
);

OR2x2_ASAP7_75t_L g4147 ( 
.A(n_3993),
.B(n_95),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_4002),
.B(n_95),
.Y(n_4148)
);

BUFx3_ASAP7_75t_L g4149 ( 
.A(n_3987),
.Y(n_4149)
);

BUFx2_ASAP7_75t_L g4150 ( 
.A(n_4033),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_4014),
.B(n_96),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4009),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3979),
.Y(n_4153)
);

NAND2x1p5_ASAP7_75t_L g4154 ( 
.A(n_4040),
.B(n_97),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3987),
.Y(n_4155)
);

INVx3_ASAP7_75t_L g4156 ( 
.A(n_3991),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3991),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3999),
.B(n_97),
.Y(n_4158)
);

AO31x2_ASAP7_75t_L g4159 ( 
.A1(n_4024),
.A2(n_101),
.A3(n_98),
.B(n_100),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4007),
.B(n_98),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4000),
.Y(n_4161)
);

AO31x2_ASAP7_75t_L g4162 ( 
.A1(n_4042),
.A2(n_103),
.A3(n_101),
.B(n_102),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3994),
.B(n_102),
.Y(n_4163)
);

BUFx3_ASAP7_75t_L g4164 ( 
.A(n_4049),
.Y(n_4164)
);

AND2x2_ASAP7_75t_L g4165 ( 
.A(n_4043),
.B(n_103),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4004),
.Y(n_4166)
);

BUFx6f_ASAP7_75t_L g4167 ( 
.A(n_4006),
.Y(n_4167)
);

BUFx2_ASAP7_75t_L g4168 ( 
.A(n_4044),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4021),
.Y(n_4169)
);

OR2x2_ASAP7_75t_L g4170 ( 
.A(n_4005),
.B(n_104),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4018),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_4058),
.B(n_4060),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_4061),
.B(n_104),
.Y(n_4173)
);

CKINVDCx16_ASAP7_75t_R g4174 ( 
.A(n_4070),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4017),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4003),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_3984),
.B(n_105),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3995),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_3980),
.B(n_106),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3976),
.B(n_107),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4076),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_3966),
.B(n_107),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_4020),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4015),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_4051),
.Y(n_4185)
);

AOI22xp33_ASAP7_75t_SL g4186 ( 
.A1(n_4001),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4013),
.Y(n_4187)
);

INVx3_ASAP7_75t_L g4188 ( 
.A(n_4053),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4011),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_4056),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_4069),
.Y(n_4191)
);

OR2x2_ASAP7_75t_L g4192 ( 
.A(n_3962),
.B(n_108),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4019),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3983),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_3978),
.B(n_109),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4016),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_4012),
.B(n_110),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_3969),
.B(n_111),
.Y(n_4198)
);

HB1xp67_ASAP7_75t_L g4199 ( 
.A(n_3965),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3977),
.Y(n_4200)
);

AOI22xp33_ASAP7_75t_L g4201 ( 
.A1(n_4010),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_4201)
);

AND2x2_ASAP7_75t_L g4202 ( 
.A(n_3961),
.B(n_112),
.Y(n_4202)
);

AND2x4_ASAP7_75t_L g4203 ( 
.A(n_4034),
.B(n_114),
.Y(n_4203)
);

INVx3_ASAP7_75t_L g4204 ( 
.A(n_3982),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3977),
.Y(n_4205)
);

AND2x4_ASAP7_75t_L g4206 ( 
.A(n_4034),
.B(n_114),
.Y(n_4206)
);

OR2x2_ASAP7_75t_L g4207 ( 
.A(n_3963),
.B(n_115),
.Y(n_4207)
);

INVx2_ASAP7_75t_SL g4208 ( 
.A(n_3982),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3977),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3977),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3977),
.Y(n_4211)
);

BUFx3_ASAP7_75t_L g4212 ( 
.A(n_4032),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3977),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_3964),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3992),
.B(n_116),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_3964),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3964),
.Y(n_4217)
);

BUFx2_ASAP7_75t_L g4218 ( 
.A(n_3965),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_3961),
.B(n_116),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_3961),
.B(n_117),
.Y(n_4220)
);

OAI21x1_ASAP7_75t_L g4221 ( 
.A1(n_3998),
.A2(n_118),
.B(n_119),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_3961),
.B(n_118),
.Y(n_4222)
);

OR2x2_ASAP7_75t_L g4223 ( 
.A(n_3963),
.B(n_119),
.Y(n_4223)
);

AND2x4_ASAP7_75t_SL g4224 ( 
.A(n_3982),
.B(n_120),
.Y(n_4224)
);

BUFx3_ASAP7_75t_L g4225 ( 
.A(n_4032),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_3961),
.B(n_121),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3977),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3977),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_3961),
.B(n_122),
.Y(n_4229)
);

INVx2_ASAP7_75t_SL g4230 ( 
.A(n_3982),
.Y(n_4230)
);

INVx1_ASAP7_75t_SL g4231 ( 
.A(n_3997),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_3964),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3977),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3977),
.Y(n_4234)
);

OR2x2_ASAP7_75t_L g4235 ( 
.A(n_3963),
.B(n_122),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_3964),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3977),
.Y(n_4237)
);

OR2x2_ASAP7_75t_L g4238 ( 
.A(n_3963),
.B(n_123),
.Y(n_4238)
);

OR2x2_ASAP7_75t_L g4239 ( 
.A(n_4116),
.B(n_123),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4132),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4088),
.B(n_124),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_4087),
.B(n_4204),
.Y(n_4242)
);

NOR2xp33_ASAP7_75t_SL g4243 ( 
.A(n_4174),
.B(n_124),
.Y(n_4243)
);

INVx4_ASAP7_75t_L g4244 ( 
.A(n_4104),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4208),
.B(n_125),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4101),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_4230),
.B(n_126),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4091),
.B(n_126),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_4218),
.B(n_127),
.Y(n_4249)
);

AND2x2_ASAP7_75t_L g4250 ( 
.A(n_4199),
.B(n_127),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4114),
.B(n_4145),
.Y(n_4251)
);

AND2x4_ASAP7_75t_SL g4252 ( 
.A(n_4104),
.B(n_128),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4084),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4090),
.Y(n_4254)
);

BUFx2_ASAP7_75t_SL g4255 ( 
.A(n_4172),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4079),
.B(n_128),
.Y(n_4256)
);

INVx2_ASAP7_75t_SL g4257 ( 
.A(n_4212),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4096),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_4152),
.B(n_129),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4178),
.B(n_129),
.Y(n_4260)
);

INVx8_ASAP7_75t_L g4261 ( 
.A(n_4165),
.Y(n_4261)
);

OR2x2_ASAP7_75t_L g4262 ( 
.A(n_4115),
.B(n_130),
.Y(n_4262)
);

HB1xp67_ASAP7_75t_L g4263 ( 
.A(n_4194),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4078),
.B(n_131),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4214),
.B(n_131),
.Y(n_4265)
);

BUFx2_ASAP7_75t_L g4266 ( 
.A(n_4093),
.Y(n_4266)
);

INVx3_ASAP7_75t_L g4267 ( 
.A(n_4225),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4137),
.B(n_132),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4098),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4139),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4094),
.B(n_132),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4216),
.B(n_133),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4106),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4107),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_4156),
.Y(n_4275)
);

BUFx2_ASAP7_75t_L g4276 ( 
.A(n_4188),
.Y(n_4276)
);

HB1xp67_ASAP7_75t_L g4277 ( 
.A(n_4185),
.Y(n_4277)
);

OR2x2_ASAP7_75t_L g4278 ( 
.A(n_4112),
.B(n_4123),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4217),
.B(n_133),
.Y(n_4279)
);

OR2x2_ASAP7_75t_L g4280 ( 
.A(n_4126),
.B(n_4130),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4108),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4200),
.Y(n_4282)
);

BUFx3_ASAP7_75t_L g4283 ( 
.A(n_4129),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4232),
.B(n_134),
.Y(n_4284)
);

OR2x2_ASAP7_75t_L g4285 ( 
.A(n_4171),
.B(n_135),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4149),
.Y(n_4286)
);

INVxp67_ASAP7_75t_SL g4287 ( 
.A(n_4105),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4205),
.Y(n_4288)
);

AND2x4_ASAP7_75t_L g4289 ( 
.A(n_4155),
.B(n_135),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4209),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4236),
.B(n_136),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4167),
.B(n_137),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4085),
.B(n_138),
.Y(n_4293)
);

AOI22xp33_ASAP7_75t_SL g4294 ( 
.A1(n_4190),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4210),
.Y(n_4295)
);

INVx3_ASAP7_75t_L g4296 ( 
.A(n_4154),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4167),
.B(n_139),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_4191),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4157),
.Y(n_4299)
);

BUFx2_ASAP7_75t_L g4300 ( 
.A(n_4113),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4211),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4213),
.Y(n_4302)
);

NAND2x1_ASAP7_75t_L g4303 ( 
.A(n_4141),
.B(n_140),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4166),
.B(n_141),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4102),
.B(n_142),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4118),
.B(n_143),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4089),
.Y(n_4307)
);

AND2x4_ASAP7_75t_L g4308 ( 
.A(n_4125),
.B(n_143),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4119),
.B(n_144),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4150),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4121),
.B(n_144),
.Y(n_4311)
);

OR2x2_ASAP7_75t_L g4312 ( 
.A(n_4169),
.B(n_145),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4227),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4168),
.Y(n_4314)
);

INVxp67_ASAP7_75t_L g4315 ( 
.A(n_4192),
.Y(n_4315)
);

BUFx2_ASAP7_75t_L g4316 ( 
.A(n_4162),
.Y(n_4316)
);

NOR2xp33_ASAP7_75t_L g4317 ( 
.A(n_4231),
.B(n_145),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4228),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4111),
.Y(n_4319)
);

HB1xp67_ASAP7_75t_L g4320 ( 
.A(n_4233),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4117),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4175),
.B(n_146),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4133),
.B(n_146),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4176),
.B(n_147),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4184),
.B(n_148),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4234),
.Y(n_4326)
);

OR2x2_ASAP7_75t_L g4327 ( 
.A(n_4237),
.B(n_150),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4153),
.B(n_150),
.Y(n_4328)
);

OR2x2_ASAP7_75t_L g4329 ( 
.A(n_4109),
.B(n_151),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4083),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4207),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4182),
.B(n_151),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4223),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4235),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4238),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4127),
.B(n_153),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4100),
.B(n_154),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4136),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4097),
.B(n_154),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4134),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4080),
.Y(n_4341)
);

AND2x4_ASAP7_75t_L g4342 ( 
.A(n_4135),
.B(n_4138),
.Y(n_4342)
);

AND2x2_ASAP7_75t_SL g4343 ( 
.A(n_4197),
.B(n_155),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4143),
.B(n_4144),
.Y(n_4344)
);

INVxp67_ASAP7_75t_SL g4345 ( 
.A(n_4196),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_4221),
.B(n_155),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4082),
.Y(n_4347)
);

HB1xp67_ASAP7_75t_L g4348 ( 
.A(n_4162),
.Y(n_4348)
);

INVxp67_ASAP7_75t_SL g4349 ( 
.A(n_4160),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4086),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4103),
.B(n_158),
.Y(n_4351)
);

BUFx6f_ASAP7_75t_L g4352 ( 
.A(n_4203),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4092),
.Y(n_4353)
);

BUFx2_ASAP7_75t_L g4354 ( 
.A(n_4161),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4095),
.B(n_158),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_4202),
.B(n_159),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4206),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_4110),
.Y(n_4358)
);

AND2x4_ASAP7_75t_L g4359 ( 
.A(n_4219),
.B(n_160),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4220),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4222),
.B(n_160),
.Y(n_4361)
);

AND2x4_ASAP7_75t_L g4362 ( 
.A(n_4226),
.B(n_161),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4229),
.B(n_161),
.Y(n_4363)
);

INVxp67_ASAP7_75t_L g4364 ( 
.A(n_4148),
.Y(n_4364)
);

AND2x4_ASAP7_75t_L g4365 ( 
.A(n_4140),
.B(n_162),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4147),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4120),
.B(n_4124),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4081),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_L g4369 ( 
.A(n_4163),
.B(n_162),
.Y(n_4369)
);

OR2x2_ASAP7_75t_L g4370 ( 
.A(n_4170),
.B(n_163),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4215),
.Y(n_4371)
);

HB1xp67_ASAP7_75t_L g4372 ( 
.A(n_4159),
.Y(n_4372)
);

BUFx2_ASAP7_75t_L g4373 ( 
.A(n_4189),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_4128),
.B(n_164),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4159),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4224),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4131),
.B(n_165),
.Y(n_4377)
);

INVxp67_ASAP7_75t_L g4378 ( 
.A(n_4195),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_4193),
.B(n_165),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4187),
.B(n_167),
.Y(n_4380)
);

BUFx2_ASAP7_75t_L g4381 ( 
.A(n_4146),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4142),
.B(n_4158),
.Y(n_4382)
);

INVx2_ASAP7_75t_L g4383 ( 
.A(n_4198),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4164),
.Y(n_4384)
);

OAI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_4122),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4151),
.Y(n_4386)
);

OR2x2_ASAP7_75t_L g4387 ( 
.A(n_4181),
.B(n_169),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4173),
.Y(n_4388)
);

INVx3_ASAP7_75t_L g4389 ( 
.A(n_4177),
.Y(n_4389)
);

INVx3_ASAP7_75t_L g4390 ( 
.A(n_4179),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4183),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4180),
.B(n_170),
.Y(n_4392)
);

INVxp67_ASAP7_75t_SL g4393 ( 
.A(n_4186),
.Y(n_4393)
);

INVx2_ASAP7_75t_L g4394 ( 
.A(n_4099),
.Y(n_4394)
);

INVx3_ASAP7_75t_L g4395 ( 
.A(n_4201),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4088),
.B(n_171),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4088),
.B(n_172),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4132),
.Y(n_4398)
);

INVxp67_ASAP7_75t_L g4399 ( 
.A(n_4093),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4101),
.Y(n_4400)
);

AND2x4_ASAP7_75t_L g4401 ( 
.A(n_4208),
.B(n_173),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4178),
.B(n_173),
.Y(n_4402)
);

OAI221xp5_ASAP7_75t_L g4403 ( 
.A1(n_4093),
.A2(n_177),
.B1(n_174),
.B2(n_176),
.C(n_178),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4132),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4088),
.B(n_178),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4101),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4088),
.B(n_179),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4101),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4088),
.B(n_179),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4101),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_4178),
.B(n_180),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4101),
.Y(n_4412)
);

AND2x4_ASAP7_75t_L g4413 ( 
.A(n_4208),
.B(n_181),
.Y(n_4413)
);

AND2x4_ASAP7_75t_L g4414 ( 
.A(n_4208),
.B(n_181),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4101),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4132),
.Y(n_4416)
);

INVx1_ASAP7_75t_SL g4417 ( 
.A(n_4113),
.Y(n_4417)
);

AND2x4_ASAP7_75t_L g4418 ( 
.A(n_4208),
.B(n_182),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4208),
.B(n_182),
.Y(n_4419)
);

OR2x2_ASAP7_75t_L g4420 ( 
.A(n_4116),
.B(n_183),
.Y(n_4420)
);

OR2x2_ASAP7_75t_L g4421 ( 
.A(n_4116),
.B(n_183),
.Y(n_4421)
);

NAND2xp33_ASAP7_75t_L g4422 ( 
.A(n_4192),
.B(n_185),
.Y(n_4422)
);

AND2x4_ASAP7_75t_L g4423 ( 
.A(n_4208),
.B(n_186),
.Y(n_4423)
);

HB1xp67_ASAP7_75t_L g4424 ( 
.A(n_4115),
.Y(n_4424)
);

INVx3_ASAP7_75t_L g4425 ( 
.A(n_4212),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4088),
.B(n_186),
.Y(n_4426)
);

INVx4_ASAP7_75t_L g4427 ( 
.A(n_4104),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4088),
.B(n_187),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_4132),
.Y(n_4429)
);

AND2x4_ASAP7_75t_L g4430 ( 
.A(n_4208),
.B(n_187),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4101),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4088),
.B(n_188),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4101),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_4283),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_4266),
.B(n_188),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4424),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4244),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4300),
.B(n_189),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4417),
.B(n_190),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_SL g4440 ( 
.A(n_4267),
.B(n_190),
.Y(n_4440)
);

HB1xp67_ASAP7_75t_L g4441 ( 
.A(n_4277),
.Y(n_4441)
);

INVx2_ASAP7_75t_SL g4442 ( 
.A(n_4352),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4276),
.B(n_192),
.Y(n_4443)
);

NAND4xp25_ASAP7_75t_L g4444 ( 
.A(n_4399),
.B(n_195),
.C(n_193),
.D(n_194),
.Y(n_4444)
);

AND2x4_ASAP7_75t_L g4445 ( 
.A(n_4257),
.B(n_193),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4427),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4263),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4425),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4287),
.B(n_4378),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4310),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4320),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4242),
.B(n_196),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4251),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4314),
.B(n_196),
.Y(n_4454)
);

OR2x2_ASAP7_75t_L g4455 ( 
.A(n_4345),
.B(n_197),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4296),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4383),
.B(n_198),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4381),
.B(n_199),
.Y(n_4458)
);

OR2x2_ASAP7_75t_L g4459 ( 
.A(n_4298),
.B(n_199),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4389),
.B(n_200),
.Y(n_4460)
);

INVx3_ASAP7_75t_L g4461 ( 
.A(n_4352),
.Y(n_4461)
);

AND2x2_ASAP7_75t_L g4462 ( 
.A(n_4240),
.B(n_200),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4388),
.Y(n_4463)
);

AND2x4_ASAP7_75t_SL g4464 ( 
.A(n_4270),
.B(n_201),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_4390),
.B(n_201),
.Y(n_4465)
);

OR2x2_ASAP7_75t_L g4466 ( 
.A(n_4315),
.B(n_202),
.Y(n_4466)
);

OR2x2_ASAP7_75t_L g4467 ( 
.A(n_4349),
.B(n_202),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4398),
.B(n_203),
.Y(n_4468)
);

NAND3xp33_ASAP7_75t_L g4469 ( 
.A(n_4348),
.B(n_4316),
.C(n_4372),
.Y(n_4469)
);

INVx2_ASAP7_75t_L g4470 ( 
.A(n_4404),
.Y(n_4470)
);

OR2x2_ASAP7_75t_L g4471 ( 
.A(n_4354),
.B(n_203),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4416),
.B(n_204),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4429),
.Y(n_4473)
);

BUFx2_ASAP7_75t_L g4474 ( 
.A(n_4261),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4253),
.Y(n_4475)
);

INVxp67_ASAP7_75t_SL g4476 ( 
.A(n_4303),
.Y(n_4476)
);

AND2x4_ASAP7_75t_L g4477 ( 
.A(n_4286),
.B(n_204),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4364),
.B(n_205),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4261),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4393),
.B(n_205),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4254),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4258),
.Y(n_4482)
);

OR2x2_ASAP7_75t_L g4483 ( 
.A(n_4299),
.B(n_207),
.Y(n_4483)
);

OR2x2_ASAP7_75t_L g4484 ( 
.A(n_4321),
.B(n_207),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4384),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4275),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4269),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4373),
.B(n_208),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4273),
.Y(n_4489)
);

OR2x2_ASAP7_75t_L g4490 ( 
.A(n_4340),
.B(n_208),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4382),
.B(n_209),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4255),
.B(n_209),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4395),
.B(n_210),
.Y(n_4493)
);

AND2x4_ASAP7_75t_L g4494 ( 
.A(n_4357),
.B(n_211),
.Y(n_4494)
);

NOR2x1_ASAP7_75t_SL g4495 ( 
.A(n_4375),
.B(n_4246),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4274),
.Y(n_4496)
);

NOR2x1_ASAP7_75t_L g4497 ( 
.A(n_4422),
.B(n_211),
.Y(n_4497)
);

OR2x2_ASAP7_75t_L g4498 ( 
.A(n_4366),
.B(n_212),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4358),
.B(n_213),
.Y(n_4499)
);

INVxp67_ASAP7_75t_L g4500 ( 
.A(n_4243),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4344),
.B(n_213),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4281),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4367),
.B(n_214),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4341),
.B(n_214),
.Y(n_4504)
);

OR2x2_ASAP7_75t_L g4505 ( 
.A(n_4330),
.B(n_215),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_4347),
.B(n_215),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4350),
.B(n_216),
.Y(n_4507)
);

AND2x4_ASAP7_75t_L g4508 ( 
.A(n_4376),
.B(n_217),
.Y(n_4508)
);

INVx2_ASAP7_75t_L g4509 ( 
.A(n_4342),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_L g4510 ( 
.A(n_4353),
.B(n_217),
.Y(n_4510)
);

INVx3_ASAP7_75t_L g4511 ( 
.A(n_4401),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4360),
.B(n_218),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4386),
.B(n_218),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4331),
.B(n_219),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4333),
.B(n_219),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4282),
.Y(n_4516)
);

OR2x2_ASAP7_75t_L g4517 ( 
.A(n_4334),
.B(n_220),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_4335),
.B(n_221),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4288),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4338),
.B(n_222),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4248),
.B(n_4249),
.Y(n_4521)
);

INVx1_ASAP7_75t_L g4522 ( 
.A(n_4290),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4295),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4301),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_4241),
.Y(n_4525)
);

INVx3_ASAP7_75t_L g4526 ( 
.A(n_4413),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4391),
.B(n_222),
.Y(n_4527)
);

OR2x2_ASAP7_75t_L g4528 ( 
.A(n_4368),
.B(n_223),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4250),
.B(n_223),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4371),
.B(n_224),
.Y(n_4530)
);

BUFx2_ASAP7_75t_L g4531 ( 
.A(n_4396),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4256),
.B(n_224),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4397),
.B(n_225),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4302),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4405),
.B(n_225),
.Y(n_4535)
);

OAI22xp5_ASAP7_75t_L g4536 ( 
.A1(n_4394),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4407),
.B(n_226),
.Y(n_4537)
);

NAND2x1p5_ASAP7_75t_L g4538 ( 
.A(n_4409),
.B(n_229),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4343),
.B(n_230),
.Y(n_4539)
);

AND2x4_ASAP7_75t_L g4540 ( 
.A(n_4426),
.B(n_231),
.Y(n_4540)
);

INVx1_ASAP7_75t_SL g4541 ( 
.A(n_4428),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4313),
.Y(n_4542)
);

OR2x2_ASAP7_75t_L g4543 ( 
.A(n_4280),
.B(n_232),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4318),
.Y(n_4544)
);

HB1xp67_ASAP7_75t_L g4545 ( 
.A(n_4400),
.Y(n_4545)
);

HB1xp67_ASAP7_75t_L g4546 ( 
.A(n_4406),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4326),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4278),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4319),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4432),
.B(n_232),
.Y(n_4550)
);

OR2x2_ASAP7_75t_L g4551 ( 
.A(n_4408),
.B(n_233),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4322),
.B(n_233),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_4245),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_SL g4554 ( 
.A(n_4260),
.B(n_234),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4247),
.Y(n_4555)
);

AND2x4_ASAP7_75t_L g4556 ( 
.A(n_4414),
.B(n_234),
.Y(n_4556)
);

OR2x2_ASAP7_75t_L g4557 ( 
.A(n_4410),
.B(n_235),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4332),
.B(n_236),
.Y(n_4558)
);

OR2x2_ASAP7_75t_L g4559 ( 
.A(n_4412),
.B(n_237),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_4418),
.B(n_237),
.Y(n_4560)
);

OR2x2_ASAP7_75t_L g4561 ( 
.A(n_4415),
.B(n_238),
.Y(n_4561)
);

OR2x2_ASAP7_75t_L g4562 ( 
.A(n_4431),
.B(n_4433),
.Y(n_4562)
);

AND2x2_ASAP7_75t_L g4563 ( 
.A(n_4323),
.B(n_239),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4306),
.B(n_240),
.Y(n_4564)
);

INVx1_ASAP7_75t_SL g4565 ( 
.A(n_4252),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4327),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4307),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4402),
.B(n_240),
.Y(n_4568)
);

HB1xp67_ASAP7_75t_L g4569 ( 
.A(n_4239),
.Y(n_4569)
);

OR2x2_ASAP7_75t_L g4570 ( 
.A(n_4411),
.B(n_241),
.Y(n_4570)
);

NOR2xp33_ASAP7_75t_L g4571 ( 
.A(n_4271),
.B(n_242),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4420),
.Y(n_4572)
);

HB1xp67_ASAP7_75t_L g4573 ( 
.A(n_4441),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4545),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4474),
.B(n_4380),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4531),
.B(n_4309),
.Y(n_4576)
);

BUFx3_ASAP7_75t_L g4577 ( 
.A(n_4511),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4461),
.B(n_4526),
.Y(n_4578)
);

OR2x2_ASAP7_75t_L g4579 ( 
.A(n_4541),
.B(n_4328),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4546),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4476),
.B(n_4311),
.Y(n_4581)
);

OR2x2_ASAP7_75t_L g4582 ( 
.A(n_4449),
.B(n_4525),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4436),
.Y(n_4583)
);

OR2x2_ASAP7_75t_L g4584 ( 
.A(n_4553),
.B(n_4421),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4447),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4495),
.Y(n_4586)
);

NOR2x1_ASAP7_75t_SL g4587 ( 
.A(n_4471),
.B(n_4262),
.Y(n_4587)
);

INVx4_ASAP7_75t_L g4588 ( 
.A(n_4445),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4442),
.B(n_4419),
.Y(n_4589)
);

OR2x2_ASAP7_75t_L g4590 ( 
.A(n_4555),
.B(n_4268),
.Y(n_4590)
);

BUFx2_ASAP7_75t_L g4591 ( 
.A(n_4500),
.Y(n_4591)
);

INVx4_ASAP7_75t_L g4592 ( 
.A(n_4477),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4479),
.B(n_4423),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4437),
.B(n_4430),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4446),
.B(n_4392),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4434),
.B(n_4304),
.Y(n_4596)
);

OR2x2_ASAP7_75t_L g4597 ( 
.A(n_4450),
.B(n_4292),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4456),
.B(n_4259),
.Y(n_4598)
);

AND2x4_ASAP7_75t_L g4599 ( 
.A(n_4448),
.B(n_4289),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4509),
.B(n_4336),
.Y(n_4600)
);

INVxp67_ASAP7_75t_SL g4601 ( 
.A(n_4497),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4565),
.B(n_4264),
.Y(n_4602)
);

AND2x4_ASAP7_75t_SL g4603 ( 
.A(n_4540),
.B(n_4556),
.Y(n_4603)
);

HB1xp67_ASAP7_75t_L g4604 ( 
.A(n_4569),
.Y(n_4604)
);

INVx4_ASAP7_75t_L g4605 ( 
.A(n_4508),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4452),
.Y(n_4606)
);

OR2x2_ASAP7_75t_L g4607 ( 
.A(n_4521),
.B(n_4297),
.Y(n_4607)
);

OR2x2_ASAP7_75t_L g4608 ( 
.A(n_4470),
.B(n_4387),
.Y(n_4608)
);

INVx2_ASAP7_75t_L g4609 ( 
.A(n_4538),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4485),
.B(n_4265),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4486),
.B(n_4272),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4443),
.B(n_4492),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4438),
.B(n_4369),
.Y(n_4613)
);

OR2x2_ASAP7_75t_L g4614 ( 
.A(n_4473),
.B(n_4324),
.Y(n_4614)
);

INVx2_ASAP7_75t_L g4615 ( 
.A(n_4484),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_SL g4616 ( 
.A(n_4467),
.B(n_4294),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4562),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4572),
.B(n_4279),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4515),
.Y(n_4619)
);

AND2x4_ASAP7_75t_L g4620 ( 
.A(n_4454),
.B(n_4462),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4566),
.B(n_4325),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4488),
.B(n_4379),
.Y(n_4622)
);

OR2x2_ASAP7_75t_L g4623 ( 
.A(n_4453),
.B(n_4285),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4490),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4520),
.Y(n_4625)
);

BUFx3_ASAP7_75t_L g4626 ( 
.A(n_4560),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_4548),
.B(n_4312),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4551),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4468),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4557),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4472),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4503),
.B(n_4284),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4458),
.B(n_4291),
.Y(n_4633)
);

OR2x2_ASAP7_75t_L g4634 ( 
.A(n_4463),
.B(n_4370),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4480),
.B(n_4308),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4501),
.B(n_4293),
.Y(n_4636)
);

AND2x4_ASAP7_75t_SL g4637 ( 
.A(n_4494),
.B(n_4365),
.Y(n_4637)
);

AND2x2_ASAP7_75t_L g4638 ( 
.A(n_4504),
.B(n_4355),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4451),
.B(n_4346),
.Y(n_4639)
);

AND2x4_ASAP7_75t_L g4640 ( 
.A(n_4464),
.B(n_4359),
.Y(n_4640)
);

OR2x2_ASAP7_75t_L g4641 ( 
.A(n_4455),
.B(n_4337),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4459),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4483),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4532),
.B(n_4356),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4558),
.B(n_4361),
.Y(n_4645)
);

OR2x2_ASAP7_75t_L g4646 ( 
.A(n_4435),
.B(n_4339),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4533),
.B(n_4363),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4559),
.Y(n_4648)
);

INVx4_ASAP7_75t_L g4649 ( 
.A(n_4535),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4537),
.B(n_4550),
.Y(n_4650)
);

INVx1_ASAP7_75t_SL g4651 ( 
.A(n_4539),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4561),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4564),
.B(n_4351),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_4543),
.Y(n_4654)
);

OR2x2_ASAP7_75t_L g4655 ( 
.A(n_4439),
.B(n_4329),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4513),
.B(n_4362),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_L g4657 ( 
.A(n_4530),
.B(n_4305),
.Y(n_4657)
);

AND2x4_ASAP7_75t_L g4658 ( 
.A(n_4457),
.B(n_4499),
.Y(n_4658)
);

HB1xp67_ASAP7_75t_L g4659 ( 
.A(n_4469),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_4498),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4552),
.B(n_4374),
.Y(n_4661)
);

OR2x2_ASAP7_75t_L g4662 ( 
.A(n_4493),
.B(n_4403),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_SL g4663 ( 
.A(n_4466),
.B(n_4377),
.Y(n_4663)
);

INVx4_ASAP7_75t_L g4664 ( 
.A(n_4563),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_SL g4665 ( 
.A(n_4528),
.B(n_4317),
.Y(n_4665)
);

HB1xp67_ASAP7_75t_L g4666 ( 
.A(n_4505),
.Y(n_4666)
);

AOI31xp33_ASAP7_75t_L g4667 ( 
.A1(n_4440),
.A2(n_4385),
.A3(n_244),
.B(n_242),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4640),
.B(n_4517),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4604),
.Y(n_4669)
);

NOR2xp33_ASAP7_75t_L g4670 ( 
.A(n_4605),
.B(n_4514),
.Y(n_4670)
);

HB1xp67_ASAP7_75t_L g4671 ( 
.A(n_4573),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4575),
.B(n_4567),
.Y(n_4672)
);

INVx1_ASAP7_75t_SL g4673 ( 
.A(n_4637),
.Y(n_4673)
);

AOI22xp5_ASAP7_75t_L g4674 ( 
.A1(n_4659),
.A2(n_4444),
.B1(n_4571),
.B2(n_4536),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4589),
.B(n_4549),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4601),
.B(n_4518),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4591),
.B(n_4527),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4666),
.Y(n_4678)
);

OR2x2_ASAP7_75t_L g4679 ( 
.A(n_4612),
.B(n_4491),
.Y(n_4679)
);

AND2x2_ASAP7_75t_L g4680 ( 
.A(n_4578),
.B(n_4506),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4602),
.B(n_4507),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4576),
.B(n_4510),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4649),
.B(n_4512),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4653),
.B(n_4554),
.Y(n_4684)
);

HB1xp67_ASAP7_75t_L g4685 ( 
.A(n_4626),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4654),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4650),
.B(n_4475),
.Y(n_4687)
);

OR2x2_ASAP7_75t_L g4688 ( 
.A(n_4581),
.B(n_4460),
.Y(n_4688)
);

AND2x4_ASAP7_75t_L g4689 ( 
.A(n_4588),
.B(n_4465),
.Y(n_4689)
);

OR2x2_ASAP7_75t_L g4690 ( 
.A(n_4651),
.B(n_4478),
.Y(n_4690)
);

OR2x2_ASAP7_75t_L g4691 ( 
.A(n_4608),
.B(n_4570),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4574),
.Y(n_4692)
);

OAI21xp5_ASAP7_75t_L g4693 ( 
.A1(n_4616),
.A2(n_4568),
.B(n_4482),
.Y(n_4693)
);

OAI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4662),
.A2(n_4586),
.B1(n_4667),
.B2(n_4633),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4580),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4594),
.B(n_4593),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4582),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4595),
.B(n_4481),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4617),
.Y(n_4699)
);

INVx2_ASAP7_75t_L g4700 ( 
.A(n_4577),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_4661),
.B(n_4487),
.Y(n_4701)
);

OR2x2_ASAP7_75t_L g4702 ( 
.A(n_4579),
.B(n_4489),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4613),
.B(n_4496),
.Y(n_4703)
);

AND2x4_ASAP7_75t_L g4704 ( 
.A(n_4592),
.B(n_4502),
.Y(n_4704)
);

NOR2x1_ASAP7_75t_L g4705 ( 
.A(n_4664),
.B(n_4529),
.Y(n_4705)
);

NOR2xp67_ASAP7_75t_L g4706 ( 
.A(n_4609),
.B(n_4516),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4634),
.Y(n_4707)
);

INVx3_ASAP7_75t_L g4708 ( 
.A(n_4603),
.Y(n_4708)
);

NAND2x1p5_ASAP7_75t_L g4709 ( 
.A(n_4620),
.B(n_4519),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_4599),
.Y(n_4710)
);

INVxp67_ASAP7_75t_L g4711 ( 
.A(n_4587),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4644),
.B(n_4522),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4596),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4619),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4647),
.B(n_4523),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4598),
.Y(n_4716)
);

AND2x2_ASAP7_75t_L g4717 ( 
.A(n_4645),
.B(n_4524),
.Y(n_4717)
);

INVx1_ASAP7_75t_SL g4718 ( 
.A(n_4638),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4632),
.B(n_4534),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4625),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4636),
.B(n_4542),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4623),
.Y(n_4722)
);

AND2x4_ASAP7_75t_L g4723 ( 
.A(n_4600),
.B(n_4544),
.Y(n_4723)
);

OR2x2_ASAP7_75t_L g4724 ( 
.A(n_4655),
.B(n_4547),
.Y(n_4724)
);

OR2x2_ASAP7_75t_L g4725 ( 
.A(n_4641),
.B(n_243),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4658),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4618),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4610),
.B(n_243),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4657),
.B(n_244),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4709),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4708),
.B(n_4611),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4671),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4696),
.B(n_4673),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4685),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4669),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4700),
.B(n_4606),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4686),
.Y(n_4737)
);

A2O1A1Ixp33_ASAP7_75t_L g4738 ( 
.A1(n_4674),
.A2(n_4665),
.B(n_4583),
.C(n_4639),
.Y(n_4738)
);

INVx2_ASAP7_75t_L g4739 ( 
.A(n_4668),
.Y(n_4739)
);

AOI21xp5_ASAP7_75t_L g4740 ( 
.A1(n_4711),
.A2(n_4622),
.B(n_4663),
.Y(n_4740)
);

AND2x4_ASAP7_75t_L g4741 ( 
.A(n_4710),
.B(n_4629),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4726),
.Y(n_4742)
);

OR2x2_ASAP7_75t_L g4743 ( 
.A(n_4718),
.B(n_4631),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4672),
.B(n_4660),
.Y(n_4744)
);

NOR2x1_ASAP7_75t_L g4745 ( 
.A(n_4705),
.B(n_4628),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4675),
.B(n_4643),
.Y(n_4746)
);

AOI22xp5_ASAP7_75t_L g4747 ( 
.A1(n_4694),
.A2(n_4648),
.B1(n_4652),
.B2(n_4630),
.Y(n_4747)
);

NAND2x1p5_ASAP7_75t_L g4748 ( 
.A(n_4704),
.B(n_4615),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4706),
.B(n_4624),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4728),
.B(n_4642),
.Y(n_4750)
);

AND2x4_ASAP7_75t_L g4751 ( 
.A(n_4727),
.B(n_4656),
.Y(n_4751)
);

INVx1_ASAP7_75t_SL g4752 ( 
.A(n_4691),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4684),
.B(n_4607),
.Y(n_4753)
);

INVx2_ASAP7_75t_L g4754 ( 
.A(n_4713),
.Y(n_4754)
);

OR2x2_ASAP7_75t_L g4755 ( 
.A(n_4678),
.B(n_4627),
.Y(n_4755)
);

OR2x2_ASAP7_75t_L g4756 ( 
.A(n_4716),
.B(n_4584),
.Y(n_4756)
);

INVxp67_ASAP7_75t_L g4757 ( 
.A(n_4670),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4681),
.B(n_4635),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4719),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4721),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4715),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4717),
.Y(n_4762)
);

NOR2xp33_ASAP7_75t_L g4763 ( 
.A(n_4682),
.B(n_4646),
.Y(n_4763)
);

INVx2_ASAP7_75t_SL g4764 ( 
.A(n_4723),
.Y(n_4764)
);

AOI21xp33_ASAP7_75t_SL g4765 ( 
.A1(n_4722),
.A2(n_4614),
.B(n_4597),
.Y(n_4765)
);

INVx2_ASAP7_75t_L g4766 ( 
.A(n_4689),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4680),
.B(n_4585),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4687),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4698),
.B(n_4590),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4707),
.B(n_4621),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4724),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4697),
.B(n_245),
.Y(n_4772)
);

NOR2xp33_ASAP7_75t_L g4773 ( 
.A(n_4677),
.B(n_245),
.Y(n_4773)
);

OR2x2_ASAP7_75t_L g4774 ( 
.A(n_4702),
.B(n_247),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4701),
.Y(n_4775)
);

NOR3xp33_ASAP7_75t_L g4776 ( 
.A(n_4676),
.B(n_248),
.C(n_249),
.Y(n_4776)
);

OAI22xp33_ASAP7_75t_L g4777 ( 
.A1(n_4752),
.A2(n_4693),
.B1(n_4690),
.B2(n_4683),
.Y(n_4777)
);

INVxp67_ASAP7_75t_SL g4778 ( 
.A(n_4748),
.Y(n_4778)
);

AOI22xp5_ASAP7_75t_L g4779 ( 
.A1(n_4733),
.A2(n_4695),
.B1(n_4692),
.B2(n_4699),
.Y(n_4779)
);

AOI31xp33_ASAP7_75t_L g4780 ( 
.A1(n_4745),
.A2(n_4714),
.A3(n_4720),
.B(n_4679),
.Y(n_4780)
);

NAND3xp33_ASAP7_75t_L g4781 ( 
.A(n_4738),
.B(n_4703),
.C(n_4688),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4731),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4744),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4764),
.B(n_4739),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4734),
.Y(n_4785)
);

OAI22xp5_ASAP7_75t_L g4786 ( 
.A1(n_4747),
.A2(n_4712),
.B1(n_4729),
.B2(n_4725),
.Y(n_4786)
);

OAI31xp33_ASAP7_75t_L g4787 ( 
.A1(n_4776),
.A2(n_253),
.A3(n_250),
.B(n_252),
.Y(n_4787)
);

AOI211xp5_ASAP7_75t_SL g4788 ( 
.A1(n_4740),
.A2(n_259),
.B(n_267),
.C(n_250),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4746),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4755),
.Y(n_4790)
);

NOR2xp33_ASAP7_75t_SL g4791 ( 
.A(n_4730),
.B(n_253),
.Y(n_4791)
);

OA21x2_ASAP7_75t_L g4792 ( 
.A1(n_4749),
.A2(n_252),
.B(n_254),
.Y(n_4792)
);

AOI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_4758),
.A2(n_255),
.B(n_256),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4743),
.Y(n_4794)
);

AO22x1_ASAP7_75t_L g4795 ( 
.A1(n_4732),
.A2(n_263),
.B1(n_275),
.B2(n_255),
.Y(n_4795)
);

XNOR2xp5_ASAP7_75t_L g4796 ( 
.A(n_4751),
.B(n_256),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4741),
.B(n_257),
.Y(n_4797)
);

AOI22xp33_ASAP7_75t_L g4798 ( 
.A1(n_4742),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4770),
.A2(n_258),
.B(n_261),
.Y(n_4799)
);

A2O1A1Ixp33_ASAP7_75t_L g4800 ( 
.A1(n_4773),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4769),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4756),
.Y(n_4802)
);

NAND4xp25_ASAP7_75t_L g4803 ( 
.A(n_4763),
.B(n_265),
.C(n_262),
.D(n_264),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4759),
.Y(n_4804)
);

BUFx2_ASAP7_75t_SL g4805 ( 
.A(n_4766),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4760),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_4750),
.A2(n_265),
.B(n_266),
.Y(n_4807)
);

XOR2x2_ASAP7_75t_L g4808 ( 
.A(n_4753),
.B(n_268),
.Y(n_4808)
);

XNOR2x1_ASAP7_75t_L g4809 ( 
.A(n_4736),
.B(n_269),
.Y(n_4809)
);

INVxp67_ASAP7_75t_L g4810 ( 
.A(n_4761),
.Y(n_4810)
);

INVx1_ASAP7_75t_SL g4811 ( 
.A(n_4774),
.Y(n_4811)
);

AOI31xp33_ASAP7_75t_L g4812 ( 
.A1(n_4757),
.A2(n_274),
.A3(n_269),
.B(n_271),
.Y(n_4812)
);

OA22x2_ASAP7_75t_L g4813 ( 
.A1(n_4762),
.A2(n_276),
.B1(n_271),
.B2(n_274),
.Y(n_4813)
);

OAI22xp33_ASAP7_75t_L g4814 ( 
.A1(n_4771),
.A2(n_4767),
.B1(n_4754),
.B2(n_4737),
.Y(n_4814)
);

AOI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4775),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_4815)
);

OAI21xp33_ASAP7_75t_L g4816 ( 
.A1(n_4735),
.A2(n_277),
.B(n_280),
.Y(n_4816)
);

INVxp67_ASAP7_75t_SL g4817 ( 
.A(n_4772),
.Y(n_4817)
);

XOR2x2_ASAP7_75t_L g4818 ( 
.A(n_4768),
.B(n_280),
.Y(n_4818)
);

OAI21xp5_ASAP7_75t_L g4819 ( 
.A1(n_4765),
.A2(n_285),
.B(n_284),
.Y(n_4819)
);

AOI21xp33_ASAP7_75t_L g4820 ( 
.A1(n_4745),
.A2(n_282),
.B(n_284),
.Y(n_4820)
);

AOI21x1_ASAP7_75t_L g4821 ( 
.A1(n_4745),
.A2(n_285),
.B(n_286),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4744),
.Y(n_4822)
);

NOR2xp33_ASAP7_75t_L g4823 ( 
.A(n_4733),
.B(n_288),
.Y(n_4823)
);

NOR2xp67_ASAP7_75t_L g4824 ( 
.A(n_4764),
.B(n_289),
.Y(n_4824)
);

NAND2x1p5_ASAP7_75t_L g4825 ( 
.A(n_4733),
.B(n_290),
.Y(n_4825)
);

XNOR2xp5_ASAP7_75t_L g4826 ( 
.A(n_4733),
.B(n_289),
.Y(n_4826)
);

AOI22x1_ASAP7_75t_L g4827 ( 
.A1(n_4778),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_4827)
);

AOI21xp5_ASAP7_75t_L g4828 ( 
.A1(n_4780),
.A2(n_291),
.B(n_292),
.Y(n_4828)
);

INVx1_ASAP7_75t_SL g4829 ( 
.A(n_4805),
.Y(n_4829)
);

OAI32xp33_ASAP7_75t_L g4830 ( 
.A1(n_4781),
.A2(n_295),
.A3(n_297),
.B1(n_294),
.B2(n_296),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_4825),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4782),
.Y(n_4832)
);

INVxp67_ASAP7_75t_L g4833 ( 
.A(n_4824),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4821),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4795),
.B(n_293),
.Y(n_4835)
);

AOI32xp33_ASAP7_75t_L g4836 ( 
.A1(n_4777),
.A2(n_4788),
.A3(n_4814),
.B1(n_4801),
.B2(n_4789),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4796),
.Y(n_4837)
);

INVxp67_ASAP7_75t_L g4838 ( 
.A(n_4791),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4826),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4784),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4783),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4822),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4817),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4790),
.B(n_293),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4792),
.Y(n_4845)
);

NAND2x1_ASAP7_75t_L g4846 ( 
.A(n_4792),
.B(n_294),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4797),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4802),
.B(n_4794),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4813),
.Y(n_4849)
);

AOI22xp5_ASAP7_75t_L g4850 ( 
.A1(n_4786),
.A2(n_298),
.B1(n_295),
.B2(n_296),
.Y(n_4850)
);

AOI32xp33_ASAP7_75t_L g4851 ( 
.A1(n_4785),
.A2(n_300),
.A3(n_298),
.B1(n_299),
.B2(n_302),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4779),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4809),
.Y(n_4853)
);

OAI21xp33_ASAP7_75t_SL g4854 ( 
.A1(n_4820),
.A2(n_303),
.B(n_304),
.Y(n_4854)
);

INVx2_ASAP7_75t_SL g4855 ( 
.A(n_4808),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4823),
.Y(n_4856)
);

O2A1O1Ixp33_ASAP7_75t_L g4857 ( 
.A1(n_4819),
.A2(n_307),
.B(n_303),
.C(n_306),
.Y(n_4857)
);

NOR2xp33_ASAP7_75t_L g4858 ( 
.A(n_4811),
.B(n_307),
.Y(n_4858)
);

INVxp67_ASAP7_75t_SL g4859 ( 
.A(n_4818),
.Y(n_4859)
);

NOR2xp33_ASAP7_75t_L g4860 ( 
.A(n_4803),
.B(n_308),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4793),
.B(n_308),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4816),
.B(n_309),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4804),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4806),
.Y(n_4864)
);

OAI21xp33_ASAP7_75t_L g4865 ( 
.A1(n_4810),
.A2(n_310),
.B(n_311),
.Y(n_4865)
);

OAI33xp33_ASAP7_75t_L g4866 ( 
.A1(n_4787),
.A2(n_312),
.A3(n_315),
.B1(n_310),
.B2(n_311),
.B3(n_313),
.Y(n_4866)
);

AND2x2_ASAP7_75t_L g4867 ( 
.A(n_4807),
.B(n_312),
.Y(n_4867)
);

OAI222xp33_ASAP7_75t_L g4868 ( 
.A1(n_4799),
.A2(n_318),
.B1(n_320),
.B2(n_313),
.C1(n_315),
.C2(n_319),
.Y(n_4868)
);

OAI21xp5_ASAP7_75t_SL g4869 ( 
.A1(n_4812),
.A2(n_318),
.B(n_319),
.Y(n_4869)
);

OAI22xp5_ASAP7_75t_L g4870 ( 
.A1(n_4798),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_4870)
);

AND2x2_ASAP7_75t_L g4871 ( 
.A(n_4800),
.B(n_321),
.Y(n_4871)
);

OR2x2_ASAP7_75t_L g4872 ( 
.A(n_4815),
.B(n_322),
.Y(n_4872)
);

NOR2xp33_ASAP7_75t_L g4873 ( 
.A(n_4778),
.B(n_323),
.Y(n_4873)
);

AND2x2_ASAP7_75t_L g4874 ( 
.A(n_4778),
.B(n_324),
.Y(n_4874)
);

INVx3_ASAP7_75t_L g4875 ( 
.A(n_4825),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4824),
.Y(n_4876)
);

O2A1O1Ixp5_ASAP7_75t_L g4877 ( 
.A1(n_4778),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4824),
.B(n_325),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4824),
.Y(n_4879)
);

INVx1_ASAP7_75t_SL g4880 ( 
.A(n_4805),
.Y(n_4880)
);

OR2x2_ASAP7_75t_L g4881 ( 
.A(n_4782),
.B(n_326),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4778),
.B(n_327),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4824),
.B(n_328),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4829),
.B(n_4880),
.Y(n_4884)
);

OR2x2_ASAP7_75t_L g4885 ( 
.A(n_4876),
.B(n_328),
.Y(n_4885)
);

INVxp67_ASAP7_75t_SL g4886 ( 
.A(n_4846),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4833),
.B(n_329),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4845),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4879),
.B(n_329),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4848),
.B(n_331),
.Y(n_4890)
);

O2A1O1Ixp33_ASAP7_75t_L g4891 ( 
.A1(n_4830),
.A2(n_341),
.B(n_352),
.C(n_332),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4849),
.B(n_332),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4874),
.Y(n_4893)
);

AND2x2_ASAP7_75t_L g4894 ( 
.A(n_4831),
.B(n_333),
.Y(n_4894)
);

OAI31xp33_ASAP7_75t_L g4895 ( 
.A1(n_4868),
.A2(n_4828),
.A3(n_4869),
.B(n_4852),
.Y(n_4895)
);

INVx2_ASAP7_75t_SL g4896 ( 
.A(n_4875),
.Y(n_4896)
);

AOI211xp5_ASAP7_75t_L g4897 ( 
.A1(n_4854),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4882),
.Y(n_4898)
);

AOI22xp5_ASAP7_75t_L g4899 ( 
.A1(n_4855),
.A2(n_338),
.B1(n_334),
.B2(n_337),
.Y(n_4899)
);

HB1xp67_ASAP7_75t_L g4900 ( 
.A(n_4875),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4834),
.B(n_337),
.Y(n_4901)
);

NOR3xp33_ASAP7_75t_L g4902 ( 
.A(n_4859),
.B(n_349),
.C(n_338),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4827),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4836),
.B(n_339),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4878),
.Y(n_4905)
);

NAND3xp33_ASAP7_75t_SL g4906 ( 
.A(n_4877),
.B(n_339),
.C(n_340),
.Y(n_4906)
);

OAI221xp5_ASAP7_75t_L g4907 ( 
.A1(n_4838),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.C(n_345),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4873),
.B(n_342),
.Y(n_4908)
);

AOI22xp5_ASAP7_75t_L g4909 ( 
.A1(n_4840),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_SL g4910 ( 
.A1(n_4843),
.A2(n_350),
.B1(n_346),
.B2(n_348),
.Y(n_4910)
);

OAI22xp5_ASAP7_75t_L g4911 ( 
.A1(n_4832),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_4911)
);

NOR2xp33_ASAP7_75t_L g4912 ( 
.A(n_4866),
.B(n_351),
.Y(n_4912)
);

OAI21xp5_ASAP7_75t_SL g4913 ( 
.A1(n_4853),
.A2(n_353),
.B(n_355),
.Y(n_4913)
);

OAI322xp33_ASAP7_75t_L g4914 ( 
.A1(n_4841),
.A2(n_360),
.A3(n_359),
.B1(n_357),
.B2(n_355),
.C1(n_356),
.C2(n_358),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4883),
.Y(n_4915)
);

AOI21xp5_ASAP7_75t_L g4916 ( 
.A1(n_4861),
.A2(n_357),
.B(n_360),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4844),
.B(n_361),
.Y(n_4917)
);

INVx2_ASAP7_75t_SL g4918 ( 
.A(n_4881),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4839),
.B(n_361),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4835),
.Y(n_4920)
);

INVx1_ASAP7_75t_L g4921 ( 
.A(n_4858),
.Y(n_4921)
);

NOR2xp33_ASAP7_75t_L g4922 ( 
.A(n_4865),
.B(n_362),
.Y(n_4922)
);

AND2x2_ASAP7_75t_L g4923 ( 
.A(n_4837),
.B(n_362),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4842),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4863),
.Y(n_4925)
);

NOR2xp33_ASAP7_75t_L g4926 ( 
.A(n_4860),
.B(n_363),
.Y(n_4926)
);

OAI22xp33_ASAP7_75t_L g4927 ( 
.A1(n_4850),
.A2(n_4872),
.B1(n_4856),
.B2(n_4864),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_4867),
.B(n_363),
.Y(n_4928)
);

AOI21xp5_ASAP7_75t_L g4929 ( 
.A1(n_4857),
.A2(n_364),
.B(n_365),
.Y(n_4929)
);

INVx1_ASAP7_75t_SL g4930 ( 
.A(n_4871),
.Y(n_4930)
);

OAI22xp33_ASAP7_75t_SL g4931 ( 
.A1(n_4847),
.A2(n_367),
.B1(n_364),
.B2(n_365),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4862),
.Y(n_4932)
);

AOI211xp5_ASAP7_75t_L g4933 ( 
.A1(n_4870),
.A2(n_4851),
.B(n_369),
.C(n_367),
.Y(n_4933)
);

OAI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4829),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_4934)
);

AOI21xp33_ASAP7_75t_L g4935 ( 
.A1(n_4829),
.A2(n_371),
.B(n_370),
.Y(n_4935)
);

AOI221xp5_ASAP7_75t_L g4936 ( 
.A1(n_4828),
.A2(n_375),
.B1(n_378),
.B2(n_374),
.C(n_377),
.Y(n_4936)
);

OAI21xp5_ASAP7_75t_SL g4937 ( 
.A1(n_4829),
.A2(n_368),
.B(n_374),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4829),
.B(n_375),
.Y(n_4938)
);

OR2x2_ASAP7_75t_L g4939 ( 
.A(n_4829),
.B(n_377),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4846),
.Y(n_4940)
);

AND2x2_ASAP7_75t_SL g4941 ( 
.A(n_4876),
.B(n_378),
.Y(n_4941)
);

NOR2xp33_ASAP7_75t_L g4942 ( 
.A(n_4829),
.B(n_379),
.Y(n_4942)
);

OAI222xp33_ASAP7_75t_L g4943 ( 
.A1(n_4829),
.A2(n_381),
.B1(n_383),
.B2(n_379),
.C1(n_380),
.C2(n_382),
.Y(n_4943)
);

AOI21xp33_ASAP7_75t_SL g4944 ( 
.A1(n_4833),
.A2(n_383),
.B(n_382),
.Y(n_4944)
);

NOR3xp33_ASAP7_75t_L g4945 ( 
.A(n_4875),
.B(n_393),
.C(n_380),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4846),
.Y(n_4946)
);

O2A1O1Ixp33_ASAP7_75t_L g4947 ( 
.A1(n_4830),
.A2(n_397),
.B(n_405),
.C(n_384),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4846),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4829),
.B(n_385),
.Y(n_4949)
);

XNOR2x2_ASAP7_75t_L g4950 ( 
.A(n_4828),
.B(n_385),
.Y(n_4950)
);

OAI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4833),
.A2(n_386),
.B(n_389),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4846),
.Y(n_4952)
);

AOI222xp33_ASAP7_75t_L g4953 ( 
.A1(n_4852),
.A2(n_390),
.B1(n_392),
.B2(n_386),
.C1(n_389),
.C2(n_391),
.Y(n_4953)
);

INVx2_ASAP7_75t_L g4954 ( 
.A(n_4875),
.Y(n_4954)
);

O2A1O1Ixp33_ASAP7_75t_L g4955 ( 
.A1(n_4830),
.A2(n_401),
.B(n_409),
.C(n_390),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4846),
.Y(n_4956)
);

NOR2x1_ASAP7_75t_L g4957 ( 
.A(n_4845),
.B(n_391),
.Y(n_4957)
);

A2O1A1Ixp33_ASAP7_75t_L g4958 ( 
.A1(n_4828),
.A2(n_397),
.B(n_398),
.C(n_393),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4875),
.Y(n_4959)
);

NOR2x1_ASAP7_75t_L g4960 ( 
.A(n_4845),
.B(n_392),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4829),
.B(n_399),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4875),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4875),
.Y(n_4963)
);

AOI22xp33_ASAP7_75t_L g4964 ( 
.A1(n_4852),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_4964)
);

NAND2xp5_ASAP7_75t_L g4965 ( 
.A(n_4829),
.B(n_400),
.Y(n_4965)
);

OAI21xp33_ASAP7_75t_L g4966 ( 
.A1(n_4836),
.A2(n_410),
.B(n_402),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4846),
.Y(n_4967)
);

O2A1O1Ixp33_ASAP7_75t_L g4968 ( 
.A1(n_4830),
.A2(n_413),
.B(n_421),
.C(n_403),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4829),
.B(n_403),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4846),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4886),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4957),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4960),
.Y(n_4973)
);

NOR2x1_ASAP7_75t_L g4974 ( 
.A(n_4940),
.B(n_404),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_SL g4975 ( 
.A(n_4946),
.B(n_405),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4900),
.Y(n_4976)
);

AOI221xp5_ASAP7_75t_SL g4977 ( 
.A1(n_4966),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.C(n_409),
.Y(n_4977)
);

NOR3xp33_ASAP7_75t_SL g4978 ( 
.A(n_4927),
.B(n_406),
.C(n_407),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4948),
.B(n_408),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4884),
.A2(n_4956),
.B(n_4952),
.Y(n_4980)
);

OAI21xp5_ASAP7_75t_L g4981 ( 
.A1(n_4891),
.A2(n_4955),
.B(n_4947),
.Y(n_4981)
);

O2A1O1Ixp5_ASAP7_75t_SL g4982 ( 
.A1(n_4888),
.A2(n_414),
.B(n_411),
.C(n_413),
.Y(n_4982)
);

OR2x2_ASAP7_75t_L g4983 ( 
.A(n_4967),
.B(n_414),
.Y(n_4983)
);

NOR2xp33_ASAP7_75t_L g4984 ( 
.A(n_4970),
.B(n_415),
.Y(n_4984)
);

NOR2xp33_ASAP7_75t_L g4985 ( 
.A(n_4893),
.B(n_415),
.Y(n_4985)
);

OAI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4968),
.A2(n_4929),
.B(n_4942),
.Y(n_4986)
);

NOR3xp33_ASAP7_75t_L g4987 ( 
.A(n_4896),
.B(n_416),
.C(n_417),
.Y(n_4987)
);

NAND3xp33_ASAP7_75t_L g4988 ( 
.A(n_4897),
.B(n_416),
.C(n_418),
.Y(n_4988)
);

BUFx2_ASAP7_75t_L g4989 ( 
.A(n_4941),
.Y(n_4989)
);

XNOR2x1_ASAP7_75t_L g4990 ( 
.A(n_4950),
.B(n_4939),
.Y(n_4990)
);

NAND3xp33_ASAP7_75t_L g4991 ( 
.A(n_4895),
.B(n_419),
.C(n_420),
.Y(n_4991)
);

NOR2xp33_ASAP7_75t_L g4992 ( 
.A(n_4898),
.B(n_420),
.Y(n_4992)
);

NAND3xp33_ASAP7_75t_SL g4993 ( 
.A(n_4933),
.B(n_421),
.C(n_422),
.Y(n_4993)
);

OR2x2_ASAP7_75t_L g4994 ( 
.A(n_4906),
.B(n_422),
.Y(n_4994)
);

INVxp33_ASAP7_75t_L g4995 ( 
.A(n_4892),
.Y(n_4995)
);

AOI221xp5_ASAP7_75t_L g4996 ( 
.A1(n_4904),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.C(n_427),
.Y(n_4996)
);

OAI21xp5_ASAP7_75t_SL g4997 ( 
.A1(n_4937),
.A2(n_4903),
.B(n_4912),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4890),
.B(n_423),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4885),
.Y(n_4999)
);

NOR2xp33_ASAP7_75t_L g5000 ( 
.A(n_4954),
.B(n_424),
.Y(n_5000)
);

OAI221xp5_ASAP7_75t_SL g5001 ( 
.A1(n_4959),
.A2(n_428),
.B1(n_425),
.B2(n_427),
.C(n_429),
.Y(n_5001)
);

AOI221xp5_ASAP7_75t_SL g5002 ( 
.A1(n_4930),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.C(n_432),
.Y(n_5002)
);

NAND2x1_ASAP7_75t_L g5003 ( 
.A(n_4962),
.B(n_430),
.Y(n_5003)
);

INVxp67_ASAP7_75t_L g5004 ( 
.A(n_4938),
.Y(n_5004)
);

AOI21xp33_ASAP7_75t_SL g5005 ( 
.A1(n_4918),
.A2(n_432),
.B(n_434),
.Y(n_5005)
);

INVxp67_ASAP7_75t_L g5006 ( 
.A(n_4949),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4963),
.B(n_435),
.Y(n_5007)
);

NOR2xp33_ASAP7_75t_L g5008 ( 
.A(n_4913),
.B(n_435),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_SL g5009 ( 
.A(n_4931),
.B(n_436),
.Y(n_5009)
);

NAND2xp5_ASAP7_75t_L g5010 ( 
.A(n_4910),
.B(n_437),
.Y(n_5010)
);

NOR2xp33_ASAP7_75t_L g5011 ( 
.A(n_4944),
.B(n_437),
.Y(n_5011)
);

INVx2_ASAP7_75t_L g5012 ( 
.A(n_4894),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4961),
.Y(n_5013)
);

OAI322xp33_ASAP7_75t_L g5014 ( 
.A1(n_4924),
.A2(n_444),
.A3(n_443),
.B1(n_441),
.B2(n_439),
.C1(n_440),
.C2(n_442),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4919),
.B(n_439),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4953),
.B(n_441),
.Y(n_5016)
);

AOI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_4928),
.A2(n_442),
.B(n_444),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4965),
.Y(n_5018)
);

NOR2xp33_ASAP7_75t_L g5019 ( 
.A(n_4969),
.B(n_445),
.Y(n_5019)
);

AND2x2_ASAP7_75t_L g5020 ( 
.A(n_4923),
.B(n_4920),
.Y(n_5020)
);

AND2x2_ASAP7_75t_L g5021 ( 
.A(n_4902),
.B(n_446),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_SL g5022 ( 
.A(n_4936),
.B(n_447),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4921),
.B(n_447),
.Y(n_5023)
);

OR2x2_ASAP7_75t_L g5024 ( 
.A(n_4887),
.B(n_448),
.Y(n_5024)
);

INVx2_ASAP7_75t_L g5025 ( 
.A(n_4917),
.Y(n_5025)
);

AOI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_4916),
.A2(n_448),
.B(n_449),
.Y(n_5026)
);

AOI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4901),
.A2(n_449),
.B(n_450),
.Y(n_5027)
);

AOI21xp5_ASAP7_75t_L g5028 ( 
.A1(n_4889),
.A2(n_4958),
.B(n_4951),
.Y(n_5028)
);

NOR2xp33_ASAP7_75t_L g5029 ( 
.A(n_4935),
.B(n_451),
.Y(n_5029)
);

NAND3xp33_ASAP7_75t_L g5030 ( 
.A(n_4925),
.B(n_452),
.C(n_453),
.Y(n_5030)
);

AOI221xp5_ASAP7_75t_L g5031 ( 
.A1(n_4932),
.A2(n_4915),
.B1(n_4905),
.B2(n_4943),
.C(n_4914),
.Y(n_5031)
);

NOR2xp33_ASAP7_75t_L g5032 ( 
.A(n_4907),
.B(n_453),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4926),
.B(n_454),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_SL g5034 ( 
.A(n_4945),
.B(n_454),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_SL g5035 ( 
.A(n_4899),
.B(n_4934),
.Y(n_5035)
);

AOI21xp5_ASAP7_75t_L g5036 ( 
.A1(n_4908),
.A2(n_4922),
.B(n_4911),
.Y(n_5036)
);

NOR2x1_ASAP7_75t_L g5037 ( 
.A(n_4964),
.B(n_455),
.Y(n_5037)
);

INVxp67_ASAP7_75t_L g5038 ( 
.A(n_4909),
.Y(n_5038)
);

NOR3xp33_ASAP7_75t_L g5039 ( 
.A(n_4884),
.B(n_456),
.C(n_457),
.Y(n_5039)
);

NOR2xp33_ASAP7_75t_L g5040 ( 
.A(n_4886),
.B(n_456),
.Y(n_5040)
);

NOR2xp67_ASAP7_75t_L g5041 ( 
.A(n_4940),
.B(n_459),
.Y(n_5041)
);

NOR2xp33_ASAP7_75t_L g5042 ( 
.A(n_4886),
.B(n_459),
.Y(n_5042)
);

NAND3xp33_ASAP7_75t_SL g5043 ( 
.A(n_4897),
.B(n_460),
.C(n_461),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4886),
.B(n_460),
.Y(n_5044)
);

NOR2xp33_ASAP7_75t_L g5045 ( 
.A(n_4886),
.B(n_462),
.Y(n_5045)
);

INVxp67_ASAP7_75t_L g5046 ( 
.A(n_4886),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4886),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4886),
.Y(n_5048)
);

NAND3xp33_ASAP7_75t_SL g5049 ( 
.A(n_4897),
.B(n_464),
.C(n_465),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4886),
.B(n_464),
.Y(n_5050)
);

OAI21xp33_ASAP7_75t_L g5051 ( 
.A1(n_4966),
.A2(n_465),
.B(n_466),
.Y(n_5051)
);

O2A1O1Ixp33_ASAP7_75t_L g5052 ( 
.A1(n_4943),
.A2(n_468),
.B(n_466),
.C(n_467),
.Y(n_5052)
);

NAND3xp33_ASAP7_75t_L g5053 ( 
.A(n_4897),
.B(n_469),
.C(n_470),
.Y(n_5053)
);

INVx1_ASAP7_75t_SL g5054 ( 
.A(n_4941),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4886),
.B(n_469),
.Y(n_5055)
);

OAI211xp5_ASAP7_75t_L g5056 ( 
.A1(n_4980),
.A2(n_5046),
.B(n_4997),
.C(n_5031),
.Y(n_5056)
);

A2O1A1Ixp33_ASAP7_75t_L g5057 ( 
.A1(n_5052),
.A2(n_474),
.B(n_471),
.C(n_472),
.Y(n_5057)
);

O2A1O1Ixp33_ASAP7_75t_SL g5058 ( 
.A1(n_4972),
.A2(n_481),
.B(n_489),
.C(n_471),
.Y(n_5058)
);

NAND3xp33_ASAP7_75t_SL g5059 ( 
.A(n_5054),
.B(n_472),
.C(n_475),
.Y(n_5059)
);

NOR3xp33_ASAP7_75t_L g5060 ( 
.A(n_4991),
.B(n_4993),
.C(n_4989),
.Y(n_5060)
);

AOI211xp5_ASAP7_75t_L g5061 ( 
.A1(n_4976),
.A2(n_477),
.B(n_475),
.C(n_476),
.Y(n_5061)
);

AOI222xp33_ASAP7_75t_L g5062 ( 
.A1(n_4971),
.A2(n_479),
.B1(n_482),
.B2(n_477),
.C1(n_478),
.C2(n_480),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_5041),
.B(n_5047),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_5048),
.B(n_478),
.Y(n_5064)
);

OAI21xp5_ASAP7_75t_SL g5065 ( 
.A1(n_4995),
.A2(n_479),
.B(n_480),
.Y(n_5065)
);

AOI22xp5_ASAP7_75t_L g5066 ( 
.A1(n_5051),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_5066)
);

AOI221xp5_ASAP7_75t_L g5067 ( 
.A1(n_5040),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.C(n_487),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_5042),
.B(n_485),
.Y(n_5068)
);

NAND4xp25_ASAP7_75t_L g5069 ( 
.A(n_4981),
.B(n_489),
.C(n_487),
.D(n_488),
.Y(n_5069)
);

AOI22xp33_ASAP7_75t_L g5070 ( 
.A1(n_5043),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_5070)
);

AO22x2_ASAP7_75t_L g5071 ( 
.A1(n_4973),
.A2(n_494),
.B1(n_490),
.B2(n_493),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_5045),
.B(n_493),
.Y(n_5072)
);

OAI21xp5_ASAP7_75t_L g5073 ( 
.A1(n_4988),
.A2(n_497),
.B(n_496),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_4983),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_L g5075 ( 
.A(n_5015),
.B(n_495),
.Y(n_5075)
);

NAND3xp33_ASAP7_75t_SL g5076 ( 
.A(n_5003),
.B(n_498),
.C(n_499),
.Y(n_5076)
);

AOI211xp5_ASAP7_75t_L g5077 ( 
.A1(n_5049),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_5077)
);

NOR2xp33_ASAP7_75t_L g5078 ( 
.A(n_4994),
.B(n_501),
.Y(n_5078)
);

AOI221xp5_ASAP7_75t_L g5079 ( 
.A1(n_5038),
.A2(n_505),
.B1(n_502),
.B2(n_503),
.C(n_506),
.Y(n_5079)
);

OAI21xp33_ASAP7_75t_L g5080 ( 
.A1(n_4990),
.A2(n_4978),
.B(n_5035),
.Y(n_5080)
);

AOI22xp5_ASAP7_75t_L g5081 ( 
.A1(n_4987),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_5081)
);

A2O1A1Ixp33_ASAP7_75t_L g5082 ( 
.A1(n_4984),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_5002),
.B(n_508),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_L g5084 ( 
.A(n_5005),
.B(n_509),
.Y(n_5084)
);

AOI221xp5_ASAP7_75t_L g5085 ( 
.A1(n_4986),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.C(n_513),
.Y(n_5085)
);

NAND4xp25_ASAP7_75t_SL g5086 ( 
.A(n_4977),
.B(n_515),
.C(n_510),
.D(n_514),
.Y(n_5086)
);

OAI21xp5_ASAP7_75t_L g5087 ( 
.A1(n_5053),
.A2(n_518),
.B(n_517),
.Y(n_5087)
);

AOI211xp5_ASAP7_75t_L g5088 ( 
.A1(n_5009),
.A2(n_518),
.B(n_515),
.C(n_517),
.Y(n_5088)
);

NOR2x1_ASAP7_75t_L g5089 ( 
.A(n_4974),
.B(n_519),
.Y(n_5089)
);

OAI22xp5_ASAP7_75t_L g5090 ( 
.A1(n_5010),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_5090)
);

AOI22xp5_ASAP7_75t_L g5091 ( 
.A1(n_5032),
.A2(n_523),
.B1(n_520),
.B2(n_522),
.Y(n_5091)
);

NOR2xp33_ASAP7_75t_L g5092 ( 
.A(n_4998),
.B(n_522),
.Y(n_5092)
);

AOI21xp5_ASAP7_75t_L g5093 ( 
.A1(n_4975),
.A2(n_524),
.B(n_525),
.Y(n_5093)
);

NOR3xp33_ASAP7_75t_L g5094 ( 
.A(n_5034),
.B(n_531),
.C(n_530),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_5024),
.Y(n_5095)
);

NAND3xp33_ASAP7_75t_SL g5096 ( 
.A(n_5039),
.B(n_529),
.C(n_530),
.Y(n_5096)
);

O2A1O1Ixp5_ASAP7_75t_SL g5097 ( 
.A1(n_4999),
.A2(n_532),
.B(n_529),
.C(n_531),
.Y(n_5097)
);

NAND4xp75_ASAP7_75t_L g5098 ( 
.A(n_5037),
.B(n_535),
.C(n_533),
.D(n_534),
.Y(n_5098)
);

AOI221xp5_ASAP7_75t_L g5099 ( 
.A1(n_5044),
.A2(n_537),
.B1(n_533),
.B2(n_534),
.C(n_538),
.Y(n_5099)
);

A2O1A1Ixp33_ASAP7_75t_L g5100 ( 
.A1(n_5011),
.A2(n_540),
.B(n_537),
.C(n_539),
.Y(n_5100)
);

OAI21xp5_ASAP7_75t_SL g5101 ( 
.A1(n_5004),
.A2(n_540),
.B(n_541),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5050),
.Y(n_5102)
);

OAI21xp5_ASAP7_75t_L g5103 ( 
.A1(n_5028),
.A2(n_543),
.B(n_542),
.Y(n_5103)
);

AOI221xp5_ASAP7_75t_L g5104 ( 
.A1(n_5055),
.A2(n_545),
.B1(n_541),
.B2(n_544),
.C(n_546),
.Y(n_5104)
);

AOI221xp5_ASAP7_75t_L g5105 ( 
.A1(n_5006),
.A2(n_549),
.B1(n_544),
.B2(n_548),
.C(n_551),
.Y(n_5105)
);

AOI21xp33_ASAP7_75t_L g5106 ( 
.A1(n_4979),
.A2(n_548),
.B(n_549),
.Y(n_5106)
);

AOI21xp5_ASAP7_75t_L g5107 ( 
.A1(n_5026),
.A2(n_551),
.B(n_552),
.Y(n_5107)
);

AOI21xp5_ASAP7_75t_L g5108 ( 
.A1(n_5017),
.A2(n_553),
.B(n_554),
.Y(n_5108)
);

AOI221x1_ASAP7_75t_L g5109 ( 
.A1(n_5007),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.C(n_558),
.Y(n_5109)
);

NOR3xp33_ASAP7_75t_L g5110 ( 
.A(n_5016),
.B(n_5022),
.C(n_5018),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_SL g5111 ( 
.A(n_4996),
.B(n_556),
.Y(n_5111)
);

OAI21xp33_ASAP7_75t_L g5112 ( 
.A1(n_5020),
.A2(n_557),
.B(n_559),
.Y(n_5112)
);

O2A1O1Ixp33_ASAP7_75t_SL g5113 ( 
.A1(n_5013),
.A2(n_569),
.B(n_578),
.C(n_559),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_5027),
.A2(n_560),
.B(n_563),
.Y(n_5114)
);

OAI211xp5_ASAP7_75t_L g5115 ( 
.A1(n_5036),
.A2(n_564),
.B(n_560),
.C(n_563),
.Y(n_5115)
);

NAND4xp75_ASAP7_75t_L g5116 ( 
.A(n_5021),
.B(n_566),
.C(n_564),
.D(n_565),
.Y(n_5116)
);

OAI221xp5_ASAP7_75t_L g5117 ( 
.A1(n_5008),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.C(n_568),
.Y(n_5117)
);

NOR3xp33_ASAP7_75t_L g5118 ( 
.A(n_5012),
.B(n_571),
.C(n_570),
.Y(n_5118)
);

AOI221xp5_ASAP7_75t_L g5119 ( 
.A1(n_5014),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.C(n_572),
.Y(n_5119)
);

NAND2xp5_ASAP7_75t_L g5120 ( 
.A(n_5000),
.B(n_5023),
.Y(n_5120)
);

NOR3xp33_ASAP7_75t_SL g5121 ( 
.A(n_5029),
.B(n_573),
.C(n_574),
.Y(n_5121)
);

INVx1_ASAP7_75t_SL g5122 ( 
.A(n_5033),
.Y(n_5122)
);

NAND2xp5_ASAP7_75t_L g5123 ( 
.A(n_4985),
.B(n_573),
.Y(n_5123)
);

OAI211xp5_ASAP7_75t_SL g5124 ( 
.A1(n_5025),
.A2(n_576),
.B(n_574),
.C(n_575),
.Y(n_5124)
);

AOI211xp5_ASAP7_75t_L g5125 ( 
.A1(n_5001),
.A2(n_578),
.B(n_575),
.C(n_576),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_SL g5126 ( 
.A(n_5030),
.B(n_4992),
.Y(n_5126)
);

AOI22xp5_ASAP7_75t_L g5127 ( 
.A1(n_5019),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.Y(n_5127)
);

NOR3xp33_ASAP7_75t_L g5128 ( 
.A(n_4982),
.B(n_581),
.C(n_580),
.Y(n_5128)
);

A2O1A1Ixp33_ASAP7_75t_L g5129 ( 
.A1(n_5052),
.A2(n_583),
.B(n_579),
.C(n_582),
.Y(n_5129)
);

AOI221xp5_ASAP7_75t_L g5130 ( 
.A1(n_5046),
.A2(n_588),
.B1(n_582),
.B2(n_584),
.C(n_589),
.Y(n_5130)
);

AOI221xp5_ASAP7_75t_L g5131 ( 
.A1(n_5046),
.A2(n_590),
.B1(n_584),
.B2(n_589),
.C(n_591),
.Y(n_5131)
);

OAI21xp5_ASAP7_75t_SL g5132 ( 
.A1(n_4997),
.A2(n_593),
.B(n_594),
.Y(n_5132)
);

NAND4xp25_ASAP7_75t_L g5133 ( 
.A(n_5031),
.B(n_596),
.C(n_593),
.D(n_594),
.Y(n_5133)
);

AOI322xp5_ASAP7_75t_L g5134 ( 
.A1(n_4993),
.A2(n_602),
.A3(n_601),
.B1(n_598),
.B2(n_596),
.C1(n_597),
.C2(n_600),
.Y(n_5134)
);

O2A1O1Ixp5_ASAP7_75t_L g5135 ( 
.A1(n_4980),
.A2(n_602),
.B(n_598),
.C(n_600),
.Y(n_5135)
);

NOR3xp33_ASAP7_75t_L g5136 ( 
.A(n_4997),
.B(n_605),
.C(n_604),
.Y(n_5136)
);

AOI221xp5_ASAP7_75t_L g5137 ( 
.A1(n_5046),
.A2(n_608),
.B1(n_603),
.B2(n_607),
.C(n_609),
.Y(n_5137)
);

AO22x1_ASAP7_75t_L g5138 ( 
.A1(n_4974),
.A2(n_610),
.B1(n_607),
.B2(n_609),
.Y(n_5138)
);

AOI22xp5_ASAP7_75t_L g5139 ( 
.A1(n_4976),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_5041),
.B(n_611),
.Y(n_5140)
);

OAI211xp5_ASAP7_75t_L g5141 ( 
.A1(n_4980),
.A2(n_616),
.B(n_614),
.C(n_615),
.Y(n_5141)
);

NOR3xp33_ASAP7_75t_L g5142 ( 
.A(n_5056),
.B(n_614),
.C(n_615),
.Y(n_5142)
);

O2A1O1Ixp33_ASAP7_75t_L g5143 ( 
.A1(n_5058),
.A2(n_618),
.B(n_616),
.C(n_617),
.Y(n_5143)
);

AOI21xp33_ASAP7_75t_L g5144 ( 
.A1(n_5080),
.A2(n_617),
.B(n_618),
.Y(n_5144)
);

AOI21xp5_ASAP7_75t_L g5145 ( 
.A1(n_5063),
.A2(n_619),
.B(n_620),
.Y(n_5145)
);

OAI21xp33_ASAP7_75t_SL g5146 ( 
.A1(n_5089),
.A2(n_5133),
.B(n_5086),
.Y(n_5146)
);

OAI22xp5_ASAP7_75t_L g5147 ( 
.A1(n_5070),
.A2(n_622),
.B1(n_619),
.B2(n_621),
.Y(n_5147)
);

NOR2xp33_ASAP7_75t_L g5148 ( 
.A(n_5069),
.B(n_621),
.Y(n_5148)
);

OAI211xp5_ASAP7_75t_SL g5149 ( 
.A1(n_5126),
.A2(n_625),
.B(n_622),
.C(n_623),
.Y(n_5149)
);

A2O1A1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_5135),
.A2(n_627),
.B(n_625),
.C(n_626),
.Y(n_5150)
);

OAI22xp5_ASAP7_75t_L g5151 ( 
.A1(n_5066),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_5151)
);

O2A1O1Ixp33_ASAP7_75t_L g5152 ( 
.A1(n_5128),
.A2(n_631),
.B(n_628),
.C(n_629),
.Y(n_5152)
);

AND2x2_ASAP7_75t_L g5153 ( 
.A(n_5122),
.B(n_631),
.Y(n_5153)
);

AOI22xp33_ASAP7_75t_L g5154 ( 
.A1(n_5060),
.A2(n_5110),
.B1(n_5074),
.B2(n_5096),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_L g5155 ( 
.A(n_5138),
.B(n_632),
.Y(n_5155)
);

NAND3xp33_ASAP7_75t_SL g5156 ( 
.A(n_5077),
.B(n_633),
.C(n_634),
.Y(n_5156)
);

AOI21xp33_ASAP7_75t_SL g5157 ( 
.A1(n_5140),
.A2(n_633),
.B(n_635),
.Y(n_5157)
);

AOI221xp5_ASAP7_75t_L g5158 ( 
.A1(n_5119),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.C(n_640),
.Y(n_5158)
);

AOI22xp5_ASAP7_75t_L g5159 ( 
.A1(n_5136),
.A2(n_641),
.B1(n_638),
.B2(n_640),
.Y(n_5159)
);

AOI21xp5_ASAP7_75t_SL g5160 ( 
.A1(n_5109),
.A2(n_641),
.B(n_642),
.Y(n_5160)
);

NOR2xp33_ASAP7_75t_SL g5161 ( 
.A(n_5098),
.B(n_643),
.Y(n_5161)
);

NOR4xp25_ASAP7_75t_L g5162 ( 
.A(n_5141),
.B(n_644),
.C(n_642),
.D(n_643),
.Y(n_5162)
);

AOI221xp5_ASAP7_75t_L g5163 ( 
.A1(n_5078),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.C(n_647),
.Y(n_5163)
);

AOI221xp5_ASAP7_75t_L g5164 ( 
.A1(n_5057),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.C(n_649),
.Y(n_5164)
);

AOI221x1_ASAP7_75t_L g5165 ( 
.A1(n_5094),
.A2(n_650),
.B1(n_648),
.B2(n_649),
.C(n_651),
.Y(n_5165)
);

NOR2xp33_ASAP7_75t_L g5166 ( 
.A(n_5112),
.B(n_650),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_5134),
.B(n_651),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5071),
.Y(n_5168)
);

INVxp67_ASAP7_75t_L g5169 ( 
.A(n_5071),
.Y(n_5169)
);

XOR2xp5_ASAP7_75t_L g5170 ( 
.A(n_5116),
.B(n_652),
.Y(n_5170)
);

AND2x2_ASAP7_75t_L g5171 ( 
.A(n_5121),
.B(n_653),
.Y(n_5171)
);

OAI211xp5_ASAP7_75t_L g5172 ( 
.A1(n_5125),
.A2(n_655),
.B(n_653),
.C(n_654),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_5129),
.B(n_656),
.Y(n_5173)
);

AOI221xp5_ASAP7_75t_L g5174 ( 
.A1(n_5059),
.A2(n_659),
.B1(n_657),
.B2(n_658),
.C(n_661),
.Y(n_5174)
);

AOI21xp5_ASAP7_75t_L g5175 ( 
.A1(n_5113),
.A2(n_5107),
.B(n_5076),
.Y(n_5175)
);

NAND4xp25_ASAP7_75t_SL g5176 ( 
.A(n_5088),
.B(n_661),
.C(n_657),
.D(n_658),
.Y(n_5176)
);

OAI21xp33_ASAP7_75t_L g5177 ( 
.A1(n_5120),
.A2(n_662),
.B(n_664),
.Y(n_5177)
);

BUFx2_ASAP7_75t_L g5178 ( 
.A(n_5103),
.Y(n_5178)
);

AND2x2_ASAP7_75t_L g5179 ( 
.A(n_5073),
.B(n_5087),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_5061),
.B(n_662),
.Y(n_5180)
);

AOI221xp5_ASAP7_75t_SL g5181 ( 
.A1(n_5111),
.A2(n_667),
.B1(n_664),
.B2(n_666),
.C(n_668),
.Y(n_5181)
);

AOI21xp33_ASAP7_75t_L g5182 ( 
.A1(n_5064),
.A2(n_666),
.B(n_667),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5075),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_5118),
.B(n_668),
.Y(n_5184)
);

AOI221x1_ASAP7_75t_L g5185 ( 
.A1(n_5090),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.C(n_672),
.Y(n_5185)
);

OR2x2_ASAP7_75t_L g5186 ( 
.A(n_5083),
.B(n_669),
.Y(n_5186)
);

AOI221xp5_ASAP7_75t_L g5187 ( 
.A1(n_5132),
.A2(n_672),
.B1(n_670),
.B2(n_671),
.C(n_673),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_5062),
.B(n_5065),
.Y(n_5188)
);

AOI221x1_ASAP7_75t_L g5189 ( 
.A1(n_5108),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.C(n_676),
.Y(n_5189)
);

OAI211xp5_ASAP7_75t_SL g5190 ( 
.A1(n_5102),
.A2(n_677),
.B(n_675),
.C(n_676),
.Y(n_5190)
);

OAI21xp5_ASAP7_75t_L g5191 ( 
.A1(n_5114),
.A2(n_677),
.B(n_678),
.Y(n_5191)
);

NAND3xp33_ASAP7_75t_L g5192 ( 
.A(n_5097),
.B(n_678),
.C(n_679),
.Y(n_5192)
);

NOR2xp33_ASAP7_75t_L g5193 ( 
.A(n_5101),
.B(n_680),
.Y(n_5193)
);

OAI211xp5_ASAP7_75t_SL g5194 ( 
.A1(n_5095),
.A2(n_683),
.B(n_681),
.C(n_682),
.Y(n_5194)
);

AOI21xp5_ASAP7_75t_L g5195 ( 
.A1(n_5093),
.A2(n_681),
.B(n_682),
.Y(n_5195)
);

NAND4xp75_ASAP7_75t_L g5196 ( 
.A(n_5091),
.B(n_685),
.C(n_683),
.D(n_684),
.Y(n_5196)
);

OAI221xp5_ASAP7_75t_SL g5197 ( 
.A1(n_5081),
.A2(n_687),
.B1(n_684),
.B2(n_686),
.C(n_688),
.Y(n_5197)
);

AOI321xp33_ASAP7_75t_L g5198 ( 
.A1(n_5092),
.A2(n_689),
.A3(n_691),
.B1(n_687),
.B2(n_688),
.C(n_690),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_5082),
.B(n_689),
.Y(n_5199)
);

OAI211xp5_ASAP7_75t_L g5200 ( 
.A1(n_5115),
.A2(n_693),
.B(n_690),
.C(n_692),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_L g5201 ( 
.A(n_5117),
.B(n_692),
.Y(n_5201)
);

NOR3xp33_ASAP7_75t_L g5202 ( 
.A(n_5084),
.B(n_693),
.C(n_694),
.Y(n_5202)
);

OAI21xp33_ASAP7_75t_L g5203 ( 
.A1(n_5068),
.A2(n_5072),
.B(n_5100),
.Y(n_5203)
);

AOI22xp33_ASAP7_75t_SL g5204 ( 
.A1(n_5123),
.A2(n_5124),
.B1(n_5106),
.B2(n_5085),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_5139),
.B(n_694),
.Y(n_5205)
);

AOI221xp5_ASAP7_75t_L g5206 ( 
.A1(n_5079),
.A2(n_697),
.B1(n_695),
.B2(n_696),
.C(n_698),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_L g5207 ( 
.A(n_5127),
.B(n_695),
.Y(n_5207)
);

AO221x1_ASAP7_75t_L g5208 ( 
.A1(n_5130),
.A2(n_698),
.B1(n_696),
.B2(n_697),
.C(n_699),
.Y(n_5208)
);

NAND2xp5_ASAP7_75t_L g5209 ( 
.A(n_5067),
.B(n_700),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_5099),
.B(n_700),
.Y(n_5210)
);

NAND2xp5_ASAP7_75t_L g5211 ( 
.A(n_5104),
.B(n_701),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_5137),
.Y(n_5212)
);

NOR3xp33_ASAP7_75t_L g5213 ( 
.A(n_5131),
.B(n_5105),
.C(n_701),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_5089),
.Y(n_5214)
);

OAI21xp33_ASAP7_75t_L g5215 ( 
.A1(n_5080),
.A2(n_702),
.B(n_703),
.Y(n_5215)
);

AOI222xp33_ASAP7_75t_L g5216 ( 
.A1(n_5080),
.A2(n_705),
.B1(n_707),
.B2(n_703),
.C1(n_704),
.C2(n_706),
.Y(n_5216)
);

NOR2x1_ASAP7_75t_L g5217 ( 
.A(n_5089),
.B(n_704),
.Y(n_5217)
);

HB1xp67_ASAP7_75t_L g5218 ( 
.A(n_5089),
.Y(n_5218)
);

NAND4xp25_ASAP7_75t_SL g5219 ( 
.A(n_5152),
.B(n_710),
.C(n_707),
.D(n_708),
.Y(n_5219)
);

NAND3xp33_ASAP7_75t_L g5220 ( 
.A(n_5142),
.B(n_5161),
.C(n_5165),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_SL g5221 ( 
.A(n_5162),
.B(n_708),
.Y(n_5221)
);

INVx2_ASAP7_75t_SL g5222 ( 
.A(n_5217),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_5153),
.B(n_710),
.Y(n_5223)
);

AOI211xp5_ASAP7_75t_L g5224 ( 
.A1(n_5144),
.A2(n_715),
.B(n_711),
.C(n_712),
.Y(n_5224)
);

INVx1_ASAP7_75t_L g5225 ( 
.A(n_5218),
.Y(n_5225)
);

OAI32xp33_ASAP7_75t_L g5226 ( 
.A1(n_5146),
.A2(n_719),
.A3(n_716),
.B1(n_718),
.B2(n_720),
.Y(n_5226)
);

AOI221xp5_ASAP7_75t_L g5227 ( 
.A1(n_5143),
.A2(n_721),
.B1(n_718),
.B2(n_719),
.C(n_722),
.Y(n_5227)
);

AOI211xp5_ASAP7_75t_SL g5228 ( 
.A1(n_5160),
.A2(n_724),
.B(n_721),
.C(n_723),
.Y(n_5228)
);

O2A1O1Ixp33_ASAP7_75t_L g5229 ( 
.A1(n_5169),
.A2(n_725),
.B(n_723),
.C(n_724),
.Y(n_5229)
);

NOR2x1_ASAP7_75t_L g5230 ( 
.A(n_5168),
.B(n_725),
.Y(n_5230)
);

AOI221xp5_ASAP7_75t_L g5231 ( 
.A1(n_5214),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.C(n_729),
.Y(n_5231)
);

AOI21xp5_ASAP7_75t_L g5232 ( 
.A1(n_5175),
.A2(n_726),
.B(n_729),
.Y(n_5232)
);

NAND3xp33_ASAP7_75t_L g5233 ( 
.A(n_5216),
.B(n_730),
.C(n_731),
.Y(n_5233)
);

OAI21xp33_ASAP7_75t_SL g5234 ( 
.A1(n_5154),
.A2(n_5188),
.B(n_5155),
.Y(n_5234)
);

OAI221xp5_ASAP7_75t_SL g5235 ( 
.A1(n_5203),
.A2(n_732),
.B1(n_730),
.B2(n_731),
.C(n_733),
.Y(n_5235)
);

AOI322xp5_ASAP7_75t_L g5236 ( 
.A1(n_5156),
.A2(n_738),
.A3(n_737),
.B1(n_735),
.B2(n_733),
.C1(n_734),
.C2(n_736),
.Y(n_5236)
);

OAI211xp5_ASAP7_75t_L g5237 ( 
.A1(n_5200),
.A2(n_5158),
.B(n_5215),
.C(n_5172),
.Y(n_5237)
);

OAI221xp5_ASAP7_75t_SL g5238 ( 
.A1(n_5213),
.A2(n_736),
.B1(n_734),
.B2(n_735),
.C(n_737),
.Y(n_5238)
);

OAI221xp5_ASAP7_75t_SL g5239 ( 
.A1(n_5212),
.A2(n_5186),
.B1(n_5204),
.B2(n_5150),
.C(n_5178),
.Y(n_5239)
);

OAI211xp5_ASAP7_75t_L g5240 ( 
.A1(n_5174),
.A2(n_740),
.B(n_738),
.C(n_739),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_L g5241 ( 
.A(n_5171),
.B(n_739),
.Y(n_5241)
);

AOI211xp5_ASAP7_75t_SL g5242 ( 
.A1(n_5167),
.A2(n_743),
.B(n_741),
.C(n_742),
.Y(n_5242)
);

INVx1_ASAP7_75t_SL g5243 ( 
.A(n_5170),
.Y(n_5243)
);

AOI321xp33_ASAP7_75t_L g5244 ( 
.A1(n_5179),
.A2(n_746),
.A3(n_748),
.B1(n_741),
.B2(n_745),
.C(n_747),
.Y(n_5244)
);

OAI22xp5_ASAP7_75t_L g5245 ( 
.A1(n_5159),
.A2(n_749),
.B1(n_747),
.B2(n_748),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_5145),
.A2(n_749),
.B(n_750),
.Y(n_5246)
);

AOI221xp5_ASAP7_75t_L g5247 ( 
.A1(n_5192),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.C(n_753),
.Y(n_5247)
);

NOR2xp33_ASAP7_75t_SL g5248 ( 
.A(n_5197),
.B(n_752),
.Y(n_5248)
);

AOI211xp5_ASAP7_75t_L g5249 ( 
.A1(n_5176),
.A2(n_756),
.B(n_754),
.C(n_755),
.Y(n_5249)
);

AOI221xp5_ASAP7_75t_L g5250 ( 
.A1(n_5157),
.A2(n_758),
.B1(n_755),
.B2(n_756),
.C(n_759),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_5208),
.B(n_758),
.Y(n_5251)
);

AOI22xp33_ASAP7_75t_L g5252 ( 
.A1(n_5183),
.A2(n_761),
.B1(n_759),
.B2(n_760),
.Y(n_5252)
);

AOI21xp33_ASAP7_75t_SL g5253 ( 
.A1(n_5147),
.A2(n_764),
.B(n_762),
.Y(n_5253)
);

AOI22xp5_ASAP7_75t_L g5254 ( 
.A1(n_5148),
.A2(n_5166),
.B1(n_5193),
.B2(n_5201),
.Y(n_5254)
);

NAND3xp33_ASAP7_75t_L g5255 ( 
.A(n_5185),
.B(n_5189),
.C(n_5206),
.Y(n_5255)
);

NOR2xp33_ASAP7_75t_L g5256 ( 
.A(n_5177),
.B(n_760),
.Y(n_5256)
);

NAND2xp5_ASAP7_75t_L g5257 ( 
.A(n_5187),
.B(n_762),
.Y(n_5257)
);

OA22x2_ASAP7_75t_L g5258 ( 
.A1(n_5191),
.A2(n_767),
.B1(n_765),
.B2(n_766),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_5181),
.B(n_766),
.Y(n_5259)
);

AOI221xp5_ASAP7_75t_L g5260 ( 
.A1(n_5195),
.A2(n_769),
.B1(n_767),
.B2(n_768),
.C(n_770),
.Y(n_5260)
);

AOI21xp33_ASAP7_75t_L g5261 ( 
.A1(n_5211),
.A2(n_768),
.B(n_770),
.Y(n_5261)
);

AOI221xp5_ASAP7_75t_L g5262 ( 
.A1(n_5202),
.A2(n_774),
.B1(n_771),
.B2(n_772),
.C(n_775),
.Y(n_5262)
);

O2A1O1Ixp33_ASAP7_75t_L g5263 ( 
.A1(n_5173),
.A2(n_777),
.B(n_772),
.C(n_776),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5184),
.Y(n_5264)
);

NAND4xp25_ASAP7_75t_SL g5265 ( 
.A(n_5164),
.B(n_779),
.C(n_776),
.D(n_778),
.Y(n_5265)
);

AOI22xp5_ASAP7_75t_L g5266 ( 
.A1(n_5149),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_5266)
);

AOI221xp5_ASAP7_75t_L g5267 ( 
.A1(n_5151),
.A2(n_5210),
.B1(n_5199),
.B2(n_5209),
.C(n_5194),
.Y(n_5267)
);

OAI21xp5_ASAP7_75t_L g5268 ( 
.A1(n_5180),
.A2(n_780),
.B(n_781),
.Y(n_5268)
);

AO21x1_ASAP7_75t_L g5269 ( 
.A1(n_5205),
.A2(n_782),
.B(n_783),
.Y(n_5269)
);

AOI21xp33_ASAP7_75t_L g5270 ( 
.A1(n_5207),
.A2(n_782),
.B(n_783),
.Y(n_5270)
);

AND2x2_ASAP7_75t_L g5271 ( 
.A(n_5196),
.B(n_785),
.Y(n_5271)
);

XNOR2x2_ASAP7_75t_L g5272 ( 
.A(n_5163),
.B(n_785),
.Y(n_5272)
);

NAND2xp33_ASAP7_75t_SL g5273 ( 
.A(n_5198),
.B(n_786),
.Y(n_5273)
);

NOR3xp33_ASAP7_75t_L g5274 ( 
.A(n_5182),
.B(n_794),
.C(n_786),
.Y(n_5274)
);

NOR2x1_ASAP7_75t_L g5275 ( 
.A(n_5230),
.B(n_5190),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_5228),
.B(n_788),
.Y(n_5276)
);

OAI22xp5_ASAP7_75t_L g5277 ( 
.A1(n_5266),
.A2(n_789),
.B1(n_787),
.B2(n_788),
.Y(n_5277)
);

NOR2xp33_ASAP7_75t_L g5278 ( 
.A(n_5251),
.B(n_787),
.Y(n_5278)
);

OAI22x1_ASAP7_75t_L g5279 ( 
.A1(n_5219),
.A2(n_792),
.B1(n_790),
.B2(n_791),
.Y(n_5279)
);

NAND4xp75_ASAP7_75t_L g5280 ( 
.A(n_5234),
.B(n_794),
.C(n_790),
.D(n_793),
.Y(n_5280)
);

NAND3xp33_ASAP7_75t_L g5281 ( 
.A(n_5247),
.B(n_793),
.C(n_795),
.Y(n_5281)
);

NAND2xp5_ASAP7_75t_L g5282 ( 
.A(n_5223),
.B(n_796),
.Y(n_5282)
);

NOR4xp75_ASAP7_75t_L g5283 ( 
.A(n_5221),
.B(n_798),
.C(n_795),
.D(n_797),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_5258),
.Y(n_5284)
);

NAND3xp33_ASAP7_75t_SL g5285 ( 
.A(n_5269),
.B(n_797),
.C(n_798),
.Y(n_5285)
);

NOR2xp33_ASAP7_75t_L g5286 ( 
.A(n_5222),
.B(n_5240),
.Y(n_5286)
);

NAND3xp33_ASAP7_75t_L g5287 ( 
.A(n_5242),
.B(n_799),
.C(n_800),
.Y(n_5287)
);

NOR2xp33_ASAP7_75t_L g5288 ( 
.A(n_5238),
.B(n_799),
.Y(n_5288)
);

OAI322xp33_ASAP7_75t_L g5289 ( 
.A1(n_5248),
.A2(n_828),
.A3(n_811),
.B1(n_837),
.B2(n_840),
.C1(n_820),
.C2(n_800),
.Y(n_5289)
);

INVxp67_ASAP7_75t_SL g5290 ( 
.A(n_5229),
.Y(n_5290)
);

NOR3xp33_ASAP7_75t_L g5291 ( 
.A(n_5239),
.B(n_802),
.C(n_803),
.Y(n_5291)
);

NOR3xp33_ASAP7_75t_L g5292 ( 
.A(n_5225),
.B(n_802),
.C(n_803),
.Y(n_5292)
);

NOR2xp67_ASAP7_75t_L g5293 ( 
.A(n_5220),
.B(n_5255),
.Y(n_5293)
);

AO22x2_ASAP7_75t_L g5294 ( 
.A1(n_5243),
.A2(n_807),
.B1(n_804),
.B2(n_806),
.Y(n_5294)
);

NOR2x1_ASAP7_75t_L g5295 ( 
.A(n_5241),
.B(n_808),
.Y(n_5295)
);

NOR2xp33_ASAP7_75t_L g5296 ( 
.A(n_5265),
.B(n_808),
.Y(n_5296)
);

NOR2x1_ASAP7_75t_L g5297 ( 
.A(n_5232),
.B(n_809),
.Y(n_5297)
);

NOR4xp25_ASAP7_75t_L g5298 ( 
.A(n_5237),
.B(n_814),
.C(n_812),
.D(n_813),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_5271),
.Y(n_5299)
);

OAI222xp33_ASAP7_75t_L g5300 ( 
.A1(n_5254),
.A2(n_814),
.B1(n_816),
.B2(n_812),
.C1(n_813),
.C2(n_815),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_5259),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_5236),
.B(n_815),
.Y(n_5302)
);

NOR2x1_ASAP7_75t_L g5303 ( 
.A(n_5233),
.B(n_816),
.Y(n_5303)
);

NOR4xp75_ASAP7_75t_L g5304 ( 
.A(n_5268),
.B(n_820),
.C(n_817),
.D(n_819),
.Y(n_5304)
);

NOR2x1_ASAP7_75t_L g5305 ( 
.A(n_5263),
.B(n_817),
.Y(n_5305)
);

NOR3xp33_ASAP7_75t_L g5306 ( 
.A(n_5261),
.B(n_819),
.C(n_821),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5272),
.Y(n_5307)
);

NAND4xp75_ASAP7_75t_L g5308 ( 
.A(n_5227),
.B(n_823),
.C(n_821),
.D(n_822),
.Y(n_5308)
);

INVx1_ASAP7_75t_SL g5309 ( 
.A(n_5273),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5294),
.Y(n_5310)
);

AND2x4_ASAP7_75t_L g5311 ( 
.A(n_5295),
.B(n_5274),
.Y(n_5311)
);

NOR2xp67_ASAP7_75t_SL g5312 ( 
.A(n_5280),
.B(n_5264),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_5294),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5276),
.Y(n_5314)
);

NAND2x1_ASAP7_75t_L g5315 ( 
.A(n_5275),
.B(n_5246),
.Y(n_5315)
);

NAND4xp75_ASAP7_75t_L g5316 ( 
.A(n_5293),
.B(n_5257),
.C(n_5267),
.D(n_5270),
.Y(n_5316)
);

NAND4xp75_ASAP7_75t_L g5317 ( 
.A(n_5303),
.B(n_5256),
.C(n_5262),
.D(n_5260),
.Y(n_5317)
);

NOR2xp33_ASAP7_75t_L g5318 ( 
.A(n_5289),
.B(n_5287),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5282),
.Y(n_5319)
);

NOR2x1_ASAP7_75t_L g5320 ( 
.A(n_5285),
.B(n_5307),
.Y(n_5320)
);

NAND3xp33_ASAP7_75t_L g5321 ( 
.A(n_5291),
.B(n_5224),
.C(n_5249),
.Y(n_5321)
);

NOR2x1_ASAP7_75t_L g5322 ( 
.A(n_5300),
.B(n_5245),
.Y(n_5322)
);

NOR3xp33_ASAP7_75t_L g5323 ( 
.A(n_5278),
.B(n_5253),
.C(n_5250),
.Y(n_5323)
);

INVx1_ASAP7_75t_SL g5324 ( 
.A(n_5283),
.Y(n_5324)
);

NAND4xp25_ASAP7_75t_L g5325 ( 
.A(n_5286),
.B(n_5244),
.C(n_5235),
.D(n_5231),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_5279),
.Y(n_5326)
);

AND4x2_ASAP7_75t_L g5327 ( 
.A(n_5297),
.B(n_5226),
.C(n_5252),
.D(n_824),
.Y(n_5327)
);

NOR2xp67_ASAP7_75t_SL g5328 ( 
.A(n_5316),
.B(n_5299),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_5310),
.B(n_5298),
.Y(n_5329)
);

NOR4xp75_ASAP7_75t_SL g5330 ( 
.A(n_5327),
.B(n_5302),
.C(n_5277),
.D(n_5309),
.Y(n_5330)
);

OR2x2_ASAP7_75t_L g5331 ( 
.A(n_5325),
.B(n_5284),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_5313),
.Y(n_5332)
);

AOI221xp5_ASAP7_75t_L g5333 ( 
.A1(n_5312),
.A2(n_5290),
.B1(n_5288),
.B2(n_5281),
.C(n_5296),
.Y(n_5333)
);

NAND4xp75_ASAP7_75t_L g5334 ( 
.A(n_5320),
.B(n_5305),
.C(n_5301),
.D(n_5306),
.Y(n_5334)
);

NOR2xp33_ASAP7_75t_L g5335 ( 
.A(n_5324),
.B(n_5308),
.Y(n_5335)
);

AOI211xp5_ASAP7_75t_L g5336 ( 
.A1(n_5321),
.A2(n_5292),
.B(n_5304),
.C(n_825),
.Y(n_5336)
);

INVx1_ASAP7_75t_L g5337 ( 
.A(n_5326),
.Y(n_5337)
);

INVx3_ASAP7_75t_SL g5338 ( 
.A(n_5311),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_5336),
.B(n_5311),
.Y(n_5339)
);

NAND2xp33_ASAP7_75t_R g5340 ( 
.A(n_5329),
.B(n_5314),
.Y(n_5340)
);

NOR2xp33_ASAP7_75t_R g5341 ( 
.A(n_5338),
.B(n_5319),
.Y(n_5341)
);

NOR2xp33_ASAP7_75t_R g5342 ( 
.A(n_5337),
.B(n_5318),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_SL g5343 ( 
.A(n_5330),
.B(n_5322),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_5332),
.B(n_5323),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_5328),
.B(n_5315),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5345),
.Y(n_5346)
);

OAI22xp5_ASAP7_75t_SL g5347 ( 
.A1(n_5344),
.A2(n_5335),
.B1(n_5331),
.B2(n_5334),
.Y(n_5347)
);

INVx3_ASAP7_75t_L g5348 ( 
.A(n_5339),
.Y(n_5348)
);

OAI22xp5_ASAP7_75t_SL g5349 ( 
.A1(n_5340),
.A2(n_5333),
.B1(n_5317),
.B2(n_825),
.Y(n_5349)
);

INVx1_ASAP7_75t_SL g5350 ( 
.A(n_5341),
.Y(n_5350)
);

OR3x2_ASAP7_75t_L g5351 ( 
.A(n_5346),
.B(n_5342),
.C(n_5343),
.Y(n_5351)
);

NOR2xp33_ASAP7_75t_L g5352 ( 
.A(n_5350),
.B(n_822),
.Y(n_5352)
);

INVxp67_ASAP7_75t_L g5353 ( 
.A(n_5352),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5353),
.Y(n_5354)
);

OAI22x1_ASAP7_75t_L g5355 ( 
.A1(n_5354),
.A2(n_5348),
.B1(n_5351),
.B2(n_5349),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_5355),
.A2(n_5347),
.B(n_823),
.Y(n_5356)
);

OAI21xp5_ASAP7_75t_L g5357 ( 
.A1(n_5356),
.A2(n_826),
.B(n_827),
.Y(n_5357)
);

AOI21xp33_ASAP7_75t_SL g5358 ( 
.A1(n_5357),
.A2(n_826),
.B(n_828),
.Y(n_5358)
);

OAI21x1_ASAP7_75t_L g5359 ( 
.A1(n_5358),
.A2(n_829),
.B(n_830),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_5359),
.Y(n_5360)
);

AOI221xp5_ASAP7_75t_L g5361 ( 
.A1(n_5360),
.A2(n_833),
.B1(n_829),
.B2(n_831),
.C(n_834),
.Y(n_5361)
);

AOI21xp5_ASAP7_75t_L g5362 ( 
.A1(n_5361),
.A2(n_831),
.B(n_833),
.Y(n_5362)
);

AOI211xp5_ASAP7_75t_L g5363 ( 
.A1(n_5362),
.A2(n_836),
.B(n_834),
.C(n_835),
.Y(n_5363)
);


endmodule