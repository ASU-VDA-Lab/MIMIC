module fake_jpeg_23119_n_325 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_37),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_20),
.C(n_24),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_27),
.B1(n_28),
.B2(n_16),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_53),
.B1(n_58),
.B2(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_27),
.B1(n_16),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_57),
.B1(n_38),
.B2(n_14),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_27),
.B1(n_16),
.B2(n_26),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_61),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_66),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_20),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_81),
.B1(n_55),
.B2(n_56),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_16),
.B1(n_26),
.B2(n_20),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_74),
.B(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_77),
.Y(n_94)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_38),
.B1(n_24),
.B2(n_30),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_83),
.B(n_88),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_57),
.B(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_89),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_24),
.B1(n_53),
.B2(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_30),
.B1(n_24),
.B2(n_46),
.Y(n_86)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_58),
.B(n_41),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_26),
.B1(n_14),
.B2(n_49),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_103),
.Y(n_125)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_102),
.Y(n_109)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_32),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_101),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_69),
.C(n_75),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_61),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_32),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_101),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_126),
.B1(n_130),
.B2(n_92),
.Y(n_143)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_104),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_39),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_82),
.B1(n_85),
.B2(n_95),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_144),
.B1(n_151),
.B2(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_103),
.B1(n_84),
.B2(n_88),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_148),
.B1(n_154),
.B2(n_147),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_90),
.B(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_118),
.B1(n_120),
.B2(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_90),
.B1(n_80),
.B2(n_78),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_87),
.B1(n_76),
.B2(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_34),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_18),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_59),
.B1(n_65),
.B2(n_33),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_59),
.B1(n_33),
.B2(n_37),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_154),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_174),
.B(n_181),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_162),
.Y(n_195)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_130),
.B1(n_117),
.B2(n_126),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_176),
.B1(n_178),
.B2(n_145),
.Y(n_200)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_173),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_125),
.C(n_110),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_144),
.C(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_115),
.B1(n_104),
.B2(n_14),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_37),
.B1(n_17),
.B2(n_19),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_177),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_104),
.B1(n_25),
.B2(n_17),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_143),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_133),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_196),
.B1(n_203),
.B2(n_204),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_151),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_135),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_205),
.C(n_207),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_166),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_201),
.B1(n_208),
.B2(n_205),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_148),
.B1(n_141),
.B2(n_137),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_132),
.C(n_139),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_137),
.C(n_136),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_148),
.B1(n_136),
.B2(n_153),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_157),
.B(n_182),
.CI(n_164),
.CON(n_209),
.SN(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_219),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_173),
.B1(n_171),
.B2(n_167),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_220),
.B1(n_19),
.B2(n_21),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_184),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_215),
.B(n_225),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_226),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_157),
.B1(n_165),
.B2(n_181),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_228),
.B1(n_17),
.B2(n_19),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_165),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_97),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_93),
.C(n_127),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_187),
.C(n_188),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_64),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_18),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_0),
.B(n_1),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_194),
.B(n_25),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_238),
.C(n_240),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_208),
.B1(n_199),
.B2(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_236),
.B1(n_243),
.B2(n_247),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_198),
.B1(n_207),
.B2(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_186),
.C(n_107),
.Y(n_238)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_63),
.C(n_62),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_230),
.B(n_18),
.C(n_216),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_63),
.C(n_62),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_232),
.C(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_60),
.B1(n_22),
.B2(n_21),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_231),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_60),
.B1(n_22),
.B2(n_33),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_18),
.B1(n_33),
.B2(n_35),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_256),
.C(n_259),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_261),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_231),
.C(n_226),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_229),
.B(n_9),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_260),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_13),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_13),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_12),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_11),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_268),
.B(n_237),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_235),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_275),
.C(n_279),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_233),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_270),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_254),
.C(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_247),
.B1(n_249),
.B2(n_248),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_283),
.B1(n_0),
.B2(n_1),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_252),
.B(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_258),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

NAND2xp67_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_261),
.B(n_8),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_290),
.A2(n_3),
.B(n_4),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_296),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_279),
.C(n_274),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_305),
.C(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_272),
.C(n_35),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_302),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_291),
.B1(n_287),
.B2(n_286),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_312),
.B(n_300),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_4),
.B(n_5),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_303),
.B(n_298),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_305),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_313),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_315),
.C(n_6),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_6),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_7),
.B(n_285),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_7),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_7),
.Y(n_325)
);


endmodule