module fake_jpeg_14853_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx14_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_24),
.Y(n_26)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_18),
.B1(n_14),
.B2(n_9),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_9),
.B1(n_23),
.B2(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_19),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_12),
.B(n_18),
.C(n_14),
.Y(n_31)
);

OAI32xp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_24),
.A3(n_11),
.B1(n_15),
.B2(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_29),
.B1(n_19),
.B2(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_11),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_37),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_20),
.B1(n_15),
.B2(n_19),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_36),
.B1(n_33),
.B2(n_39),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_20),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_3),
.B(n_4),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_34),
.Y(n_56)
);

OA21x2_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_4),
.B(n_6),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_36),
.B(n_32),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_28),
.C(n_6),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_45),
.C(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_49),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_60),
.B1(n_51),
.B2(n_54),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_44),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_58),
.C(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_69),
.Y(n_73)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_65),
.B(n_62),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_65),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_4),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_68),
.B(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_7),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_8),
.B(n_61),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_76),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_78),
.Y(n_81)
);


endmodule