module real_jpeg_10333_n_16 (n_5, n_4, n_8, n_0, n_12, n_318, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_318;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_1),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_141),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_141),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_141),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_2),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_159),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_159),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_159),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_32),
.B1(n_48),
.B2(n_50),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_32),
.B1(n_64),
.B2(n_65),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_10),
.A2(n_35),
.B1(n_48),
.B2(n_50),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_35),
.B1(n_64),
.B2(n_65),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_11),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_168),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_168),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_168),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_13),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_53),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_13),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_15),
.A2(n_50),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_15),
.B(n_50),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_15),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_15),
.A2(n_88),
.B1(n_91),
.B2(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_15),
.B(n_103),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_15),
.A2(n_25),
.B(n_27),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_177),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_104),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_84),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_21),
.A2(n_72),
.B1(n_73),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_21),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_22),
.A2(n_23),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_23),
.B(n_58),
.C(n_71),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_33),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_28),
.B(n_31),
.C(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_24),
.A2(n_29),
.B1(n_37),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_24),
.A2(n_37),
.B1(n_260),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_24),
.A2(n_37),
.B1(n_140),
.B2(n_269),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_44),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g202 ( 
.A(n_27),
.B(n_177),
.CON(n_202),
.SN(n_202)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_28),
.A2(n_31),
.B(n_177),
.C(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_34),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_36),
.A2(n_103),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_37),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_37),
.A2(n_140),
.B(n_142),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_58),
.B1(n_59),
.B2(n_71),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_51),
.B(n_54),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_42),
.A2(n_57),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_42),
.A2(n_57),
.B1(n_220),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_42),
.A2(n_113),
.B(n_256),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_47),
.B1(n_52),
.B2(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_43),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_43),
.A2(n_47),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_43),
.A2(n_55),
.B(n_114),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_44),
.B(n_50),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_46),
.A2(n_48),
.B1(n_202),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_56),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_57),
.A2(n_76),
.B(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_57),
.B(n_177),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_59),
.B1(n_112),
.B2(n_117),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_68),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_63),
.B1(n_95),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_60),
.A2(n_63),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_60),
.A2(n_63),
.B1(n_167),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_60),
.A2(n_63),
.B1(n_192),
.B2(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_60),
.A2(n_78),
.B(n_200),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_63),
.B(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_63),
.A2(n_80),
.B(n_137),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_64),
.B(n_67),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_64),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_65),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_169)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_69),
.A2(n_83),
.B(n_97),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_98),
.B(n_99),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_86),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_98),
.B1(n_99),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_87),
.A2(n_94),
.B1(n_98),
.B2(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_88),
.A2(n_91),
.B1(n_158),
.B2(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_88),
.A2(n_135),
.B(n_161),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_88),
.A2(n_92),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_88),
.A2(n_91),
.B1(n_224),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_88),
.A2(n_210),
.B(n_246),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_89),
.B(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_89),
.A2(n_90),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_90),
.B(n_134),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_91),
.B(n_177),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_91),
.A2(n_133),
.B(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_94),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_101),
.B(n_103),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_119),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_118),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_148),
.B(n_316),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_145),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_123),
.B(n_145),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_124),
.B(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_124),
.B(n_308),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_129),
.CI(n_130),
.CON(n_124),
.SN(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.C(n_143),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_131),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_132),
.B(n_136),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

AOI321xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_295),
.A3(n_307),
.B1(n_309),
.B2(n_315),
.C(n_318),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_262),
.C(n_291),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_236),
.B(n_261),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_213),
.B(n_235),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_195),
.B(n_212),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_186),
.B(n_194),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_174),
.B(n_185),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_162),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_169),
.B2(n_173),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_180),
.B(n_184),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_196),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.CI(n_193),
.CON(n_189),
.SN(n_189)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_206),
.B2(n_211),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_199),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_205),
.C(n_211),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_203),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_215),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_229),
.B2(n_230),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_232),
.C(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_228),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.C(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_231),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_238),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_250),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_249),
.C(n_250),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_245),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_254),
.C(n_257),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_278),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_278),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_272),
.C(n_276),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_267),
.C(n_271),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_270),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_273),
.B1(n_276),
.B2(n_277),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_278)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_287),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_287),
.C(n_288),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_283),
.C(n_286),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_293),
.Y(n_312)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_298),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_306),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_304),
.C(n_306),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_310)
);


endmodule