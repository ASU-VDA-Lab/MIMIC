module fake_jpeg_22103_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_23),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_1),
.C(n_3),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_4),
.C(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_5),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_4),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_6),
.C(n_8),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_14),
.B1(n_17),
.B2(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_15),
.B1(n_24),
.B2(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_13),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_42),
.B1(n_47),
.B2(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_17),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_30),
.C(n_36),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_15),
.B(n_6),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_35),
.C(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_59),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_48),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.C(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_46),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_39),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_63),
.B(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_61),
.C(n_58),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_66),
.B(n_65),
.Y(n_71)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_49),
.B1(n_55),
.B2(n_31),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_31),
.B1(n_42),
.B2(n_33),
.Y(n_73)
);


endmodule