module fake_jpeg_8439_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx13_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_3),
.B(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_23),
.B1(n_24),
.B2(n_14),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp33_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_4),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_15),
.B1(n_20),
.B2(n_24),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_10),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_34),
.B1(n_26),
.B2(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_28),
.B1(n_15),
.B2(n_29),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.C(n_38),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_31),
.C(n_27),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_23),
.B1(n_20),
.B2(n_24),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_40),
.B(n_7),
.C(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_43),
.Y(n_44)
);


endmodule