module real_aes_8857_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g507 ( .A(n_1), .Y(n_507) );
INVx1_ASAP7_75t_L g264 ( .A(n_2), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_3), .A2(n_39), .B1(n_183), .B2(n_535), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g171 ( .A1(n_4), .A2(n_172), .B(n_173), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_5), .B(n_170), .Y(n_484) );
AND2x6_ASAP7_75t_L g145 ( .A(n_6), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_8), .B(n_40), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_8), .B(n_40), .Y(n_448) );
INVx1_ASAP7_75t_L g180 ( .A(n_9), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_10), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g142 ( .A(n_11), .Y(n_142) );
INVx1_ASAP7_75t_L g503 ( .A(n_12), .Y(n_503) );
INVx1_ASAP7_75t_L g246 ( .A(n_13), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_14), .B(n_148), .Y(n_541) );
AOI222xp33_ASAP7_75t_SL g452 ( .A1(n_15), .A2(n_453), .B1(n_454), .B2(n_463), .C1(n_751), .C2(n_752), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_16), .B(n_138), .Y(n_512) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_17), .B(n_121), .Y(n_120) );
AO32x2_ASAP7_75t_L g532 ( .A1(n_17), .A2(n_137), .A3(n_170), .B1(n_495), .B2(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_18), .B(n_183), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_19), .B(n_191), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_20), .B(n_138), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_21), .A2(n_51), .B1(n_183), .B2(n_535), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_22), .B(n_172), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_23), .A2(n_78), .B1(n_148), .B2(n_183), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_24), .B(n_183), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_25), .B(n_168), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_26), .A2(n_455), .B1(n_456), .B2(n_462), .Y(n_454) );
INVx1_ASAP7_75t_L g462 ( .A(n_26), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_27), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_28), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_29), .B(n_185), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_30), .B(n_178), .Y(n_265) );
INVx1_ASAP7_75t_L g156 ( .A(n_31), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_32), .A2(n_105), .B1(n_113), .B2(n_756), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_33), .B(n_185), .Y(n_529) );
INVx2_ASAP7_75t_L g150 ( .A(n_34), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_35), .B(n_183), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_36), .B(n_185), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_37), .A2(n_43), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_37), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_38), .A2(n_145), .B(n_157), .C(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g154 ( .A(n_41), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_42), .B(n_178), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_43), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_44), .B(n_183), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_45), .A2(n_88), .B1(n_208), .B2(n_535), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_46), .B(n_183), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_47), .B(n_183), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g160 ( .A(n_48), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_49), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_50), .B(n_172), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_52), .A2(n_61), .B1(n_148), .B2(n_183), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_53), .A2(n_148), .B1(n_151), .B2(n_157), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_54), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_55), .B(n_183), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_56), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_57), .B(n_183), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_58), .A2(n_177), .B(n_179), .C(n_182), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_59), .Y(n_221) );
INVx1_ASAP7_75t_L g174 ( .A(n_60), .Y(n_174) );
INVx1_ASAP7_75t_L g146 ( .A(n_62), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_63), .B(n_183), .Y(n_508) );
INVx1_ASAP7_75t_L g141 ( .A(n_64), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
AO32x2_ASAP7_75t_L g552 ( .A1(n_66), .A2(n_170), .A3(n_226), .B1(n_495), .B2(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g492 ( .A(n_67), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_68), .A2(n_124), .B1(n_125), .B2(n_128), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_68), .Y(n_128) );
INVx1_ASAP7_75t_L g524 ( .A(n_69), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_SL g190 ( .A1(n_70), .A2(n_182), .B(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g193 ( .A(n_71), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_72), .B(n_148), .Y(n_525) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_74), .Y(n_165) );
INVx1_ASAP7_75t_L g214 ( .A(n_75), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_76), .A2(n_102), .B1(n_460), .B2(n_461), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_76), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_77), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_79), .A2(n_145), .B(n_157), .C(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_80), .B(n_535), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_81), .B(n_148), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_82), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_84), .B(n_191), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_85), .B(n_148), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_86), .A2(n_145), .B(n_157), .C(n_263), .Y(n_262) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_87), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g445 ( .A(n_87), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g466 ( .A(n_87), .B(n_447), .Y(n_466) );
INVx2_ASAP7_75t_L g750 ( .A(n_87), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_89), .A2(n_103), .B1(n_148), .B2(n_149), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_90), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_91), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_92), .A2(n_145), .B(n_157), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_93), .Y(n_236) );
INVx1_ASAP7_75t_L g189 ( .A(n_94), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_95), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_96), .B(n_204), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_97), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_97), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_98), .B(n_148), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_99), .B(n_170), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_101), .A2(n_172), .B(n_188), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_102), .Y(n_461) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g756 ( .A(n_106), .Y(n_756) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g447 ( .A(n_109), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_451), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g755 ( .A(n_118), .Y(n_755) );
OAI21x1_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_442), .B(n_449), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_129), .B2(n_130), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_129), .A2(n_464), .B1(n_467), .B2(n_747), .Y(n_463) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_130), .A2(n_464), .B1(n_753), .B2(n_754), .Y(n_752) );
AND3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_367), .C(n_416), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_274), .C(n_312), .Y(n_131) );
OAI222xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_195), .B1(n_249), .B2(n_255), .C1(n_269), .C2(n_272), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_166), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_134), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_134), .B(n_317), .Y(n_408) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g285 ( .A(n_135), .B(n_186), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_135), .B(n_167), .Y(n_293) );
AND2x2_ASAP7_75t_L g328 ( .A(n_135), .B(n_305), .Y(n_328) );
OR2x2_ASAP7_75t_L g352 ( .A(n_135), .B(n_167), .Y(n_352) );
OR2x2_ASAP7_75t_L g360 ( .A(n_135), .B(n_259), .Y(n_360) );
AND2x2_ASAP7_75t_L g363 ( .A(n_135), .B(n_186), .Y(n_363) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g257 ( .A(n_136), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g271 ( .A(n_136), .B(n_186), .Y(n_271) );
AND2x2_ASAP7_75t_L g321 ( .A(n_136), .B(n_259), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_136), .B(n_167), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_136), .B(n_420), .Y(n_441) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_164), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_137), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g209 ( .A(n_137), .Y(n_209) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_137), .A2(n_260), .B(n_267), .Y(n_259) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_139), .B(n_140), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B1(n_160), .B2(n_161), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_144), .A2(n_174), .B(n_175), .C(n_176), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_144), .A2(n_175), .B(n_189), .C(n_190), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_144), .A2(n_175), .B(n_242), .C(n_243), .Y(n_241) );
INVx4_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_145), .B(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g172 ( .A(n_145), .B(n_162), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_145), .A2(n_476), .B(n_479), .Y(n_475) );
BUFx3_ASAP7_75t_L g495 ( .A(n_145), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_145), .A2(n_502), .B(n_506), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_145), .A2(n_523), .B(n_526), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_145), .A2(n_539), .B(n_543), .Y(n_538) );
INVx2_ASAP7_75t_L g266 ( .A(n_148), .Y(n_266) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVx1_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_154), .B1(n_155), .B2(n_156), .Y(n_151) );
INVx2_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx4_ASAP7_75t_L g244 ( .A(n_152), .Y(n_244) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
AND2x2_ASAP7_75t_L g162 ( .A(n_153), .B(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
INVx3_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
INVx1_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
INVx5_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
BUFx3_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
INVx1_ASAP7_75t_L g535 ( .A(n_158), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_161), .A2(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_161), .A2(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g482 ( .A(n_163), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_166), .A2(n_360), .B(n_361), .C(n_364), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_166), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_166), .B(n_304), .Y(n_426) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_186), .Y(n_166) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_167), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
AND2x2_ASAP7_75t_L g311 ( .A(n_167), .B(n_305), .Y(n_311) );
INVx1_ASAP7_75t_SL g319 ( .A(n_167), .Y(n_319) );
AND2x2_ASAP7_75t_L g342 ( .A(n_167), .B(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g420 ( .A(n_167), .Y(n_420) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_184), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g210 ( .A(n_169), .B(n_211), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_169), .B(n_495), .C(n_514), .Y(n_513) );
AO21x1_ASAP7_75t_L g558 ( .A1(n_169), .A2(n_514), .B(n_559), .Y(n_558) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_170), .A2(n_187), .B(n_194), .Y(n_186) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_170), .A2(n_475), .B(n_484), .Y(n_474) );
BUFx2_ASAP7_75t_L g240 ( .A(n_172), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g491 ( .A1(n_177), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_177), .A2(n_544), .B(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx4_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_178), .A2(n_483), .B1(n_515), .B2(n_516), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_178), .A2(n_483), .B1(n_534), .B2(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g553 ( .A1(n_178), .A2(n_181), .B1(n_554), .B2(n_555), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_181), .B(n_193), .Y(n_192) );
INVx5_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_SL g523 ( .A1(n_182), .A2(n_204), .B(n_524), .C(n_525), .Y(n_523) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
INVx1_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
INVx2_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_185), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_185), .A2(n_522), .B(n_529), .Y(n_521) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_185), .A2(n_538), .B(n_546), .Y(n_537) );
BUFx2_ASAP7_75t_L g256 ( .A(n_186), .Y(n_256) );
INVx1_ASAP7_75t_L g318 ( .A(n_186), .Y(n_318) );
INVx3_ASAP7_75t_L g343 ( .A(n_186), .Y(n_343) );
INVx1_ASAP7_75t_L g542 ( .A(n_191), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_195), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_223), .Y(n_195) );
INVx1_ASAP7_75t_L g339 ( .A(n_196), .Y(n_339) );
OAI32xp33_ASAP7_75t_L g345 ( .A1(n_196), .A2(n_284), .A3(n_346), .B1(n_347), .B2(n_348), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_196), .A2(n_350), .B1(n_353), .B2(n_358), .Y(n_349) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g287 ( .A(n_197), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g365 ( .A(n_197), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g435 ( .A(n_197), .B(n_381), .Y(n_435) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_212), .Y(n_197) );
AND2x2_ASAP7_75t_L g250 ( .A(n_198), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g280 ( .A(n_198), .Y(n_280) );
INVx1_ASAP7_75t_L g299 ( .A(n_198), .Y(n_299) );
OR2x2_ASAP7_75t_L g307 ( .A(n_198), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g314 ( .A(n_198), .B(n_288), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_198), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g335 ( .A(n_198), .B(n_253), .Y(n_335) );
INVx3_ASAP7_75t_L g357 ( .A(n_198), .Y(n_357) );
AND2x2_ASAP7_75t_L g382 ( .A(n_198), .B(n_254), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_198), .B(n_347), .Y(n_430) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_210), .Y(n_198) );
AOI21xp5_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_201), .B(n_209), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B(n_206), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_204), .A2(n_264), .B(n_265), .C(n_266), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_204), .A2(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g483 ( .A(n_204), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_204), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_206), .A2(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g247 ( .A(n_208), .Y(n_247) );
INVx1_ASAP7_75t_L g219 ( .A(n_209), .Y(n_219) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_209), .A2(n_487), .B(n_496), .Y(n_486) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_209), .A2(n_501), .B(n_509), .Y(n_500) );
INVx2_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
AND2x2_ASAP7_75t_L g386 ( .A(n_212), .B(n_224), .Y(n_386) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_220), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_222), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_222), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g428 ( .A(n_223), .Y(n_428) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
INVx1_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
AND2x2_ASAP7_75t_L g300 ( .A(n_224), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_224), .B(n_254), .Y(n_308) );
AND2x2_ASAP7_75t_L g366 ( .A(n_224), .B(n_289), .Y(n_366) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g252 ( .A(n_225), .Y(n_252) );
AND2x2_ASAP7_75t_L g279 ( .A(n_225), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g288 ( .A(n_225), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_225), .B(n_254), .Y(n_354) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_237), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_237), .B(n_254), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_237), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g381 ( .A(n_237), .Y(n_381) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g253 ( .A(n_238), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g289 ( .A(n_238), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g505 ( .A(n_244), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_244), .A2(n_527), .B(n_528), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_249), .A2(n_259), .B1(n_418), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OAI21xp5_ASAP7_75t_SL g440 ( .A1(n_251), .A2(n_362), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_252), .B(n_357), .Y(n_374) );
INVx1_ASAP7_75t_L g399 ( .A(n_252), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_253), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g326 ( .A(n_253), .B(n_279), .Y(n_326) );
INVx2_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
INVx1_ASAP7_75t_L g332 ( .A(n_254), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_255), .A2(n_407), .B1(n_424), .B2(n_427), .C(n_429), .Y(n_423) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g294 ( .A(n_256), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_256), .B(n_305), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_257), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g348 ( .A(n_257), .B(n_294), .Y(n_348) );
INVx3_ASAP7_75t_SL g389 ( .A(n_257), .Y(n_389) );
AND2x2_ASAP7_75t_L g333 ( .A(n_258), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g362 ( .A(n_258), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_258), .B(n_271), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_258), .B(n_317), .Y(n_403) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
OAI322xp33_ASAP7_75t_L g400 ( .A1(n_259), .A2(n_331), .A3(n_353), .B1(n_401), .B2(n_403), .C1(n_404), .C2(n_405), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_266), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_270), .A2(n_273), .B(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_SL g350 ( .A(n_271), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g372 ( .A(n_271), .B(n_284), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_271), .B(n_311), .Y(n_387) );
INVxp67_ASAP7_75t_L g338 ( .A(n_273), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_273), .A2(n_345), .B(n_349), .C(n_359), .Y(n_344) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_283), .B1(n_286), .B2(n_290), .C(n_295), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g415 ( .A(n_282), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_283), .A2(n_432), .B1(n_437), .B2(n_438), .C(n_440), .Y(n_431) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_284), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g331 ( .A(n_284), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_284), .B(n_362), .Y(n_369) );
AND2x2_ASAP7_75t_L g411 ( .A(n_284), .B(n_389), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_285), .B(n_310), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_285), .A2(n_297), .B1(n_407), .B2(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g437 ( .A(n_285), .B(n_305), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g414 ( .A(n_288), .Y(n_414) );
AND2x2_ASAP7_75t_L g439 ( .A(n_288), .B(n_382), .Y(n_439) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_SL g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g303 ( .A(n_293), .B(n_304), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_302), .B1(n_306), .B2(n_309), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g370 ( .A(n_298), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_298), .B(n_338), .Y(n_405) );
AOI322xp5_ASAP7_75t_L g329 ( .A1(n_300), .A2(n_330), .A3(n_332), .B1(n_333), .B2(n_335), .C1(n_336), .C2(n_340), .Y(n_329) );
INVxp67_ASAP7_75t_L g323 ( .A(n_301), .Y(n_323) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_303), .A2(n_308), .B1(n_325), .B2(n_327), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_304), .B(n_317), .Y(n_404) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_305), .B(n_343), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_305), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g401 ( .A(n_307), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
NAND3xp33_ASAP7_75t_SL g312 ( .A(n_313), .B(n_329), .C(n_344), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_320), .B2(n_322), .C(n_324), .Y(n_313) );
AND2x2_ASAP7_75t_L g320 ( .A(n_316), .B(n_321), .Y(n_320) );
INVx3_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g330 ( .A(n_321), .B(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_323), .Y(n_402) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_328), .B(n_342), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_331), .B(n_389), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_332), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g407 ( .A(n_335), .Y(n_407) );
AND2x2_ASAP7_75t_L g422 ( .A(n_335), .B(n_399), .Y(n_422) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_346), .A2(n_417), .B(n_423), .C(n_431), .Y(n_416) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_386), .Y(n_385) );
NAND2x1_ASAP7_75t_SL g427 ( .A(n_357), .B(n_428), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_360), .Y(n_397) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
AND2x2_ASAP7_75t_L g396 ( .A(n_366), .B(n_382), .Y(n_396) );
NOR5xp2_ASAP7_75t_L g367 ( .A(n_368), .B(n_383), .C(n_400), .D(n_406), .E(n_409), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_373), .C(n_375), .Y(n_368) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_372), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g398 ( .A(n_382), .B(n_399), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_387), .B1(n_388), .B2(n_390), .C(n_393), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B1(n_397), .B2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
AOI211xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_412), .B(n_414), .C(n_415), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g450 ( .A(n_445), .Y(n_450) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_446), .B(n_750), .Y(n_751) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g749 ( .A(n_447), .B(n_750), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_449), .B(n_452), .C(n_755), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g753 ( .A(n_467), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g467 ( .A(n_468), .B(n_671), .Y(n_467) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_469), .B(n_629), .Y(n_468) );
NOR4xp25_ASAP7_75t_L g469 ( .A(n_470), .B(n_569), .C(n_605), .D(n_619), .Y(n_469) );
OAI221xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_517), .B1(n_547), .B2(n_556), .C(n_560), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_471), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_497), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_485), .Y(n_473) );
AND2x2_ASAP7_75t_L g566 ( .A(n_474), .B(n_486), .Y(n_566) );
INVx3_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g628 ( .A(n_474), .B(n_500), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_474), .B(n_499), .Y(n_664) );
AND2x2_ASAP7_75t_L g722 ( .A(n_474), .B(n_584), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_483), .Y(n_479) );
INVx2_ASAP7_75t_L g493 ( .A(n_482), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_483), .A2(n_493), .B(n_507), .C(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g557 ( .A(n_485), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g571 ( .A(n_485), .B(n_500), .Y(n_571) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_486), .B(n_500), .Y(n_586) );
AND2x2_ASAP7_75t_L g598 ( .A(n_486), .B(n_574), .Y(n_598) );
OR2x2_ASAP7_75t_L g600 ( .A(n_486), .B(n_558), .Y(n_600) );
AND2x2_ASAP7_75t_L g635 ( .A(n_486), .B(n_558), .Y(n_635) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_486), .Y(n_680) );
INVx1_ASAP7_75t_L g688 ( .A(n_486), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_491), .B(n_495), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_497), .A2(n_606), .B1(n_610), .B2(n_614), .C(n_615), .Y(n_605) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
INVx2_ASAP7_75t_L g564 ( .A(n_499), .Y(n_564) );
AND2x2_ASAP7_75t_L g617 ( .A(n_499), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g636 ( .A(n_499), .B(n_574), .Y(n_636) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g699 ( .A(n_500), .B(n_574), .Y(n_699) );
AND2x2_ASAP7_75t_L g621 ( .A(n_510), .B(n_566), .Y(n_621) );
OAI322xp33_ASAP7_75t_L g689 ( .A1(n_510), .A2(n_645), .A3(n_690), .B1(n_692), .B2(n_695), .C1(n_697), .C2(n_701), .Y(n_689) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_511), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g585 ( .A(n_511), .Y(n_585) );
AND2x2_ASAP7_75t_L g694 ( .A(n_511), .B(n_574), .Y(n_694) );
AND2x2_ASAP7_75t_L g726 ( .A(n_511), .B(n_598), .Y(n_726) );
OR2x2_ASAP7_75t_L g729 ( .A(n_511), .B(n_730), .Y(n_729) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g559 ( .A(n_512), .Y(n_559) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
INVx1_ASAP7_75t_L g742 ( .A(n_519), .Y(n_742) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g549 ( .A(n_520), .B(n_537), .Y(n_549) );
INVx2_ASAP7_75t_L g582 ( .A(n_520), .Y(n_582) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g604 ( .A(n_521), .Y(n_604) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_521), .Y(n_612) );
OR2x2_ASAP7_75t_L g736 ( .A(n_521), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g561 ( .A(n_530), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g601 ( .A(n_530), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g653 ( .A(n_530), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_537), .Y(n_530) );
AND2x2_ASAP7_75t_L g550 ( .A(n_531), .B(n_551), .Y(n_550) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_531), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g662 ( .A(n_531), .B(n_552), .Y(n_662) );
OR2x2_ASAP7_75t_L g670 ( .A(n_531), .B(n_604), .Y(n_670) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g579 ( .A(n_532), .Y(n_579) );
AND2x2_ASAP7_75t_L g589 ( .A(n_532), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g613 ( .A(n_532), .B(n_537), .Y(n_613) );
AND2x2_ASAP7_75t_L g677 ( .A(n_532), .B(n_552), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_537), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_537), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g590 ( .A(n_537), .Y(n_590) );
INVx1_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
AND2x2_ASAP7_75t_L g607 ( .A(n_537), .B(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_537), .Y(n_685) );
INVx1_ASAP7_75t_L g737 ( .A(n_537), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_542), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g714 ( .A(n_548), .B(n_623), .Y(n_714) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g641 ( .A(n_550), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g740 ( .A(n_550), .B(n_675), .Y(n_740) );
INVx1_ASAP7_75t_L g562 ( .A(n_551), .Y(n_562) );
AND2x2_ASAP7_75t_L g588 ( .A(n_551), .B(n_582), .Y(n_588) );
BUFx2_ASAP7_75t_L g647 ( .A(n_551), .Y(n_647) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_552), .Y(n_568) );
INVx1_ASAP7_75t_L g578 ( .A(n_552), .Y(n_578) );
NOR2xp67_ASAP7_75t_L g716 ( .A(n_556), .B(n_563), .Y(n_716) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI32xp33_ASAP7_75t_L g560 ( .A1(n_557), .A2(n_561), .A3(n_563), .B1(n_565), .B2(n_567), .Y(n_560) );
AND2x2_ASAP7_75t_L g700 ( .A(n_557), .B(n_573), .Y(n_700) );
AND2x2_ASAP7_75t_L g738 ( .A(n_557), .B(n_636), .Y(n_738) );
INVx1_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_562), .B(n_624), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_563), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_563), .B(n_566), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_563), .B(n_635), .Y(n_717) );
OR2x2_ASAP7_75t_L g731 ( .A(n_563), .B(n_600), .Y(n_731) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g658 ( .A(n_564), .B(n_566), .Y(n_658) );
OR2x2_ASAP7_75t_L g667 ( .A(n_564), .B(n_654), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_566), .B(n_617), .Y(n_639) );
INVx2_ASAP7_75t_L g654 ( .A(n_568), .Y(n_654) );
OR2x2_ASAP7_75t_L g669 ( .A(n_568), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g684 ( .A(n_568), .B(n_685), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_568), .A2(n_661), .B(n_742), .C(n_743), .Y(n_741) );
OAI321xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_575), .A3(n_580), .B1(n_583), .B2(n_587), .C(n_591), .Y(n_569) );
INVx1_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g693 ( .A(n_571), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g645 ( .A(n_573), .Y(n_645) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_574), .B(n_688), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_575), .A2(n_713), .B1(n_715), .B2(n_717), .C(n_718), .Y(n_712) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
AND2x2_ASAP7_75t_L g650 ( .A(n_577), .B(n_624), .Y(n_650) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_578), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g623 ( .A(n_579), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_580), .A2(n_621), .B(n_666), .C(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g632 ( .A(n_582), .B(n_589), .Y(n_632) );
BUFx2_ASAP7_75t_L g642 ( .A(n_582), .Y(n_642) );
INVx1_ASAP7_75t_L g657 ( .A(n_582), .Y(n_657) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g663 ( .A(n_585), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g746 ( .A(n_585), .Y(n_746) );
INVx1_ASAP7_75t_L g739 ( .A(n_586), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g592 ( .A(n_588), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g696 ( .A(n_588), .B(n_613), .Y(n_696) );
INVx1_ASAP7_75t_L g625 ( .A(n_589), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B1(n_599), .B2(n_601), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_593), .B(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g661 ( .A(n_594), .B(n_662), .Y(n_661) );
BUFx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_SL g624 ( .A(n_595), .B(n_604), .Y(n_624) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g616 ( .A(n_598), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g626 ( .A(n_600), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_603), .A2(n_721), .B1(n_723), .B2(n_724), .C(n_725), .Y(n_720) );
INVx1_ASAP7_75t_L g609 ( .A(n_604), .Y(n_609) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_604), .Y(n_675) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_607), .B(n_726), .Y(n_725) );
OAI21xp5_ASAP7_75t_L g615 ( .A1(n_608), .A2(n_613), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_611), .B(n_621), .Y(n_718) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g687 ( .A(n_612), .Y(n_687) );
AND2x2_ASAP7_75t_L g646 ( .A(n_613), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g735 ( .A(n_613), .Y(n_735) );
INVx1_ASAP7_75t_L g651 ( .A(n_616), .Y(n_651) );
INVx1_ASAP7_75t_L g706 ( .A(n_617), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B1(n_625), .B2(n_626), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_623), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g691 ( .A(n_624), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_624), .B(n_662), .Y(n_728) );
OR2x2_ASAP7_75t_L g701 ( .A(n_625), .B(n_654), .Y(n_701) );
INVx1_ASAP7_75t_L g640 ( .A(n_626), .Y(n_640) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_628), .B(n_679), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_648), .C(n_659), .Y(n_629) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B(n_637), .C(n_643), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_632), .A2(n_703), .B1(n_707), .B2(n_710), .C(n_712), .Y(n_702) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
AND2x2_ASAP7_75t_L g644 ( .A(n_635), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g698 ( .A(n_635), .B(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g683 ( .A1(n_636), .A2(n_684), .B(n_686), .C(n_688), .Y(n_683) );
INVx2_ASAP7_75t_L g730 ( .A(n_636), .Y(n_730) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_640), .B(n_641), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g709 ( .A(n_642), .B(n_662), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_651), .B(n_652), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_655), .B(n_658), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_653), .B(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_658), .B(n_745), .Y(n_744) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_665), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g686 ( .A(n_662), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND4x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_702), .C(n_719), .D(n_741), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_689), .Y(n_672) );
OAI211xp5_ASAP7_75t_SL g673 ( .A1(n_674), .A2(n_678), .B(n_681), .C(n_683), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_677), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_688), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g723 ( .A(n_698), .Y(n_723) );
INVx2_ASAP7_75t_SL g711 ( .A(n_699), .Y(n_711) );
OR2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g724 ( .A(n_709), .Y(n_724) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_727), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
OAI221xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_732), .C(n_733), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g754 ( .A(n_748), .Y(n_754) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule