module fake_aes_10208_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_3), .B(n_1), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_10), .B(n_1), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_7), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_16), .B(n_0), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_17), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_15), .B(n_2), .Y(n_21) );
OA21x2_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_13), .B(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_20), .B1(n_19), .B2(n_14), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_22), .Y(n_26) );
NAND2xp33_ASAP7_75t_SL g27 ( .A(n_25), .B(n_14), .Y(n_27) );
NOR2xp33_ASAP7_75t_SL g28 ( .A(n_26), .B(n_13), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_22), .B1(n_23), .B2(n_19), .Y(n_29) );
INVxp67_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
AOI322xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_19), .A3(n_18), .B1(n_3), .B2(n_4), .C1(n_5), .C2(n_22), .Y(n_31) );
A2O1A1Ixp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_18), .B(n_22), .C(n_5), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_8), .B1(n_9), .B2(n_11), .C1(n_22), .C2(n_32), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
INVx4_ASAP7_75t_L g35 ( .A(n_31), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_35), .B(n_22), .Y(n_36) );
BUFx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
AOI22x1_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_33), .B1(n_34), .B2(n_36), .Y(n_39) );
endmodule