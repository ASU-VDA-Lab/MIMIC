module fake_jpeg_13822_n_197 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_25),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_11),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_68),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_26),
.C(n_48),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_84),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_64),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_76),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_58),
.B1(n_66),
.B2(n_74),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_58),
.B1(n_66),
.B2(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_109),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_77),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_117),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_73),
.B1(n_75),
.B2(n_74),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_73),
.B1(n_75),
.B2(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_67),
.B1(n_62),
.B2(n_63),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_71),
.B1(n_72),
.B2(n_60),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_125),
.Y(n_137)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_65),
.B1(n_59),
.B2(n_81),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_87),
.B1(n_56),
.B2(n_31),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_65),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_22),
.C(n_47),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_117),
.Y(n_142)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_142),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_81),
.A3(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_6),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_10),
.B(n_12),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_42),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_115),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_29),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_150),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_2),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_5),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_32),
.C(n_44),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_127),
.B(n_5),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_7),
.B(n_10),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_139),
.B1(n_132),
.B2(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_162),
.Y(n_176)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_164),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_37),
.C(n_43),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_150),
.C(n_140),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_167),
.A2(n_13),
.B(n_16),
.Y(n_177)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_175),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_177),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_144),
.C(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

AOI221xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_159),
.B1(n_161),
.B2(n_168),
.C(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_185),
.B1(n_176),
.B2(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_156),
.C(n_170),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_180),
.B1(n_181),
.B2(n_186),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_182),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_192),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_154),
.C(n_163),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_160),
.B1(n_35),
.B2(n_38),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_18),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_39),
.Y(n_197)
);


endmodule