module real_jpeg_26346_n_6 (n_5, n_4, n_36, n_0, n_37, n_1, n_2, n_33, n_34, n_35, n_3, n_6);

input n_5;
input n_4;
input n_36;
input n_0;
input n_37;
input n_1;
input n_2;
input n_33;
input n_34;
input n_35;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

FAx1_ASAP7_75t_SL g6 ( 
.A(n_0),
.B(n_7),
.CI(n_11),
.CON(n_6),
.SN(n_6)
);

INVx6_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_14),
.C(n_24),
.Y(n_13)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_16),
.Y(n_15)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_9),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g9 ( 
.A(n_10),
.Y(n_9)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_27),
.C(n_28),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_19),
.C(n_20),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_33),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_34),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_35),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_36),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_37),
.Y(n_30)
);


endmodule