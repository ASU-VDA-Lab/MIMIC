module real_jpeg_32656_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_1),
.A2(n_339),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_1),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_66),
.B2(n_68),
.Y(n_60)
);

INVx2_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_2),
.A2(n_68),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_2),
.A2(n_68),
.B1(n_273),
.B2(n_277),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g421 ( 
.A1(n_2),
.A2(n_68),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_3),
.A2(n_37),
.B1(n_114),
.B2(n_120),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_37),
.B1(n_244),
.B2(n_248),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_3),
.A2(n_37),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_4),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_4),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_4),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_6),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_7),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_7),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_7),
.A2(n_285),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_9),
.A2(n_97),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_9),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_9),
.A2(n_139),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_9),
.A2(n_139),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_10),
.A2(n_155),
.B1(n_261),
.B2(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_10),
.A2(n_155),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_13),
.A2(n_406),
.B1(n_408),
.B2(n_411),
.Y(n_405)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_13),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_14),
.Y(n_209)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_14),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_14),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_15),
.A2(n_194),
.B1(n_199),
.B2(n_200),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_15),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_15),
.A2(n_199),
.B1(n_376),
.B2(n_378),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_28),
.B1(n_38),
.B2(n_43),
.Y(n_27)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_16),
.A2(n_203),
.A3(n_205),
.B1(n_210),
.B2(n_215),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_16),
.A2(n_51),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_16),
.B(n_330),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_16),
.A2(n_329),
.B(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_391),
.B1(n_434),
.B2(n_435),
.Y(n_18)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_19),
.Y(n_435)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_304),
.B(n_390),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_253),
.B(n_303),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_182),
.B(n_252),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_145),
.Y(n_23)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_81),
.B(n_142),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_58),
.B(n_80),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_49),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_28),
.A2(n_43),
.B1(n_60),
.B2(n_69),
.Y(n_59)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_32),
.Y(n_341)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_32),
.Y(n_410)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_42),
.Y(n_149)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_42),
.Y(n_415)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_43),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_43),
.A2(n_137),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_43),
.A2(n_338),
.B1(n_405),
.B2(n_412),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_46),
.Y(n_192)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_46),
.Y(n_336)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_48),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_93),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_SL g125 ( 
.A1(n_51),
.A2(n_92),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_51),
.B(n_211),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_R g289 ( 
.A(n_51),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_53),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_71),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_71),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_64),
.Y(n_287)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_72),
.A2(n_130),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_72),
.A2(n_130),
.B1(n_260),
.B2(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_72),
.A2(n_130),
.B1(n_375),
.B2(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AO21x2_ASAP7_75t_L g130 ( 
.A1(n_73),
.A2(n_102),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_135),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_110),
.B1(n_111),
.B2(n_134),
.Y(n_82)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_83),
.B(n_110),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_91),
.B1(n_96),
.B2(n_101),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_106),
.Y(n_382)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_110),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_134),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_125),
.B2(n_129),
.Y(n_111)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_162),
.Y(n_161)
);

AOI22x1_ASAP7_75t_L g224 ( 
.A1(n_112),
.A2(n_129),
.B1(n_162),
.B2(n_225),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_129),
.Y(n_160)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_124),
.Y(n_264)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_140),
.A2(n_151),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_140),
.A2(n_193),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_140),
.A2(n_284),
.B1(n_334),
.B2(n_337),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_183),
.B(n_184),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_159),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_169),
.C(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B(n_169),
.C(n_181),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_161),
.C(n_169),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_R g186 ( 
.A(n_160),
.B(n_161),
.Y(n_186)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_165),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_167),
.Y(n_266)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_168),
.Y(n_403)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AO21x2_ASAP7_75t_L g230 ( 
.A1(n_171),
.A2(n_215),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_178),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_172),
.Y(n_377)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2x1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_187),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_222),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_188),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_202),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_189),
.B(n_202),
.Y(n_257)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_SL g241 ( 
.A(n_207),
.Y(n_241)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_208),
.Y(n_430)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_217),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_224),
.B(n_228),
.C(n_302),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_230),
.A2(n_242),
.B1(n_243),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_230),
.A2(n_242),
.B1(n_272),
.B2(n_384),
.Y(n_383)
);

OA22x2_ASAP7_75t_L g428 ( 
.A1(n_230),
.A2(n_242),
.B1(n_384),
.B2(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_244),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_246),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_301),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_301),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_269),
.B2(n_270),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_267),
.B2(n_268),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_258),
.B(n_268),
.C(n_269),
.Y(n_389)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_280),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_271),
.B(n_289),
.C(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_279),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

BUFx4f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_290),
.A2(n_352),
.B1(n_356),
.B2(n_367),
.Y(n_351)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_290),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_295),
.B1(n_299),
.B2(n_300),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_389),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_305),
.B(n_389),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_349),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_347),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_307),
.B(n_347),
.C(n_349),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_333),
.B1(n_345),
.B2(n_346),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_308),
.B(n_346),
.Y(n_417)
);

OAI32xp33_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_311),
.A3(n_314),
.B1(n_321),
.B2(n_328),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_318),
.Y(n_359)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_319),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_341),
.Y(n_344)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

BUFx2_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_373),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_SL g396 ( 
.A(n_351),
.B(n_374),
.C(n_383),
.Y(n_396)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_357),
.A2(n_420),
.B1(n_421),
.B2(n_427),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_364),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_366),
.Y(n_372)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_367),
.Y(n_427)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_391),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_432),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_393),
.B(n_394),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_416),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_404),
.Y(n_397)
);

BUFx6f_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_428),
.Y(n_418)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);


endmodule