module fake_jpeg_1315_n_210 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_210);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g69 ( 
.A(n_14),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_81),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_62),
.B1(n_61),
.B2(n_63),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_80),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_56),
.B1(n_53),
.B2(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_93),
.B1(n_66),
.B2(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_66),
.B1(n_72),
.B2(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_98),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_57),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_71),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_33),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_74),
.B(n_79),
.Y(n_116)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_111),
.B1(n_75),
.B2(n_77),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_65),
.B(n_58),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_121),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_108),
.C(n_110),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_133),
.C(n_51),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_78),
.B1(n_90),
.B2(n_53),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_73),
.B1(n_52),
.B2(n_22),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_90),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_54),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_1),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_98),
.B1(n_79),
.B2(n_59),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_74),
.B1(n_73),
.B2(n_52),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_73),
.C(n_52),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_3),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_20),
.B1(n_50),
.B2(n_47),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_151),
.B1(n_27),
.B2(n_39),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_4),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_150),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_19),
.B1(n_42),
.B2(n_40),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_120),
.B(n_26),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_8),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_156),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_153),
.C(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_169),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_131),
.B(n_129),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_156),
.B(n_151),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_174),
.B1(n_146),
.B2(n_142),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_170),
.B(n_140),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_9),
.B(n_10),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_31),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_182),
.Y(n_190)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_165),
.B(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_185),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_152),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_168),
.B1(n_176),
.B2(n_165),
.Y(n_187)
);

AO221x1_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_185),
.B1(n_167),
.B2(n_178),
.C(n_180),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_162),
.B1(n_159),
.B2(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_185),
.C(n_32),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_158),
.C(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_198),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_193),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_192),
.B1(n_196),
.B2(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_203),
.B(n_201),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_200),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_186),
.A3(n_17),
.B1(n_34),
.B2(n_44),
.C1(n_38),
.C2(n_37),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_12),
.B(n_13),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_13),
.B(n_14),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_15),
.Y(n_210)
);


endmodule