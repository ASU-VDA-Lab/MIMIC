module fake_netlist_1_2736_n_477 (n_117, n_44, n_133, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_139, n_16, n_13, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_132, n_51, n_140, n_96, n_39, n_477);
input n_117;
input n_44;
input n_133;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_139;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_51;
input n_140;
input n_96;
input n_39;
output n_477;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_431;
wire n_161;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_245;
wire n_357;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g143 ( .A(n_32), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_24), .Y(n_144) );
BUFx2_ASAP7_75t_L g145 ( .A(n_46), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_71), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_37), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_64), .Y(n_148) );
INVxp67_ASAP7_75t_SL g149 ( .A(n_68), .Y(n_149) );
INVxp33_ASAP7_75t_L g150 ( .A(n_79), .Y(n_150) );
INVxp33_ASAP7_75t_L g151 ( .A(n_78), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_35), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_72), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_48), .Y(n_154) );
BUFx5_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_117), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_14), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_67), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_84), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_22), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_27), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_75), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_121), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_77), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_96), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_97), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_106), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_38), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_76), .Y(n_172) );
INVxp33_ASAP7_75t_L g173 ( .A(n_25), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_105), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_98), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_83), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_110), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_93), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_62), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_142), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_94), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_17), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_55), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_34), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_123), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_116), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_60), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_58), .Y(n_189) );
CKINVDCx14_ASAP7_75t_R g190 ( .A(n_129), .Y(n_190) );
INVxp33_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_61), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_119), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_90), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_111), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_45), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_6), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_19), .Y(n_199) );
BUFx5_ASAP7_75t_L g200 ( .A(n_13), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_26), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_23), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_138), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_99), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_15), .Y(n_206) );
CKINVDCx14_ASAP7_75t_R g207 ( .A(n_115), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_51), .Y(n_208) );
BUFx2_ASAP7_75t_SL g209 ( .A(n_101), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_13), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_44), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_44), .Y(n_212) );
BUFx2_ASAP7_75t_SL g213 ( .A(n_120), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_200), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_196), .B(n_0), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_145), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_200), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_168), .B(n_1), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_155), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_195), .B(n_2), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_201), .B(n_2), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_155), .B(n_3), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_167), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_167), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_167), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_150), .B(n_3), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_173), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_144), .B(n_4), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_159), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_169), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_143), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_173), .B(n_5), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_171), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_240) );
INVx5_ASAP7_75t_L g241 ( .A(n_169), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_153), .A2(n_54), .B(n_53), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_153), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_203), .B(n_7), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_234), .B(n_211), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_214), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
CKINVDCx8_ASAP7_75t_R g249 ( .A(n_218), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_229), .Y(n_250) );
OR2x6_ASAP7_75t_L g251 ( .A(n_239), .B(n_209), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_234), .B(n_151), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_218), .B(n_191), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_216), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_226), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_216), .B(n_162), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_239), .B(n_190), .Y(n_259) );
BUFx10_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_239), .B(n_190), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_226), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_226), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_226), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_238), .B(n_160), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_226), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_152), .B1(n_154), .B2(n_147), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_230), .Y(n_273) );
OR2x6_ASAP7_75t_L g274 ( .A(n_240), .B(n_213), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_223), .B(n_207), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_215), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_259), .B(n_223), .Y(n_277) );
INVx4_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_261), .B(n_225), .Y(n_279) );
INVx4_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_266), .B(n_225), .Y(n_281) );
INVxp67_ASAP7_75t_SL g282 ( .A(n_252), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_275), .B(n_227), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_275), .B(n_227), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_254), .B(n_220), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_260), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_249), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_246), .B(n_245), .Y(n_290) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_266), .B(n_184), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_260), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_260), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_246), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_257), .B(n_238), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_270), .B(n_204), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g297 ( .A(n_257), .B(n_233), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_268), .A2(n_243), .B(n_221), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_251), .B(n_163), .Y(n_299) );
NOR2xp33_ASAP7_75t_SL g300 ( .A(n_274), .B(n_158), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_248), .Y(n_302) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_247), .B(n_148), .Y(n_303) );
BUFx8_ASAP7_75t_L g304 ( .A(n_250), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_258), .A2(n_243), .B(n_228), .Y(n_305) );
NOR2xp33_ASAP7_75t_SL g306 ( .A(n_258), .B(n_166), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_256), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_263), .B(n_236), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_305), .B(n_219), .C(n_217), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_298), .A2(n_222), .B(n_219), .Y(n_311) );
INVx4_ASAP7_75t_L g312 ( .A(n_278), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_277), .A2(n_224), .B(n_170), .Y(n_313) );
AND2x6_ASAP7_75t_L g314 ( .A(n_292), .B(n_182), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_279), .A2(n_149), .B(n_264), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_280), .B(n_236), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_290), .B(n_185), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_283), .A2(n_267), .B(n_264), .Y(n_318) );
AOI22x1_ASAP7_75t_L g319 ( .A1(n_305), .A2(n_244), .B1(n_231), .B2(n_237), .Y(n_319) );
O2A1O1Ixp5_ASAP7_75t_L g320 ( .A1(n_285), .A2(n_161), .B(n_165), .C(n_160), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_292), .B(n_164), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_284), .A2(n_269), .B(n_267), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_289), .B(n_299), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_295), .A2(n_271), .B(n_146), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_300), .A2(n_244), .B1(n_202), .B2(n_206), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_302), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_302), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_296), .A2(n_212), .B(n_210), .C(n_197), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_287), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_291), .A2(n_244), .B1(n_156), .B2(n_157), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_301), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_281), .A2(n_198), .B1(n_208), .B2(n_199), .Y(n_333) );
NOR2xp33_ASAP7_75t_SL g334 ( .A(n_306), .B(n_172), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_297), .B(n_181), .Y(n_335) );
INVx4_ASAP7_75t_L g336 ( .A(n_286), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_288), .B(n_183), .Y(n_337) );
NOR2xp67_ASAP7_75t_L g338 ( .A(n_308), .B(n_8), .Y(n_338) );
OAI21xp33_ASAP7_75t_L g339 ( .A1(n_303), .A2(n_176), .B(n_174), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_307), .A2(n_178), .B(n_179), .C(n_177), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_298), .A2(n_187), .B(n_186), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_298), .A2(n_189), .B(n_188), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_294), .B(n_192), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_282), .A2(n_194), .B(n_193), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_304), .B(n_205), .Y(n_345) );
AO31x2_ASAP7_75t_L g346 ( .A1(n_341), .A2(n_232), .A3(n_237), .B(n_231), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_320), .A2(n_180), .B(n_175), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_331), .A2(n_241), .B1(n_242), .B2(n_230), .Y(n_348) );
AO31x2_ASAP7_75t_L g349 ( .A1(n_342), .A2(n_242), .A3(n_230), .B(n_241), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_SL g350 ( .A1(n_340), .A2(n_57), .B(n_59), .C(n_56), .Y(n_350) );
AO32x2_ASAP7_75t_L g351 ( .A1(n_333), .A2(n_242), .A3(n_12), .B1(n_10), .B2(n_11), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_310), .A2(n_241), .B(n_63), .Y(n_352) );
AOI31xp67_ASAP7_75t_L g353 ( .A1(n_327), .A2(n_256), .A3(n_265), .B(n_262), .Y(n_353) );
OAI22x1_ASAP7_75t_L g354 ( .A1(n_325), .A2(n_18), .B1(n_16), .B2(n_17), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_334), .B(n_241), .Y(n_355) );
AO31x2_ASAP7_75t_L g356 ( .A1(n_311), .A2(n_265), .A3(n_272), .B(n_262), .Y(n_356) );
AOI31xp67_ASAP7_75t_L g357 ( .A1(n_328), .A2(n_272), .A3(n_273), .B(n_265), .Y(n_357) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_344), .A2(n_272), .B(n_273), .C(n_265), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_329), .A2(n_273), .B(n_272), .C(n_21), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_323), .B(n_20), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_318), .A2(n_66), .B(n_65), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_317), .B(n_28), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_324), .A2(n_70), .B(n_69), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_343), .B(n_28), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_322), .A2(n_74), .B(n_73), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_SL g369 ( .A1(n_345), .A2(n_95), .B(n_141), .C(n_140), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_337), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_338), .A2(n_81), .B(n_80), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_330), .A2(n_85), .B(n_82), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_315), .A2(n_87), .B(n_86), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_313), .A2(n_89), .B(n_88), .Y(n_375) );
AOI221x1_ASAP7_75t_L g376 ( .A1(n_339), .A2(n_29), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_332), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_339), .A2(n_30), .B(n_31), .C(n_33), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_335), .A2(n_92), .B(n_91), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_SL g380 ( .A1(n_321), .A2(n_104), .B(n_135), .C(n_134), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
AO31x2_ASAP7_75t_L g382 ( .A1(n_336), .A2(n_314), .A3(n_326), .B(n_34), .Y(n_382) );
AO21x1_ASAP7_75t_L g383 ( .A1(n_341), .A2(n_107), .B(n_133), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_309), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_309), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_309), .Y(n_386) );
AO21x1_ASAP7_75t_L g387 ( .A1(n_341), .A2(n_103), .B(n_131), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_319), .A2(n_102), .B(n_130), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_359), .A2(n_36), .B(n_38), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_347), .A2(n_39), .B(n_40), .Y(n_390) );
AO31x2_ASAP7_75t_L g391 ( .A1(n_383), .A2(n_41), .A3(n_42), .B(n_43), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_384), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_358), .A2(n_108), .B(n_127), .Y(n_393) );
OA21x2_ASAP7_75t_L g394 ( .A1(n_352), .A2(n_100), .B(n_126), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_385), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_366), .B(n_47), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_388), .A2(n_109), .B(n_124), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_386), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_379), .A2(n_363), .B(n_387), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_370), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_364), .B(n_49), .Y(n_401) );
AO31x2_ASAP7_75t_L g402 ( .A1(n_376), .A2(n_50), .A3(n_51), .B(n_52), .Y(n_402) );
AO31x2_ASAP7_75t_L g403 ( .A1(n_378), .A2(n_348), .A3(n_354), .B(n_361), .Y(n_403) );
AO31x2_ASAP7_75t_L g404 ( .A1(n_367), .A2(n_112), .A3(n_113), .B(n_114), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_360), .A2(n_362), .B(n_365), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_374), .B(n_370), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_368), .A2(n_372), .B(n_373), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_350), .B(n_357), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_371), .A2(n_353), .B(n_355), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_380), .A2(n_369), .B(n_381), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_356), .A2(n_349), .B(n_346), .Y(n_412) );
AO31x2_ASAP7_75t_L g413 ( .A1(n_356), .A2(n_346), .A3(n_349), .B(n_351), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_377), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_382), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_384), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_412), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_415), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_400), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_392), .B(n_395), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_413), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_398), .B(n_416), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_413), .Y(n_423) );
OR2x6_ASAP7_75t_L g424 ( .A(n_401), .B(n_396), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_406), .A2(n_389), .B(n_411), .Y(n_425) );
OR2x6_ASAP7_75t_L g426 ( .A(n_401), .B(n_396), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_405), .B(n_408), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_414), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_402), .Y(n_430) );
AO21x2_ASAP7_75t_L g431 ( .A1(n_409), .A2(n_410), .B(n_399), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_414), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
AOI21xp5_ASAP7_75t_SL g435 ( .A1(n_394), .A2(n_393), .B(n_397), .Y(n_435) );
AOI21xp5_ASAP7_75t_SL g436 ( .A1(n_394), .A2(n_393), .B(n_397), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_403), .B(n_404), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_417), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_420), .B(n_422), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_424), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_419), .B(n_427), .Y(n_441) );
INVx5_ASAP7_75t_L g442 ( .A(n_426), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_437), .B(n_434), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_426), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_418), .B(n_429), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_429), .B(n_432), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_432), .B(n_430), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_421), .B(n_423), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_438), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_443), .B(n_431), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_443), .B(n_431), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_439), .B(n_428), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_442), .B(n_433), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_441), .B(n_425), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_449), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_452), .B(n_448), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_450), .B(n_445), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_451), .B(n_447), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_457), .B(n_454), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_457), .B(n_454), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_456), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_455), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_459), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_460), .B(n_461), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_464), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_463), .Y(n_466) );
AOI22x1_ASAP7_75t_L g467 ( .A1(n_465), .A2(n_453), .B1(n_444), .B2(n_440), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_466), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_468), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_469), .B(n_467), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_470), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_471), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_472), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_473), .A2(n_435), .B(n_436), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_474), .B(n_458), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_475), .Y(n_476) );
AOI21xp33_ASAP7_75t_SL g477 ( .A1(n_476), .A2(n_446), .B(n_462), .Y(n_477) );
endmodule