module fake_jpeg_29992_n_468 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_468);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_468;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_SL g49 ( 
.A(n_43),
.Y(n_49)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_54),
.Y(n_101)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_53),
.B(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_14),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_29),
.C(n_31),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_67),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_64),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_0),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_72),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_34),
.B(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_81),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_34),
.B(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_1),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_23),
.A2(n_1),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_3),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_86),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_84),
.B(n_19),
.Y(n_153)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_85),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_42),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_2),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_94),
.Y(n_143)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_96),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_3),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_27),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_32),
.CON(n_103),
.SN(n_103)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_107),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_150),
.B(n_145),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_44),
.B1(n_39),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_130),
.B1(n_136),
.B2(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_17),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_111),
.B(n_68),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_48),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_127),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_58),
.A2(n_45),
.B1(n_44),
.B2(n_39),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_124),
.A2(n_128),
.B1(n_134),
.B2(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_48),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_45),
.B1(n_31),
.B2(n_47),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_31),
.B1(n_19),
.B2(n_35),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_70),
.A2(n_47),
.B1(n_17),
.B2(n_32),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_133),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_83),
.A2(n_30),
.B1(n_33),
.B2(n_26),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_95),
.B1(n_73),
.B2(n_80),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_19),
.B1(n_94),
.B2(n_59),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_89),
.A2(n_30),
.B1(n_33),
.B2(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_153),
.Y(n_175)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_91),
.B(n_19),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_61),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_25),
.B1(n_24),
.B2(n_65),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_154),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_170),
.Y(n_211)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_164),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_197),
.B1(n_202),
.B2(n_141),
.Y(n_208)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_51),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_165),
.B(n_171),
.Y(n_239)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

BUFx4f_ASAP7_75t_SL g210 ( 
.A(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_24),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_185),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_128),
.A2(n_85),
.B1(n_74),
.B2(n_62),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_177),
.B(n_186),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_183),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_111),
.B(n_25),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_182),
.B(n_192),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_135),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_129),
.A2(n_92),
.B1(n_50),
.B2(n_76),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_196),
.B1(n_125),
.B2(n_151),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_127),
.A2(n_91),
.B(n_24),
.C(n_49),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_150),
.B(n_149),
.C(n_131),
.Y(n_226)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_109),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_19),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_134),
.B(n_88),
.C(n_87),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_143),
.Y(n_218)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_129),
.A2(n_86),
.B1(n_56),
.B2(n_55),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_106),
.A2(n_79),
.B1(n_78),
.B2(n_71),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_121),
.B(n_64),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_199),
.Y(n_229)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_142),
.B(n_64),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_113),
.A2(n_86),
.B1(n_56),
.B2(n_55),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_100),
.A2(n_37),
.B1(n_64),
.B2(n_63),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_125),
.B1(n_113),
.B2(n_114),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_204),
.B(n_208),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_150),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_198),
.B(n_201),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_133),
.B(n_107),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_226),
.B(n_233),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_238),
.B1(n_202),
.B2(n_170),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_216),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_103),
.Y(n_219)
);

A2O1A1O1Ixp25_ASAP7_75t_L g268 ( 
.A1(n_219),
.A2(n_244),
.B(n_172),
.C(n_115),
.D(n_98),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_157),
.A2(n_148),
.B1(n_100),
.B2(n_137),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_236),
.B1(n_179),
.B2(n_176),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_173),
.A2(n_149),
.B(n_148),
.C(n_131),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_230),
.B(n_188),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_191),
.A2(n_137),
.B1(n_123),
.B2(n_118),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_123),
.B1(n_118),
.B2(n_104),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_159),
.B(n_110),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_242),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_159),
.B(n_104),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_161),
.B(n_120),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_191),
.Y(n_247)
);

AOI32xp33_ASAP7_75t_L g244 ( 
.A1(n_155),
.A2(n_98),
.A3(n_99),
.B1(n_152),
.B2(n_115),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_262),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_249),
.A2(n_256),
.B1(n_267),
.B2(n_271),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_207),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_252),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_233),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_266),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_160),
.B1(n_181),
.B2(n_177),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_205),
.B(n_160),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_160),
.Y(n_259)
);

AO21x2_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_193),
.B(n_186),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_223),
.B(n_229),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_265),
.B1(n_275),
.B2(n_217),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_205),
.B(n_178),
.C(n_175),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_277),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_232),
.A2(n_185),
.B1(n_194),
.B2(n_163),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_156),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_211),
.A2(n_169),
.B1(n_195),
.B2(n_199),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_209),
.B(n_219),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_189),
.C(n_99),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_269),
.B(n_276),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_207),
.B(n_172),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_211),
.A2(n_184),
.B1(n_183),
.B2(n_174),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_166),
.B1(n_172),
.B2(n_37),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_212),
.B(n_114),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_279),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_208),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_4),
.C(n_6),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_4),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_6),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_242),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_221),
.B(n_7),
.C(n_8),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_209),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_285),
.B(n_293),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_226),
.B1(n_209),
.B2(n_227),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_291),
.B(n_299),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_271),
.B1(n_280),
.B2(n_276),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_290),
.A2(n_301),
.B(n_206),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_230),
.B(n_227),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_229),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_295),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_252),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_298),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_234),
.B(n_236),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_247),
.A2(n_234),
.B(n_224),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_246),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_314),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_272),
.A2(n_235),
.B1(n_220),
.B2(n_215),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_303),
.A2(n_315),
.B(n_210),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_304),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_272),
.A2(n_240),
.B1(n_220),
.B2(n_214),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_261),
.B1(n_265),
.B2(n_275),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_215),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_259),
.A2(n_210),
.B(n_237),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_264),
.C(n_269),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_318),
.C(n_325),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_317),
.A2(n_340),
.B1(n_303),
.B2(n_286),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_289),
.A2(n_256),
.B1(n_260),
.B2(n_249),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_319),
.A2(n_320),
.B1(n_330),
.B2(n_290),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_289),
.A2(n_260),
.B1(n_257),
.B2(n_267),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_322),
.Y(n_346)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_326),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_262),
.C(n_260),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_300),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_260),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_332),
.C(n_338),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_293),
.C(n_298),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_281),
.C(n_268),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_333),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_285),
.Y(n_366)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_278),
.C(n_279),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_206),
.Y(n_339)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_339),
.Y(n_354)
);

AO21x2_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_210),
.B(n_222),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_342),
.A2(n_345),
.B(n_315),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_343),
.Y(n_357)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_317),
.A2(n_286),
.B1(n_294),
.B2(n_282),
.Y(n_351)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_352),
.A2(n_345),
.B1(n_340),
.B2(n_342),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_340),
.A2(n_299),
.B(n_298),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_359),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_335),
.B(n_302),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_365),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_337),
.A2(n_299),
.B(n_290),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_360),
.B(n_366),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_327),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_367),
.B1(n_368),
.B2(n_306),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_328),
.A2(n_294),
.B1(n_282),
.B2(n_302),
.Y(n_363)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_363),
.Y(n_391)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_335),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_328),
.A2(n_288),
.B1(n_284),
.B2(n_303),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_341),
.A2(n_288),
.B1(n_284),
.B2(n_291),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_310),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_320),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_325),
.B(n_318),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_372),
.C(n_332),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_316),
.B(n_338),
.C(n_329),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_352),
.B(n_360),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_362),
.A2(n_369),
.B1(n_365),
.B2(n_354),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_376),
.A2(n_379),
.B1(n_384),
.B2(n_333),
.Y(n_398)
);

AOI21xp33_ASAP7_75t_L g378 ( 
.A1(n_346),
.A2(n_287),
.B(n_340),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_378),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_340),
.B1(n_322),
.B2(n_324),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_382),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_385),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_354),
.A2(n_333),
.B1(n_319),
.B2(n_291),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_312),
.C(n_344),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_312),
.C(n_344),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_388),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_355),
.B(n_295),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_392),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_307),
.Y(n_390)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_390),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_333),
.C(n_343),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_368),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_367),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_370),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_399),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_404),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_370),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_351),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_410),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_371),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_407),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_361),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_363),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_383),
.B1(n_375),
.B2(n_358),
.Y(n_427)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_349),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_413),
.B(n_374),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_400),
.B(n_386),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_416),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_387),
.C(n_386),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_401),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_396),
.B(n_391),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_422),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_377),
.Y(n_420)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_347),
.C(n_384),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_379),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_411),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_347),
.C(n_383),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_426),
.B(n_428),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_427),
.B(n_398),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_307),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_429),
.B(n_437),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_438),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_422),
.A2(n_408),
.B(n_375),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_431),
.A2(n_432),
.B(n_421),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_415),
.A2(n_394),
.B(n_413),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_421),
.B(n_407),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_439),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_417),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_425),
.A2(n_409),
.B1(n_364),
.B2(n_357),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_424),
.A2(n_306),
.B1(n_348),
.B2(n_357),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_429),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_416),
.C(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_445),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_434),
.B(n_353),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_433),
.A2(n_348),
.B(n_423),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_L g453 ( 
.A1(n_446),
.A2(n_432),
.B(n_450),
.C(n_437),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_423),
.C(n_313),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_451),
.C(n_309),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_304),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_449),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_453),
.B(n_456),
.Y(n_459)
);

NAND4xp25_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_430),
.C(n_297),
.D(n_313),
.Y(n_454)
);

AOI322xp5_ASAP7_75t_L g462 ( 
.A1(n_454),
.A2(n_458),
.A3(n_241),
.B1(n_222),
.B2(n_10),
.C1(n_11),
.C2(n_13),
.Y(n_462)
);

AOI322xp5_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_309),
.A3(n_222),
.B1(n_241),
.B2(n_11),
.C1(n_7),
.C2(n_10),
.Y(n_458)
);

MAJx2_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_452),
.C(n_447),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g465 ( 
.A(n_460),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_457),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_461),
.B(n_458),
.C(n_222),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_462),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_463),
.A2(n_9),
.B1(n_13),
.B2(n_464),
.Y(n_467)
);

OAI221xp5_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_459),
.B1(n_9),
.B2(n_13),
.C(n_7),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_467),
.Y(n_468)
);


endmodule