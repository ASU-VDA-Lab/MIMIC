module fake_netlist_6_1810_n_72 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_72);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_72;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_21;
wire n_24;
wire n_18;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_19;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_40;
wire n_25;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx11_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

AND2x4_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_5),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_30),
.B(n_31),
.C(n_27),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_28),
.B(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_29),
.B(n_20),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_24),
.C(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OAI21x1_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_24),
.B(n_18),
.Y(n_43)
);

OA21x2_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_19),
.B(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_19),
.B(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_23),
.C(n_48),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

XOR2x2_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_48),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_57),
.B(n_50),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_51),
.B(n_43),
.C(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_60),
.B1(n_52),
.B2(n_43),
.Y(n_64)
);

OAI211xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_46),
.B(n_44),
.C(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_10),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

AOI22x1_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_25),
.B1(n_17),
.B2(n_44),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_69),
.Y(n_71)
);

OR2x6_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_69),
.Y(n_72)
);


endmodule