module fake_jpeg_29607_n_334 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_334);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_18),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_48),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_61),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_2),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_56),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_3),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_27),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_24),
.C(n_23),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_37),
.C(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_84),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_34),
.B1(n_22),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_81),
.B1(n_91),
.B2(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_34),
.B1(n_22),
.B2(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_82),
.B(n_100),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_41),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_87),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_96),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_34),
.B1(n_22),
.B2(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_31),
.B1(n_63),
.B2(n_55),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_31),
.B1(n_39),
.B2(n_29),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_57),
.B1(n_55),
.B2(n_51),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_59),
.B(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_99),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_19),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_30),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_30),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_39),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_113),
.A2(n_122),
.B1(n_131),
.B2(n_150),
.Y(n_178)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_20),
.B(n_38),
.C(n_35),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_138),
.Y(n_155)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_20),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_103),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_31),
.B(n_38),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_139),
.B(n_146),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_57),
.B1(n_51),
.B2(n_50),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_112),
.A2(n_34),
.B1(n_22),
.B2(n_35),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_128),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_50),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_130),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_39),
.B1(n_29),
.B2(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_140),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_103),
.B(n_76),
.C(n_72),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_24),
.B(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_39),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_102),
.Y(n_157)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_81),
.A2(n_29),
.B1(n_41),
.B2(n_5),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_91),
.A2(n_29),
.B(n_4),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_147),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_74),
.A2(n_3),
.B(n_4),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_97),
.B(n_111),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_153),
.B(n_163),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_143),
.B1(n_149),
.B2(n_147),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_141),
.B(n_71),
.Y(n_160)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_78),
.A3(n_70),
.B1(n_111),
.B2(n_79),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_176),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_95),
.B(n_107),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_164),
.A2(n_183),
.B(n_143),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_104),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_95),
.B(n_106),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_139),
.B(n_128),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_101),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_133),
.B(n_6),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_78),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_79),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_163),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_70),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_185),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_206),
.B(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_146),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_174),
.C(n_184),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_128),
.B1(n_143),
.B2(n_113),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_189),
.A2(n_209),
.B1(n_166),
.B2(n_156),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_192),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_135),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_207),
.B1(n_210),
.B2(n_191),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_204),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_143),
.B1(n_118),
.B2(n_114),
.Y(n_207)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_167),
.A2(n_114),
.A3(n_117),
.B1(n_116),
.B2(n_125),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_116),
.B1(n_144),
.B2(n_123),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_145),
.B1(n_142),
.B2(n_136),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_215),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_129),
.B(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_129),
.C(n_9),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_181),
.B1(n_174),
.B2(n_183),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_221),
.A2(n_200),
.B(n_180),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_157),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_231),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_172),
.B(n_155),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_224),
.A2(n_227),
.B(n_231),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_151),
.B1(n_173),
.B2(n_160),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_228),
.B1(n_229),
.B2(n_203),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_174),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_189),
.B1(n_213),
.B2(n_173),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_164),
.B1(n_162),
.B2(n_155),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_175),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_208),
.B1(n_209),
.B2(n_186),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_190),
.A2(n_179),
.B(n_182),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_240),
.B(n_206),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_153),
.B(n_152),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_201),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_193),
.B(n_171),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_205),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_194),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_250),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_233),
.B1(n_239),
.B2(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_257),
.B(n_261),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_252),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_236),
.B1(n_223),
.B2(n_218),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_215),
.C(n_156),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_264),
.C(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_259),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_8),
.Y(n_281)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_202),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_185),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_232),
.Y(n_272)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_263),
.B1(n_230),
.B2(n_233),
.Y(n_270)
);

OAI321xp33_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_170),
.A3(n_180),
.B1(n_161),
.B2(n_145),
.C(n_13),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_241),
.C(n_218),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.C(n_277),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_216),
.C(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

OAI322xp33_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_226),
.A3(n_222),
.B1(n_228),
.B2(n_240),
.C1(n_219),
.C2(n_221),
.Y(n_274)
);

OA21x2_ASAP7_75t_SL g290 ( 
.A1(n_274),
.A2(n_251),
.B(n_258),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_216),
.C(n_223),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_280),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_259),
.Y(n_288)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_290),
.B1(n_271),
.B2(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_257),
.C(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_264),
.C(n_261),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_258),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_246),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_244),
.C(n_252),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_300),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_275),
.B1(n_273),
.B2(n_279),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_301),
.B1(n_283),
.B2(n_263),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_276),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_273),
.B1(n_247),
.B2(n_245),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_278),
.B(n_262),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_288),
.B(n_287),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_17),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_282),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_309),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_282),
.C(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_305),
.C(n_301),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_286),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_312),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_255),
.B(n_281),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

OAI321xp33_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_306),
.A3(n_299),
.B1(n_13),
.B2(n_14),
.C(n_11),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_298),
.B(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_317),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_310),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_12),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_311),
.B(n_313),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_321),
.B(n_317),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_318),
.C(n_322),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

OAI311xp33_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.A3(n_15),
.B1(n_16),
.C1(n_330),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_318),
.C(n_327),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_15),
.Y(n_334)
);


endmodule