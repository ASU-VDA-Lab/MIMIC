module fake_jpeg_13262_n_180 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_33),
.Y(n_84)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_35),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_15),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_31),
.B(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_12),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

OR2x4_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_2),
.Y(n_62)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_56),
.B(n_50),
.Y(n_70)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_14),
.B1(n_38),
.B2(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_68),
.B1(n_74),
.B2(n_84),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_62),
.C(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_16),
.B1(n_53),
.B2(n_44),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_14),
.B(n_28),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_23),
.B(n_22),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_25),
.B1(n_16),
.B2(n_32),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g105 ( 
.A(n_70),
.B(n_71),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_33),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_33),
.B(n_26),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_34),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_25),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_93),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_101),
.B1(n_106),
.B2(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_6),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_96),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_6),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_98),
.C(n_78),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_4),
.C(n_5),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_4),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_4),
.B1(n_6),
.B2(n_60),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_103),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_88),
.B(n_91),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_128),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_84),
.A3(n_80),
.B1(n_73),
.B2(n_59),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_129),
.B(n_118),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_114),
.CON(n_142),
.SN(n_142)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_90),
.B(n_98),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_95),
.B(n_94),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_107),
.C(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_144),
.C(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_141),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_129),
.B1(n_119),
.B2(n_116),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_134),
.B(n_146),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_142),
.C(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_120),
.C(n_113),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_131),
.C(n_123),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_127),
.C(n_135),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_153),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_145),
.C(n_144),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_163),
.B1(n_143),
.B2(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_156),
.C(n_154),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_161),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_154),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_168),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_162),
.B1(n_159),
.B2(n_156),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_165),
.B(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_172),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_138),
.B1(n_139),
.B2(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_166),
.B(n_140),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_171),
.B(n_177),
.C(n_175),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_170),
.Y(n_180)
);


endmodule