module fake_netlist_6_4882_n_2142 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2142);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2142;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_56),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_151),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_69),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_130),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_80),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_37),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_7),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_126),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_32),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_160),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_100),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_80),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_154),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_7),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_82),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_206),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_23),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_88),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_157),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_123),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_12),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_106),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_202),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_70),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_199),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_51),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_171),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_169),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_141),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_60),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_57),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_125),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_163),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_78),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_190),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_120),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_78),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_111),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_197),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_65),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_182),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_178),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_21),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_51),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_115),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_31),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_35),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_217),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_91),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_207),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_196),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_90),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_53),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_63),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_134),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_221),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_92),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_2),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_113),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_39),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_133),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_35),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_48),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_166),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_128),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_97),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_74),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_155),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_59),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_83),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_153),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_55),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_50),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_77),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_187),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_95),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_10),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_42),
.Y(n_316)
);

BUFx8_ASAP7_75t_SL g317 ( 
.A(n_98),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_13),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_116),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_108),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_76),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_25),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_14),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_117),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_124),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_156),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_94),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_81),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_42),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_86),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_203),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_37),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_29),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_107),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_38),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_192),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_49),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_185),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_65),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_214),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_105),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_219),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_140),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_101),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_189),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_201),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_16),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_82),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_129),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_148),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_61),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_209),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_53),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_58),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_23),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_52),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_77),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_44),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_4),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_20),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_6),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_48),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_121),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_8),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_174),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_71),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_0),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_15),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_127),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_66),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_114),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_49),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_56),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_96),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_112),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_54),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_85),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_172),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_64),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_118),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_99),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_180),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_204),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_138),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_186),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_76),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_59),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_122),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_60),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_139),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_19),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_29),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_213),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_181),
.Y(n_398)
);

BUFx8_ASAP7_75t_SL g399 ( 
.A(n_143),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_179),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_194),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_150),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_170),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_152),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_61),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_46),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_142),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_83),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_70),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_64),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_66),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_84),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_68),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_18),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_33),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_12),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_183),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_41),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_191),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_131),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_198),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_87),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_40),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_167),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_57),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_45),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_13),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_32),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_188),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_144),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_119),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_75),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_20),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_44),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_102),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_215),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_146),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_223),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_241),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_241),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_241),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_241),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_241),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_241),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_241),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_244),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_244),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_296),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_244),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_244),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_244),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_317),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_310),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_310),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_399),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_275),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_310),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_310),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_310),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_420),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_276),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_306),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_365),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_223),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_303),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_236),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_230),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_236),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_388),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_295),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_295),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_227),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_341),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_341),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_283),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_358),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_230),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_261),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_368),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_368),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_363),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_232),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_284),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_377),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_289),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_248),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_232),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_257),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_271),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_312),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_332),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_333),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_336),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_363),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_290),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_343),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_314),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_355),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_357),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_238),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_359),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_360),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_320),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_266),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_364),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_323),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_371),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_326),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_327),
.Y(n_519)
);

INVxp33_ASAP7_75t_SL g520 ( 
.A(n_233),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_378),
.Y(n_521)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_233),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_376),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_329),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_334),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_406),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_363),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_234),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_234),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_261),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_427),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_340),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_288),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_288),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_346),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_266),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_259),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_347),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_261),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_321),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_321),
.Y(n_543)
);

INVxp33_ASAP7_75t_SL g544 ( 
.A(n_243),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_383),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_383),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_243),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_335),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_225),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_353),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_335),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_229),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_268),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_231),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_354),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_237),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_239),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_250),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_457),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_255),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_245),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_338),
.Y(n_563)
);

AND2x2_ASAP7_75t_R g564 ( 
.A(n_541),
.B(n_251),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_449),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_467),
.A2(n_318),
.B1(n_339),
.B2(n_278),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_439),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_501),
.B(n_254),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_439),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_440),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_447),
.Y(n_571)
);

NOR2x1_ASAP7_75t_L g572 ( 
.A(n_514),
.B(n_270),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_483),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_440),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_492),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_255),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_448),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_470),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_448),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_450),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_450),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_441),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_441),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_494),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_451),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_451),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_505),
.B(n_299),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_507),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_442),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_469),
.B(n_277),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_452),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_443),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_443),
.B(n_254),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_454),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_444),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_454),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_299),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_471),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_273),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_444),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_555),
.B(n_557),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_455),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_445),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_445),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_446),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_455),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_446),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_516),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_458),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_539),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_459),
.B(n_254),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_510),
.B(n_338),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_459),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_557),
.B(n_279),
.Y(n_618)
);

BUFx8_ASAP7_75t_L g619 ( 
.A(n_469),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_514),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_541),
.B(n_338),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_460),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_460),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_461),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_482),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_486),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_461),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_462),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_453),
.B(n_367),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_462),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_518),
.B(n_282),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_463),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_538),
.A2(n_286),
.B(n_285),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_554),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_463),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_535),
.B(n_302),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_466),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_466),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_525),
.B(n_291),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_514),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_474),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_519),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_534),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_474),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_484),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_484),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_475),
.A2(n_416),
.B1(n_253),
.B2(n_263),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_496),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_488),
.Y(n_651)
);

NOR2x1_ASAP7_75t_L g652 ( 
.A(n_538),
.B(n_294),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_488),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_540),
.B(n_300),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_600),
.B(n_556),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_568),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_643),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_560),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_571),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_568),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_643),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_634),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_568),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_567),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_643),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_567),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_643),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_614),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_573),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_571),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_569),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_563),
.B(n_501),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_620),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_563),
.B(n_545),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_569),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_614),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_561),
.B(n_464),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_575),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_570),
.Y(n_681)
);

OAI21xp33_ASAP7_75t_SL g682 ( 
.A1(n_621),
.A2(n_536),
.B(n_535),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_570),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_626),
.B(n_547),
.Y(n_684)
);

BUFx8_ASAP7_75t_SL g685 ( 
.A(n_565),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_570),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_643),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_590),
.B(n_558),
.Y(n_688)
);

CKINVDCx6p67_ASAP7_75t_R g689 ( 
.A(n_601),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_620),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_574),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_620),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_643),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_631),
.B(n_558),
.Y(n_694)
);

INVxp33_ASAP7_75t_L g695 ( 
.A(n_593),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_626),
.B(n_438),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_579),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_640),
.B(n_559),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_574),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_574),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_616),
.B(n_485),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_616),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_584),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_624),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_583),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_585),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_591),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_636),
.B(n_559),
.C(n_543),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_593),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_611),
.B(n_520),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_583),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_580),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_654),
.B(n_522),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_589),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_589),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_602),
.A2(n_490),
.B1(n_473),
.B2(n_529),
.Y(n_718)
);

AND3x2_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_264),
.C(n_489),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_589),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_592),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_592),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_645),
.B(n_544),
.Y(n_723)
);

AND2x6_ASAP7_75t_L g724 ( 
.A(n_584),
.B(n_254),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_561),
.B(n_542),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_592),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_644),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_584),
.B(n_603),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_584),
.B(n_542),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_595),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_629),
.B(n_524),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_595),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_625),
.B(n_537),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_619),
.Y(n_734)
);

AOI21x1_ASAP7_75t_L g735 ( 
.A1(n_595),
.A2(n_549),
.B(n_543),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_596),
.B(n_254),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_R g737 ( 
.A(n_636),
.B(n_473),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_602),
.B(n_552),
.C(n_549),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_603),
.B(n_552),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_602),
.A2(n_490),
.B1(n_530),
.B2(n_528),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_602),
.A2(n_478),
.B1(n_301),
.B2(n_421),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_603),
.B(n_486),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_598),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_603),
.B(n_607),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_607),
.B(n_531),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_649),
.B(n_551),
.Y(n_746)
);

AND2x2_ASAP7_75t_SL g747 ( 
.A(n_633),
.B(n_292),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_607),
.B(n_580),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_598),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_571),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_561),
.Y(n_751)
);

BUFx10_ASAP7_75t_L g752 ( 
.A(n_618),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_604),
.B(n_456),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_598),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_562),
.B(n_548),
.C(n_527),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_624),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_606),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_607),
.B(n_531),
.Y(n_758)
);

NOR2x1p5_ASAP7_75t_L g759 ( 
.A(n_561),
.B(n_245),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_606),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_618),
.B(n_497),
.C(n_495),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_606),
.Y(n_762)
);

OAI22x1_ASAP7_75t_L g763 ( 
.A1(n_566),
.A2(n_504),
.B1(n_546),
.B2(n_263),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_627),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_619),
.B(n_521),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_627),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_627),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_635),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_580),
.B(n_319),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_635),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_576),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_608),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_608),
.Y(n_773)
);

INVx6_ASAP7_75t_L g774 ( 
.A(n_620),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_576),
.B(n_503),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_608),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_610),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_597),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_610),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_576),
.Y(n_780)
);

AND3x1_ASAP7_75t_L g781 ( 
.A(n_566),
.B(n_536),
.C(n_497),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_610),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_597),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_635),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_641),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_599),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_641),
.Y(n_787)
);

CKINVDCx11_ASAP7_75t_R g788 ( 
.A(n_564),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_618),
.A2(n_414),
.B1(n_433),
.B2(n_423),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_571),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_652),
.A2(n_381),
.B1(n_280),
.B2(n_281),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_618),
.B(n_498),
.C(n_495),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_599),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_641),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_577),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_652),
.A2(n_313),
.B(n_308),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_571),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_599),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_619),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_633),
.B(n_499),
.C(n_498),
.Y(n_800)
);

AO21x2_ASAP7_75t_L g801 ( 
.A1(n_576),
.A2(n_330),
.B(n_328),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_571),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_604),
.B(n_379),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_577),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_604),
.B(n_503),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_578),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_604),
.B(n_224),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_578),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_582),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_581),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_581),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_582),
.B(n_392),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_586),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_715),
.B(n_619),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_656),
.A2(n_633),
.B1(n_596),
.B2(n_344),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_751),
.B(n_586),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_783),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_771),
.B(n_342),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_771),
.B(n_587),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_669),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_735),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_780),
.B(n_655),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_656),
.B(n_292),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_660),
.B(n_292),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_735),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_695),
.B(n_703),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_660),
.A2(n_633),
.B1(n_596),
.B2(n_348),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_783),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_663),
.B(n_292),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_780),
.B(n_588),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_747),
.A2(n_572),
.B(n_596),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_669),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_663),
.B(n_292),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_678),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_710),
.Y(n_836)
);

BUFx6f_ASAP7_75t_SL g837 ( 
.A(n_708),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_703),
.B(n_301),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_725),
.B(n_646),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_747),
.B(n_301),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_694),
.B(n_588),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_795),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_662),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_698),
.B(n_594),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_688),
.B(n_594),
.Y(n_845)
);

OAI22xp33_ASAP7_75t_L g846 ( 
.A1(n_803),
.A2(n_419),
.B1(n_349),
.B2(n_350),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_704),
.B(n_786),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_747),
.B(n_301),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_795),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_793),
.B(n_605),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_806),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_662),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_806),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_742),
.B(n_605),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_805),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_702),
.B(n_224),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_745),
.B(n_609),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_759),
.A2(n_373),
.B1(n_382),
.B2(n_369),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_758),
.B(n_609),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_804),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_752),
.B(n_301),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_804),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_710),
.B(n_499),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_805),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_659),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_725),
.B(n_646),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_679),
.B(n_808),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_808),
.B(n_809),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_697),
.B(n_675),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_809),
.B(n_623),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_775),
.B(n_647),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_759),
.A2(n_737),
.B1(n_673),
.B2(n_755),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_813),
.B(n_628),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_775),
.B(n_647),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_658),
.B(n_226),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_728),
.A2(n_744),
.B(n_748),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_714),
.B(n_628),
.Y(n_878)
);

OAI22xp33_ASAP7_75t_L g879 ( 
.A1(n_789),
.A2(n_356),
.B1(n_375),
.B2(n_345),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_676),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_727),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_685),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_724),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_723),
.B(n_226),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_714),
.B(n_630),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_778),
.B(n_630),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_778),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_778),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_752),
.B(n_421),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_670),
.B(n_648),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_791),
.A2(n_523),
.B(n_508),
.C(n_637),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_752),
.B(n_421),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_798),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_798),
.B(n_637),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_798),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_812),
.B(n_639),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_676),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_740),
.B(n_648),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_676),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_741),
.B(n_639),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_696),
.B(n_228),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_769),
.B(n_572),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_664),
.B(n_581),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_682),
.A2(n_385),
.B1(n_386),
.B2(n_384),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_684),
.B(n_228),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_733),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_682),
.B(n_235),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_781),
.A2(n_395),
.B1(n_274),
.B2(n_265),
.C(n_253),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_664),
.B(n_581),
.Y(n_909)
);

INVx4_ASAP7_75t_SL g910 ( 
.A(n_724),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_718),
.A2(n_397),
.B1(n_398),
.B2(n_387),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_664),
.B(n_700),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_664),
.B(n_581),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_700),
.B(n_581),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_708),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_801),
.A2(n_596),
.B1(n_431),
.B2(n_430),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_807),
.B(n_711),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_681),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_746),
.A2(n_389),
.B1(n_437),
.B2(n_235),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_784),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_801),
.A2(n_596),
.B1(n_404),
.B2(n_421),
.Y(n_921)
);

BUFx8_ASAP7_75t_L g922 ( 
.A(n_765),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_784),
.Y(n_923)
);

AOI221xp5_ASAP7_75t_L g924 ( 
.A1(n_781),
.A2(n_274),
.B1(n_265),
.B2(n_395),
.C(n_396),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_800),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_689),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_681),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_731),
.B(n_240),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_752),
.B(n_421),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_709),
.B(n_651),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_753),
.B(n_240),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_657),
.B(n_620),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_680),
.B(n_242),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_800),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_707),
.B(n_242),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_789),
.B(n_246),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_700),
.B(n_612),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_761),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_709),
.B(n_761),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_729),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_700),
.B(n_726),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_681),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_L g943 ( 
.A(n_734),
.B(n_396),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_L g944 ( 
.A(n_738),
.B(n_651),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_739),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_736),
.A2(n_508),
.B(n_523),
.C(n_502),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_738),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_792),
.A2(n_269),
.B1(n_246),
.B2(n_436),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_686),
.Y(n_949)
);

AND2x6_ASAP7_75t_SL g950 ( 
.A(n_788),
.B(n_500),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_792),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_763),
.B(n_500),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_666),
.A2(n_506),
.B(n_502),
.C(n_509),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_708),
.B(n_247),
.Y(n_954)
);

XNOR2xp5_ASAP7_75t_L g955 ( 
.A(n_763),
.B(n_405),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_708),
.Y(n_956)
);

AOI221xp5_ASAP7_75t_L g957 ( 
.A1(n_799),
.A2(n_413),
.B1(n_405),
.B2(n_409),
.C(n_410),
.Y(n_957)
);

AND2x4_ASAP7_75t_SL g958 ( 
.A(n_689),
.B(n_506),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_726),
.B(n_612),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_726),
.B(n_612),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_726),
.B(n_612),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_657),
.B(n_620),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_666),
.B(n_612),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_811),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_668),
.A2(n_596),
.B1(n_615),
.B2(n_642),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_719),
.B(n_247),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_686),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_661),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_668),
.B(n_612),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_661),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_672),
.A2(n_509),
.B(n_511),
.C(n_533),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_672),
.A2(n_260),
.B1(n_436),
.B2(n_429),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_699),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_659),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_699),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_677),
.B(n_613),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_665),
.A2(n_642),
.B(n_653),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_706),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_706),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_677),
.A2(n_526),
.B(n_511),
.C(n_533),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_829),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_855),
.B(n_512),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_833),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_833),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_829),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_860),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_823),
.A2(n_796),
.B1(n_691),
.B2(n_701),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_864),
.B(n_512),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_860),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_867),
.B(n_683),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_821),
.B(n_515),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_940),
.B(n_683),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_974),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_862),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_862),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_839),
.B(n_515),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_842),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_881),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_821),
.B(n_843),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_822),
.A2(n_811),
.B(n_667),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_835),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_816),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_842),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_852),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_849),
.Y(n_1005)
);

AO22x1_ASAP7_75t_L g1006 ( 
.A1(n_936),
.A2(n_410),
.B1(n_411),
.B2(n_409),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_917),
.A2(n_701),
.B1(n_712),
.B2(n_691),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_816),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_839),
.B(n_517),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_849),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_SL g1011 ( 
.A1(n_955),
.A2(n_413),
.B1(n_415),
.B2(n_411),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_851),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_851),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_945),
.B(n_712),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_906),
.B(n_713),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_866),
.B(n_517),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_816),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_853),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_827),
.B(n_526),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_845),
.B(n_713),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_882),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_925),
.B(n_934),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_866),
.B(n_532),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_826),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_SL g1025 ( 
.A(n_879),
.B(n_418),
.C(n_415),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_896),
.B(n_722),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_836),
.B(n_722),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_863),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_853),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_840),
.A2(n_732),
.B(n_730),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_816),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_871),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_951),
.B(n_732),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_939),
.B(n_249),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_841),
.B(n_743),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_832),
.B(n_797),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_872),
.B(n_797),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_844),
.B(n_743),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_907),
.A2(n_749),
.B(n_757),
.C(n_754),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_974),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_974),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_840),
.A2(n_848),
.B1(n_939),
.B2(n_947),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_876),
.B(n_749),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_938),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_863),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_871),
.B(n_754),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_848),
.A2(n_760),
.B1(n_762),
.B2(n_757),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_874),
.B(n_760),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_915),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_964),
.Y(n_1050)
);

INVx5_ASAP7_75t_L g1051 ( 
.A(n_883),
.Y(n_1051)
);

CKINVDCx11_ASAP7_75t_R g1052 ( 
.A(n_950),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_874),
.B(n_930),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_958),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_964),
.Y(n_1055)
);

AND3x2_ASAP7_75t_SL g1056 ( 
.A(n_955),
.B(n_425),
.C(n_418),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_930),
.B(n_762),
.Y(n_1057)
);

O2A1O1Ixp5_ASAP7_75t_L g1058 ( 
.A1(n_824),
.A2(n_796),
.B(n_772),
.C(n_720),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_974),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_884),
.B(n_773),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_974),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_818),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_L g1063 ( 
.A(n_954),
.B(n_532),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_915),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_826),
.B(n_706),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_880),
.Y(n_1066)
);

INVx5_ASAP7_75t_L g1067 ( 
.A(n_883),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_898),
.B(n_472),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_880),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_952),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_868),
.B(n_773),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_933),
.B(n_665),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_814),
.B(n_252),
.C(n_249),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_877),
.A2(n_779),
.B(n_777),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_869),
.B(n_779),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_952),
.B(n_425),
.Y(n_1076)
);

NAND3xp33_ASAP7_75t_SL g1077 ( 
.A(n_957),
.B(n_428),
.C(n_426),
.Y(n_1077)
);

BUFx8_ASAP7_75t_L g1078 ( 
.A(n_837),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_SL g1079 ( 
.A(n_837),
.B(n_815),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_897),
.Y(n_1080)
);

OR2x4_ASAP7_75t_L g1081 ( 
.A(n_966),
.B(n_472),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_SL g1082 ( 
.A(n_956),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_898),
.B(n_426),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_956),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_935),
.B(n_782),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_875),
.B(n_782),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_920),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_888),
.B(n_716),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_902),
.B(n_797),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_887),
.Y(n_1090)
);

O2A1O1Ixp5_ASAP7_75t_L g1091 ( 
.A1(n_824),
.A2(n_721),
.B(n_717),
.C(n_720),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_856),
.B(n_716),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_828),
.B(n_802),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_819),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_SL g1095 ( 
.A(n_908),
.B(n_434),
.C(n_428),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_920),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_847),
.B(n_716),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_893),
.B(n_802),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_895),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_819),
.B(n_802),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_928),
.B(n_717),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_883),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_923),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_890),
.B(n_811),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_901),
.B(n_476),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_819),
.B(n_667),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_943),
.B(n_687),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_899),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_899),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_905),
.B(n_717),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_926),
.B(n_434),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_865),
.B(n_790),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_865),
.B(n_687),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_924),
.A2(n_721),
.B1(n_720),
.B2(n_772),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_931),
.A2(n_790),
.B1(n_693),
.B2(n_776),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_854),
.B(n_721),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_865),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_918),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_857),
.B(n_859),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_817),
.B(n_772),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_919),
.B(n_476),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_972),
.B(n_825),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_927),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_883),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_870),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_927),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_911),
.B(n_293),
.C(n_287),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_968),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_SL g1129 ( 
.A(n_858),
.B(n_298),
.C(n_297),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_825),
.A2(n_776),
.B(n_693),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_820),
.B(n_790),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_830),
.B(n_304),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_922),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_822),
.B(n_790),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_L g1135 ( 
.A(n_830),
.B(n_784),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_922),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_822),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_942),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_831),
.B(n_705),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_942),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_949),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_949),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_904),
.A2(n_407),
.B1(n_256),
.B2(n_258),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_967),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_834),
.B(n_705),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_944),
.B(n_477),
.Y(n_1146)
);

NOR2x1p5_ASAP7_75t_L g1147 ( 
.A(n_922),
.B(n_305),
.Y(n_1147)
);

CKINVDCx6p67_ASAP7_75t_R g1148 ( 
.A(n_838),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_967),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_861),
.A2(n_671),
.B(n_659),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_834),
.B(n_873),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_838),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_978),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_878),
.B(n_756),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_921),
.A2(n_724),
.B1(n_794),
.B2(n_787),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_SL g1156 ( 
.A1(n_948),
.A2(n_307),
.B1(n_393),
.B2(n_390),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_861),
.A2(n_422),
.B1(n_256),
.B2(n_258),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_978),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_979),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1045),
.B(n_891),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1117),
.A2(n_892),
.B(n_889),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1053),
.B(n_968),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1042),
.A2(n_892),
.B(n_889),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1001),
.B(n_885),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_998),
.B(n_846),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1059),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_991),
.B(n_900),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_SL g1169 ( 
.A1(n_1022),
.A2(n_929),
.B(n_932),
.C(n_962),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1019),
.B(n_886),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_999),
.Y(n_1171)
);

BUFx12f_ASAP7_75t_L g1172 ( 
.A(n_1078),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1119),
.B(n_970),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1051),
.B(n_1067),
.Y(n_1174)
);

OAI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1095),
.A2(n_980),
.B1(n_971),
.B2(n_953),
.C(n_850),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1137),
.B(n_970),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1151),
.A2(n_929),
.B(n_912),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1122),
.A2(n_894),
.B(n_975),
.C(n_973),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1036),
.A2(n_941),
.B(n_909),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1004),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1073),
.B(n_311),
.C(n_309),
.Y(n_1181)
);

OAI22x1_ASAP7_75t_L g1182 ( 
.A1(n_1070),
.A2(n_374),
.B1(n_315),
.B2(n_316),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1011),
.A2(n_1021),
.B1(n_999),
.B2(n_1133),
.Y(n_1183)
);

BUFx4f_ASAP7_75t_SL g1184 ( 
.A(n_1078),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_1077),
.B(n_324),
.C(n_322),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1137),
.B(n_979),
.Y(n_1186)
);

O2A1O1Ixp5_ASAP7_75t_SL g1187 ( 
.A1(n_1037),
.A2(n_491),
.B(n_487),
.C(n_480),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_963),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1117),
.A2(n_913),
.B(n_903),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1057),
.A2(n_937),
.B(n_914),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1042),
.A2(n_916),
.B1(n_965),
.B2(n_959),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_R g1192 ( 
.A(n_1079),
.B(n_252),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_999),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_1039),
.A2(n_976),
.B(n_969),
.Y(n_1194)
);

BUFx4f_ASAP7_75t_L g1195 ( 
.A(n_1136),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1122),
.A2(n_961),
.B1(n_960),
.B2(n_932),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1125),
.B(n_962),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1060),
.A2(n_260),
.B1(n_262),
.B2(n_267),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1073),
.A2(n_946),
.B(n_977),
.C(n_794),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1129),
.A2(n_262),
.B1(n_267),
.B2(n_424),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1149),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1025),
.B(n_331),
.C(n_325),
.Y(n_1202)
);

INVx1_ASAP7_75t_SL g1203 ( 
.A(n_983),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1060),
.A2(n_269),
.B1(n_407),
.B2(n_417),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_985),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1052),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1085),
.A2(n_272),
.B1(n_422),
.B2(n_424),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1036),
.A2(n_671),
.B(n_659),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1125),
.B(n_337),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1026),
.B(n_756),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1059),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1052),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1094),
.A2(n_272),
.B1(n_417),
.B2(n_403),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1070),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1093),
.A2(n_671),
.B(n_810),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_R g1216 ( 
.A(n_1079),
.B(n_394),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1002),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1085),
.A2(n_401),
.B1(n_394),
.B2(n_400),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1093),
.A2(n_810),
.B(n_659),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_984),
.B(n_1063),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1075),
.A2(n_1092),
.B1(n_1110),
.B2(n_1101),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_986),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_984),
.B(n_400),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1037),
.A2(n_787),
.B(n_785),
.C(n_770),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1102),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1082),
.B(n_401),
.Y(n_1226)
);

CKINVDCx14_ASAP7_75t_R g1227 ( 
.A(n_1111),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1132),
.A2(n_785),
.B(n_770),
.C(n_768),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1044),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1132),
.A2(n_768),
.B(n_767),
.C(n_766),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1095),
.B(n_362),
.C(n_380),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1044),
.A2(n_767),
.B(n_766),
.C(n_764),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1032),
.B(n_764),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1075),
.B(n_659),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1092),
.A2(n_1086),
.B(n_1034),
.C(n_1110),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1028),
.B(n_477),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1101),
.A2(n_810),
.B(n_671),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1054),
.A2(n_351),
.B1(n_352),
.B2(n_361),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1034),
.A2(n_402),
.B1(n_429),
.B2(n_403),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1059),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1020),
.B(n_671),
.Y(n_1241)
);

BUFx4_ASAP7_75t_SL g1242 ( 
.A(n_1049),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_993),
.A2(n_671),
.B(n_810),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_996),
.B(n_910),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1083),
.A2(n_653),
.B(n_481),
.C(n_487),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_996),
.B(n_910),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1155),
.A2(n_493),
.B(n_491),
.Y(n_1247)
);

NOR2x1_ASAP7_75t_R g1248 ( 
.A(n_1049),
.B(n_1064),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1009),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_990),
.A2(n_810),
.B(n_750),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1035),
.B(n_750),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1080),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1155),
.A2(n_1015),
.B(n_1152),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1039),
.A2(n_642),
.B(n_481),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1118),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1000),
.A2(n_479),
.B(n_480),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_993),
.A2(n_750),
.B1(n_810),
.B2(n_370),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1015),
.A2(n_1121),
.B(n_1086),
.C(n_1076),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1081),
.Y(n_1259)
);

BUFx4f_ASAP7_75t_SL g1260 ( 
.A(n_1081),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1038),
.B(n_750),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1027),
.B(n_366),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1071),
.A2(n_750),
.B(n_674),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1027),
.B(n_372),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_989),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1009),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1064),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1118),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1062),
.A2(n_493),
.B(n_479),
.C(n_2),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1016),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1046),
.A2(n_674),
.B(n_690),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_994),
.Y(n_1272)
);

AO32x1_ASAP7_75t_L g1273 ( 
.A1(n_987),
.A2(n_724),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1048),
.A2(n_674),
.B(n_690),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1016),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1143),
.A2(n_638),
.B(n_632),
.C(n_622),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1023),
.B(n_910),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1074),
.A2(n_690),
.B(n_692),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_995),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1134),
.A2(n_690),
.B(n_692),
.Y(n_1280)
);

INVx5_ASAP7_75t_L g1281 ( 
.A(n_1102),
.Y(n_1281)
);

NOR3xp33_ASAP7_75t_SL g1282 ( 
.A(n_1156),
.B(n_0),
.C(n_1),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1102),
.Y(n_1283)
);

BUFx4f_ASAP7_75t_L g1284 ( 
.A(n_1148),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1087),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1105),
.B(n_3),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1134),
.A2(n_692),
.B(n_910),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1158),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1023),
.B(n_5),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1097),
.A2(n_692),
.B(n_613),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_R g1291 ( 
.A(n_1082),
.B(n_89),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1090),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1068),
.B(n_982),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1107),
.A2(n_1104),
.B1(n_988),
.B2(n_982),
.Y(n_1294)
);

INVx5_ASAP7_75t_L g1295 ( 
.A(n_1102),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1107),
.B(n_93),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1090),
.B(n_5),
.Y(n_1297)
);

OR2x6_ASAP7_75t_L g1298 ( 
.A(n_1084),
.B(n_774),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1096),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1099),
.B(n_6),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1099),
.B(n_8),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_992),
.A2(n_774),
.B1(n_638),
.B2(n_632),
.Y(n_1302)
);

NOR3xp33_ASAP7_75t_SL g1303 ( 
.A(n_1127),
.B(n_9),
.C(n_10),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_988),
.B(n_9),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1104),
.B(n_613),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1089),
.A2(n_622),
.B(n_617),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1084),
.B(n_1124),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1103),
.Y(n_1308)
);

CKINVDCx8_ASAP7_75t_R g1309 ( 
.A(n_1146),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1089),
.A2(n_622),
.B(n_617),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1146),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1128),
.B(n_613),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1006),
.B(n_11),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1050),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1158),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1170),
.B(n_1014),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1221),
.B(n_1116),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1164),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1258),
.A2(n_1072),
.B(n_1043),
.C(n_1007),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1168),
.B(n_1033),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1293),
.B(n_1147),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1262),
.B(n_1264),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1173),
.A2(n_1050),
.B1(n_1055),
.B2(n_1128),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1208),
.A2(n_1091),
.B(n_1058),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1205),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1177),
.A2(n_1030),
.B(n_1130),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1167),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1281),
.B(n_1040),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1215),
.A2(n_1150),
.B(n_1098),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1285),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1309),
.B(n_1128),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1286),
.A2(n_1100),
.B(n_1139),
.C(n_1115),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1266),
.B(n_1157),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1181),
.A2(n_1055),
.B1(n_1100),
.B2(n_1106),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1289),
.A2(n_1106),
.B1(n_1018),
.B2(n_997),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1229),
.B(n_1012),
.Y(n_1336)
);

NOR4xp25_ASAP7_75t_L g1337 ( 
.A(n_1269),
.B(n_1313),
.C(n_1253),
.D(n_1202),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1180),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1160),
.B(n_1024),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1163),
.A2(n_1113),
.B(n_1131),
.Y(n_1340)
);

OA21x2_ASAP7_75t_L g1341 ( 
.A1(n_1237),
.A2(n_1154),
.B(n_1120),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1161),
.A2(n_1067),
.B(n_1051),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1225),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1189),
.A2(n_1088),
.B(n_1135),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1234),
.A2(n_1051),
.B(n_1067),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1214),
.B(n_1013),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1209),
.B(n_1024),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1276),
.A2(n_1145),
.A3(n_1029),
.B(n_1005),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_SL g1349 ( 
.A(n_1284),
.B(n_1124),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1167),
.Y(n_1350)
);

OAI22x1_ASAP7_75t_L g1351 ( 
.A1(n_1294),
.A2(n_1056),
.B1(n_1010),
.B2(n_1003),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1177),
.A2(n_1114),
.B(n_1047),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1306),
.A2(n_1112),
.B(n_1153),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1183),
.A2(n_1056),
.B1(n_1114),
.B2(n_1047),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1162),
.B(n_1066),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1236),
.B(n_1069),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1197),
.B(n_1138),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1179),
.A2(n_1190),
.B(n_1196),
.Y(n_1358)
);

INVx5_ASAP7_75t_L g1359 ( 
.A(n_1167),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1179),
.A2(n_1140),
.B(n_1144),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1197),
.B(n_1141),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1237),
.A2(n_1061),
.B(n_1041),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1165),
.B(n_1249),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1200),
.B(n_1123),
.C(n_1108),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1281),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1178),
.A2(n_1109),
.A3(n_1126),
.B(n_1159),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1242),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1270),
.B(n_1142),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1275),
.B(n_1008),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1299),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1311),
.B(n_1008),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1241),
.A2(n_1124),
.B(n_1031),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1267),
.B(n_1017),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1187),
.A2(n_1065),
.B(n_1031),
.Y(n_1374)
);

NAND3xp33_ASAP7_75t_L g1375 ( 
.A(n_1303),
.B(n_1017),
.C(n_638),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1250),
.A2(n_1224),
.B(n_1191),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1281),
.Y(n_1377)
);

CKINVDCx6p67_ASAP7_75t_R g1378 ( 
.A(n_1172),
.Y(n_1378)
);

AO31x2_ASAP7_75t_L g1379 ( 
.A1(n_1250),
.A2(n_1065),
.A3(n_724),
.B(n_615),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1225),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1282),
.B(n_638),
.C(n_632),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1166),
.B(n_613),
.Y(n_1382)
);

O2A1O1Ixp5_ASAP7_75t_L g1383 ( 
.A1(n_1220),
.A2(n_1065),
.B(n_724),
.C(n_15),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1228),
.A2(n_1065),
.B(n_724),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1310),
.A2(n_173),
.B(n_104),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1283),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_R g1387 ( 
.A(n_1227),
.B(n_103),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1310),
.A2(n_175),
.B(n_110),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_SL g1389 ( 
.A(n_1171),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1188),
.A2(n_1261),
.A3(n_1251),
.B(n_1278),
.Y(n_1390)
);

NOR2x1_ASAP7_75t_SL g1391 ( 
.A(n_1281),
.B(n_617),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1185),
.A2(n_632),
.B(n_622),
.C(n_617),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1278),
.A2(n_622),
.B(n_617),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1304),
.B(n_11),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1199),
.A2(n_1175),
.B(n_1297),
.C(n_1300),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_SL g1396 ( 
.A1(n_1188),
.A2(n_222),
.B(n_218),
.Y(n_1396)
);

AOI31xp67_ASAP7_75t_L g1397 ( 
.A1(n_1175),
.A2(n_615),
.A3(n_617),
.B(n_212),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1243),
.A2(n_161),
.B(n_132),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1176),
.Y(n_1399)
);

AOI221x1_ASAP7_75t_L g1400 ( 
.A1(n_1182),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_1400)
);

AO22x2_ASAP7_75t_L g1401 ( 
.A1(n_1231),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_1401)
);

INVx8_ASAP7_75t_L g1402 ( 
.A(n_1307),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1211),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1174),
.A2(n_168),
.B(n_135),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1203),
.B(n_22),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1292),
.B(n_24),
.Y(n_1406)
);

CKINVDCx6p67_ASAP7_75t_R g1407 ( 
.A(n_1212),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1283),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1307),
.Y(n_1409)
);

AOI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1290),
.A2(n_615),
.B(n_211),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1308),
.B(n_26),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1290),
.A2(n_149),
.B(n_195),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1176),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1210),
.B(n_28),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1314),
.B(n_30),
.Y(n_1415)
);

BUFx10_ASAP7_75t_L g1416 ( 
.A(n_1301),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1302),
.A2(n_615),
.A3(n_33),
.B(n_34),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1256),
.A2(n_177),
.B(n_159),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1263),
.A2(n_145),
.B(n_137),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1222),
.B(n_30),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1169),
.A2(n_109),
.B(n_615),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1259),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1186),
.A2(n_615),
.B(n_36),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1307),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1265),
.B(n_40),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1193),
.B(n_1296),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1272),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1207),
.B(n_41),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1245),
.A2(n_43),
.B(n_45),
.C(n_47),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1230),
.A2(n_43),
.B(n_47),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1271),
.A2(n_50),
.B(n_54),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1186),
.A2(n_55),
.B(n_62),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1271),
.A2(n_62),
.B(n_63),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1274),
.A2(n_67),
.B(n_68),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1218),
.B(n_67),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1238),
.B(n_69),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1279),
.B(n_86),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_SL g1438 ( 
.A1(n_1244),
.A2(n_71),
.B(n_72),
.C(n_73),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1296),
.B(n_72),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1257),
.A2(n_75),
.A3(n_79),
.B(n_81),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1233),
.B(n_1204),
.Y(n_1441)
);

OAI22x1_ASAP7_75t_L g1442 ( 
.A1(n_1239),
.A2(n_85),
.B1(n_79),
.B2(n_84),
.Y(n_1442)
);

BUFx10_ASAP7_75t_L g1443 ( 
.A(n_1298),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1298),
.B(n_1246),
.Y(n_1444)
);

AO21x1_ASAP7_75t_L g1445 ( 
.A1(n_1312),
.A2(n_1232),
.B(n_1305),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1254),
.A2(n_1274),
.B(n_1247),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1194),
.A2(n_1287),
.B(n_1280),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1254),
.A2(n_1233),
.B(n_1315),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1252),
.A2(n_1288),
.B(n_1268),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1198),
.B(n_1255),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1277),
.A2(n_1201),
.B(n_1223),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1194),
.A2(n_1295),
.B(n_1217),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1217),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1195),
.Y(n_1454)
);

AND2x6_ASAP7_75t_L g1455 ( 
.A(n_1211),
.B(n_1240),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_L g1456 ( 
.A(n_1295),
.B(n_1216),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1273),
.A2(n_1192),
.A3(n_1211),
.B(n_1240),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1240),
.A2(n_1273),
.B1(n_1260),
.B2(n_1213),
.C(n_1284),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1248),
.B(n_1226),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1295),
.B(n_1195),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1295),
.A2(n_1291),
.B(n_1184),
.C(n_1206),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1235),
.A2(n_1177),
.B(n_1039),
.Y(n_1462)
);

CKINVDCx6p67_ASAP7_75t_R g1463 ( 
.A(n_1172),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1170),
.B(n_1221),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1225),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1164),
.Y(n_1466)
);

CKINVDCx6p67_ASAP7_75t_R g1467 ( 
.A(n_1172),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1180),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1221),
.A2(n_1235),
.B1(n_1053),
.B2(n_1042),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1164),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1208),
.A2(n_1219),
.B(n_1215),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1170),
.B(n_1221),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1293),
.B(n_669),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1242),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1281),
.B(n_1295),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1214),
.B(n_669),
.Y(n_1476)
);

AO31x2_ASAP7_75t_L g1477 ( 
.A1(n_1276),
.A2(n_1039),
.A3(n_1235),
.B(n_1221),
.Y(n_1477)
);

AO21x1_ASAP7_75t_L g1478 ( 
.A1(n_1221),
.A2(n_1163),
.B(n_1122),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1366),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1322),
.A2(n_1395),
.B1(n_1476),
.B2(n_1354),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1329),
.A2(n_1344),
.B(n_1446),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1446),
.A2(n_1342),
.B(n_1353),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1318),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1325),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1428),
.A2(n_1435),
.B1(n_1436),
.B2(n_1337),
.C(n_1469),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1358),
.A2(n_1462),
.B(n_1376),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1478),
.A2(n_1354),
.B1(n_1442),
.B2(n_1401),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1330),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1473),
.B(n_1316),
.Y(n_1490)
);

INVx3_ASAP7_75t_SL g1491 ( 
.A(n_1367),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1320),
.B(n_1464),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1358),
.A2(n_1462),
.B(n_1376),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1333),
.B(n_1426),
.Y(n_1494)
);

AOI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1345),
.A2(n_1452),
.B(n_1410),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1346),
.B(n_1368),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1366),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1472),
.B(n_1382),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1324),
.A2(n_1419),
.B(n_1362),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1360),
.A2(n_1412),
.B(n_1421),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1399),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1366),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1360),
.A2(n_1418),
.B(n_1398),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1402),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1401),
.A2(n_1413),
.B1(n_1430),
.B2(n_1469),
.Y(n_1505)
);

AOI222xp33_ASAP7_75t_L g1506 ( 
.A1(n_1413),
.A2(n_1430),
.B1(n_1424),
.B2(n_1405),
.C1(n_1394),
.C2(n_1439),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1370),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1338),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1347),
.B(n_1339),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1431),
.A2(n_1385),
.B(n_1372),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1466),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1365),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1444),
.B(n_1373),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1432),
.A2(n_1352),
.B1(n_1416),
.B2(n_1317),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1336),
.Y(n_1515)
);

OAI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1319),
.A2(n_1332),
.B(n_1337),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1402),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1407),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1369),
.B(n_1441),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1409),
.A2(n_1389),
.B1(n_1363),
.B2(n_1334),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1470),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1326),
.A2(n_1458),
.B(n_1374),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1392),
.A2(n_1414),
.B(n_1364),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1384),
.A2(n_1433),
.B(n_1434),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1409),
.A2(n_1460),
.B1(n_1335),
.B2(n_1331),
.Y(n_1525)
);

CKINVDCx6p67_ASAP7_75t_R g1526 ( 
.A(n_1378),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1429),
.A2(n_1438),
.B1(n_1406),
.B2(n_1411),
.C(n_1425),
.Y(n_1527)
);

CKINVDCx14_ASAP7_75t_R g1528 ( 
.A(n_1463),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1335),
.A2(n_1454),
.B1(n_1356),
.B2(n_1450),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1427),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1387),
.A2(n_1402),
.B1(n_1349),
.B2(n_1381),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1381),
.A2(n_1437),
.B1(n_1420),
.B2(n_1375),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1357),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1474),
.B(n_1349),
.Y(n_1534)
);

OAI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1400),
.A2(n_1415),
.B1(n_1375),
.B2(n_1361),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1341),
.A2(n_1384),
.B(n_1451),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1371),
.B(n_1422),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1468),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1341),
.A2(n_1449),
.B(n_1396),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1444),
.B(n_1373),
.Y(n_1540)
);

INVx6_ASAP7_75t_L g1541 ( 
.A(n_1468),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1355),
.Y(n_1542)
);

AOI222xp33_ASAP7_75t_L g1543 ( 
.A1(n_1321),
.A2(n_1459),
.B1(n_1364),
.B2(n_1456),
.C1(n_1461),
.C2(n_1449),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_SL g1544 ( 
.A(n_1467),
.B(n_1377),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1458),
.A2(n_1423),
.B(n_1445),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1453),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1327),
.B(n_1403),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1365),
.B(n_1377),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1323),
.A2(n_1465),
.B1(n_1408),
.B2(n_1386),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1440),
.Y(n_1550)
);

NOR3xp33_ASAP7_75t_SL g1551 ( 
.A(n_1443),
.B(n_1440),
.C(n_1404),
.Y(n_1551)
);

NOR2xp67_ASAP7_75t_L g1552 ( 
.A(n_1343),
.B(n_1408),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1440),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1383),
.A2(n_1477),
.B(n_1465),
.C(n_1343),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1475),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1380),
.B(n_1386),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1328),
.A2(n_1475),
.B(n_1380),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1390),
.Y(n_1558)
);

INVx6_ASAP7_75t_L g1559 ( 
.A(n_1359),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1359),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1328),
.A2(n_1397),
.B(n_1348),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1350),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1348),
.A2(n_1477),
.B(n_1390),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1348),
.A2(n_1390),
.B(n_1477),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1359),
.A2(n_1457),
.B(n_1388),
.C(n_1403),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1350),
.A2(n_1443),
.B1(n_1457),
.B2(n_1417),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1417),
.B(n_1457),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_SL g1568 ( 
.A1(n_1391),
.A2(n_1417),
.B(n_1388),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1340),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1340),
.B(n_1455),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1455),
.Y(n_1571)
);

OAI211xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1379),
.A2(n_1322),
.B(n_872),
.C(n_1282),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1455),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1455),
.B(n_1322),
.Y(n_1574)
);

A2O1A1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1322),
.A2(n_1286),
.B(n_1235),
.C(n_1258),
.Y(n_1575)
);

AOI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1322),
.A2(n_936),
.B1(n_879),
.B2(n_814),
.C(n_1006),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1318),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1358),
.A2(n_1221),
.B(n_1322),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1322),
.B(n_449),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1358),
.A2(n_1221),
.B(n_1322),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1367),
.Y(n_1581)
);

NOR2xp67_ASAP7_75t_L g1582 ( 
.A(n_1476),
.B(n_678),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1322),
.A2(n_814),
.B1(n_1395),
.B2(n_884),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1322),
.B(n_1473),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1402),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1322),
.A2(n_884),
.B(n_1395),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1322),
.A2(n_884),
.B(n_1395),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1318),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1359),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1322),
.B(n_1473),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1318),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1468),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1365),
.B(n_1377),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1322),
.A2(n_884),
.B(n_1395),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1448),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1318),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1448),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1318),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1318),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1448),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1322),
.A2(n_884),
.B(n_1395),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1358),
.A2(n_1462),
.B(n_1376),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1358),
.A2(n_1376),
.B(n_1446),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1365),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1322),
.B(n_449),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1468),
.Y(n_1607)
);

AO31x2_ASAP7_75t_L g1608 ( 
.A1(n_1478),
.A2(n_1447),
.A3(n_1469),
.B(n_1039),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1318),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1402),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1473),
.B(n_1293),
.Y(n_1611)
);

BUFx4f_ASAP7_75t_L g1612 ( 
.A(n_1468),
.Y(n_1612)
);

AO31x2_ASAP7_75t_L g1613 ( 
.A1(n_1478),
.A2(n_1447),
.A3(n_1469),
.B(n_1039),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1322),
.A2(n_814),
.B1(n_715),
.B2(n_621),
.C(n_1166),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1616)
);

OAI22x1_ASAP7_75t_L g1617 ( 
.A1(n_1322),
.A2(n_1435),
.B1(n_1428),
.B2(n_814),
.Y(n_1617)
);

NOR2xp67_ASAP7_75t_L g1618 ( 
.A(n_1476),
.B(n_678),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1448),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1358),
.A2(n_1376),
.B(n_1446),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1318),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_SL g1623 ( 
.A(n_1367),
.B(n_669),
.Y(n_1623)
);

NAND2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1365),
.B(n_1377),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1473),
.B(n_1293),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1322),
.B(n_1473),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1468),
.Y(n_1627)
);

INVx6_ASAP7_75t_L g1628 ( 
.A(n_1468),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1448),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1318),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1318),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1468),
.Y(n_1634)
);

AOI22x1_ASAP7_75t_L g1635 ( 
.A1(n_1351),
.A2(n_1430),
.B1(n_1434),
.B2(n_1433),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1473),
.B(n_1293),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1318),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1448),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1358),
.A2(n_1462),
.B(n_1376),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1322),
.B(n_449),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1365),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1393),
.A2(n_1447),
.B(n_1471),
.Y(n_1643)
);

AO32x2_ASAP7_75t_L g1644 ( 
.A1(n_1469),
.A2(n_1413),
.A3(n_1354),
.B1(n_1221),
.B2(n_911),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1338),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1513),
.B(n_1540),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1583),
.A2(n_1615),
.B(n_1587),
.C(n_1595),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1501),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1576),
.A2(n_1486),
.B(n_1602),
.C(n_1586),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_SL g1651 ( 
.A1(n_1567),
.A2(n_1574),
.B(n_1509),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1508),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1494),
.B(n_1611),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1625),
.B(n_1636),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_R g1655 ( 
.A(n_1612),
.B(n_1534),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1490),
.B(n_1519),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1519),
.B(n_1584),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1607),
.B(n_1627),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1591),
.B(n_1626),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1612),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1578),
.A2(n_1580),
.B(n_1493),
.Y(n_1661)
);

AOI21x1_ASAP7_75t_SL g1662 ( 
.A1(n_1556),
.A2(n_1540),
.B(n_1513),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1575),
.A2(n_1481),
.B(n_1505),
.C(n_1527),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1484),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1487),
.A2(n_1603),
.B(n_1493),
.Y(n_1665)
);

O2A1O1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1572),
.A2(n_1506),
.B(n_1523),
.C(n_1535),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1557),
.B(n_1590),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1496),
.B(n_1542),
.Y(n_1668)
);

AOI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1579),
.A2(n_1606),
.B(n_1640),
.C(n_1520),
.Y(n_1669)
);

BUFx2_ASAP7_75t_SL g1670 ( 
.A(n_1538),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1537),
.B(n_1488),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1617),
.A2(n_1505),
.B1(n_1488),
.B2(n_1514),
.C(n_1535),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1561),
.A2(n_1500),
.B(n_1536),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1529),
.A2(n_1560),
.B(n_1554),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1531),
.A2(n_1582),
.B1(n_1618),
.B2(n_1640),
.Y(n_1675)
);

AOI221x1_ASAP7_75t_SL g1676 ( 
.A1(n_1498),
.A2(n_1606),
.B1(n_1579),
.B2(n_1550),
.C(n_1553),
.Y(n_1676)
);

O2A1O1Ixp5_ASAP7_75t_L g1677 ( 
.A1(n_1563),
.A2(n_1566),
.B(n_1495),
.C(n_1570),
.Y(n_1677)
);

AOI21x1_ASAP7_75t_SL g1678 ( 
.A1(n_1556),
.A2(n_1635),
.B(n_1644),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1485),
.B(n_1489),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1525),
.A2(n_1554),
.B(n_1549),
.C(n_1543),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1507),
.B(n_1511),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1645),
.B(n_1533),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1521),
.B(n_1530),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1480),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1538),
.Y(n_1685)
);

O2A1O1Ixp5_ASAP7_75t_L g1686 ( 
.A1(n_1566),
.A2(n_1570),
.B(n_1558),
.C(n_1565),
.Y(n_1686)
);

NOR2xp67_ASAP7_75t_L g1687 ( 
.A(n_1589),
.B(n_1593),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1639),
.A2(n_1620),
.B(n_1604),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1577),
.B(n_1588),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1592),
.B(n_1597),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1599),
.B(n_1600),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1549),
.A2(n_1532),
.B(n_1609),
.C(n_1621),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1631),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1632),
.B(n_1637),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1571),
.A2(n_1569),
.B1(n_1541),
.B2(n_1628),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1546),
.B(n_1639),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1562),
.B(n_1504),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1497),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1504),
.B(n_1517),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1551),
.A2(n_1568),
.B(n_1524),
.C(n_1623),
.Y(n_1700)
);

AOI21x1_ASAP7_75t_SL g1701 ( 
.A1(n_1556),
.A2(n_1644),
.B(n_1524),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1589),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1571),
.A2(n_1569),
.B1(n_1541),
.B2(n_1628),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1545),
.A2(n_1544),
.B(n_1573),
.C(n_1502),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1541),
.A2(n_1628),
.B1(n_1585),
.B2(n_1504),
.Y(n_1705)
);

AOI21x1_ASAP7_75t_SL g1706 ( 
.A1(n_1644),
.A2(n_1545),
.B(n_1613),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1547),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1517),
.B(n_1610),
.Y(n_1708)
);

NOR2xp67_ASAP7_75t_L g1709 ( 
.A(n_1593),
.B(n_1634),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1610),
.B(n_1644),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1608),
.B(n_1613),
.Y(n_1711)
);

O2A1O1Ixp5_ASAP7_75t_L g1712 ( 
.A1(n_1596),
.A2(n_1619),
.B(n_1598),
.C(n_1629),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1601),
.A2(n_1638),
.B(n_1629),
.C(n_1555),
.Y(n_1713)
);

O2A1O1Ixp5_ASAP7_75t_L g1714 ( 
.A1(n_1601),
.A2(n_1555),
.B(n_1512),
.C(n_1642),
.Y(n_1714)
);

AOI21x1_ASAP7_75t_SL g1715 ( 
.A1(n_1608),
.A2(n_1613),
.B(n_1522),
.Y(n_1715)
);

O2A1O1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1528),
.A2(n_1548),
.B(n_1624),
.C(n_1594),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1608),
.B(n_1610),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1559),
.A2(n_1528),
.B1(n_1552),
.B2(n_1518),
.Y(n_1718)
);

OR2x2_ASAP7_75t_SL g1719 ( 
.A(n_1559),
.B(n_1560),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1564),
.B(n_1539),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1491),
.B(n_1581),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1491),
.A2(n_1539),
.B(n_1503),
.C(n_1581),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1560),
.A2(n_1590),
.B(n_1624),
.Y(n_1723)
);

O2A1O1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1548),
.A2(n_1594),
.B(n_1605),
.C(n_1642),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1479),
.A2(n_1643),
.B(n_1641),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1526),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1560),
.B(n_1590),
.Y(n_1727)
);

O2A1O1Ixp5_ASAP7_75t_L g1728 ( 
.A1(n_1483),
.A2(n_1510),
.B(n_1482),
.C(n_1499),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1518),
.Y(n_1729)
);

AOI21x1_ASAP7_75t_SL g1730 ( 
.A1(n_1614),
.A2(n_1616),
.B(n_1622),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1616),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1630),
.A2(n_1322),
.B(n_1583),
.C(n_1615),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1633),
.A2(n_1221),
.B(n_1586),
.Y(n_1733)
);

AOI221x1_ASAP7_75t_SL g1734 ( 
.A1(n_1481),
.A2(n_879),
.B1(n_936),
.B2(n_1322),
.C(n_1583),
.Y(n_1734)
);

CKINVDCx6p67_ASAP7_75t_R g1735 ( 
.A(n_1491),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1496),
.B(n_1490),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1615),
.A2(n_1322),
.B1(n_1486),
.B2(n_1576),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1615),
.A2(n_1322),
.B1(n_1486),
.B2(n_1576),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1496),
.B(n_1490),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1494),
.B(n_1611),
.Y(n_1741)
);

O2A1O1Ixp5_ASAP7_75t_L g1742 ( 
.A1(n_1583),
.A2(n_1516),
.B(n_1587),
.C(n_1586),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1583),
.A2(n_1322),
.B(n_1615),
.C(n_1587),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_SL g1744 ( 
.A1(n_1567),
.A2(n_1322),
.B(n_1574),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1586),
.A2(n_837),
.B(n_1587),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1583),
.A2(n_1322),
.B(n_1615),
.C(n_1587),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1516),
.A2(n_1561),
.B(n_1500),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1586),
.A2(n_837),
.B(n_1587),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1515),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1579),
.B(n_727),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1494),
.B(n_1611),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1586),
.A2(n_837),
.B(n_1587),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1615),
.A2(n_1322),
.B1(n_1486),
.B2(n_1576),
.Y(n_1756)
);

O2A1O1Ixp5_ASAP7_75t_L g1757 ( 
.A1(n_1583),
.A2(n_1516),
.B(n_1587),
.C(n_1586),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1586),
.A2(n_1221),
.B(n_1587),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1504),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1494),
.B(n_1611),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1516),
.A2(n_1561),
.B(n_1500),
.Y(n_1762)
);

AOI21x1_ASAP7_75t_SL g1763 ( 
.A1(n_1567),
.A2(n_1322),
.B(n_1574),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1494),
.B(n_1611),
.Y(n_1765)
);

AOI21x1_ASAP7_75t_SL g1766 ( 
.A1(n_1567),
.A2(n_1322),
.B(n_1574),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1496),
.B(n_1490),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1586),
.A2(n_1221),
.B(n_1587),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1496),
.B(n_1490),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1513),
.B(n_1540),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1494),
.B(n_1611),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1667),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1696),
.B(n_1711),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1649),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1646),
.B(n_1736),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1752),
.B(n_1657),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1746),
.B(n_1749),
.Y(n_1778)
);

BUFx12f_ASAP7_75t_L g1779 ( 
.A(n_1726),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1717),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1710),
.B(n_1671),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1684),
.Y(n_1782)
);

AO21x2_ASAP7_75t_L g1783 ( 
.A1(n_1688),
.A2(n_1768),
.B(n_1758),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1664),
.B(n_1693),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1652),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1677),
.A2(n_1686),
.B(n_1742),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1674),
.B(n_1745),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1663),
.A2(n_1650),
.B(n_1648),
.Y(n_1788)
);

CKINVDCx6p67_ASAP7_75t_R g1789 ( 
.A(n_1735),
.Y(n_1789)
);

AO21x2_ASAP7_75t_L g1790 ( 
.A1(n_1733),
.A2(n_1661),
.B(n_1665),
.Y(n_1790)
);

OA21x2_ASAP7_75t_L g1791 ( 
.A1(n_1677),
.A2(n_1686),
.B(n_1742),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1698),
.Y(n_1792)
);

INVx4_ASAP7_75t_L g1793 ( 
.A(n_1667),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1712),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1719),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1751),
.Y(n_1796)
);

CKINVDCx6p67_ASAP7_75t_R g1797 ( 
.A(n_1660),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1751),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1689),
.B(n_1691),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1743),
.A2(n_1747),
.B(n_1648),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1738),
.A2(n_1739),
.B(n_1756),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1679),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1681),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1682),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1683),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1707),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1690),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1743),
.A2(n_1747),
.B(n_1757),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1757),
.A2(n_1666),
.B(n_1750),
.Y(n_1809)
);

OR2x6_ASAP7_75t_L g1810 ( 
.A(n_1755),
.B(n_1680),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_R g1811 ( 
.A(n_1685),
.B(n_1702),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1694),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1668),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1753),
.B(n_1761),
.Y(n_1814)
);

AO21x1_ASAP7_75t_SL g1815 ( 
.A1(n_1720),
.A2(n_1771),
.B(n_1764),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1656),
.B(n_1737),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1713),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1713),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1740),
.B(n_1767),
.Y(n_1819)
);

BUFx4f_ASAP7_75t_SL g1820 ( 
.A(n_1729),
.Y(n_1820)
);

OA21x2_ASAP7_75t_L g1821 ( 
.A1(n_1728),
.A2(n_1714),
.B(n_1672),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1769),
.B(n_1748),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1666),
.A2(n_1732),
.B(n_1680),
.Y(n_1823)
);

NAND2x1_ASAP7_75t_L g1824 ( 
.A(n_1723),
.B(n_1748),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1714),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1659),
.B(n_1676),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1704),
.Y(n_1827)
);

INVxp67_ASAP7_75t_SL g1828 ( 
.A(n_1692),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1653),
.B(n_1772),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1704),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1731),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1692),
.Y(n_1832)
);

OR2x6_ASAP7_75t_L g1833 ( 
.A(n_1700),
.B(n_1716),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1700),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1762),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1734),
.B(n_1760),
.Y(n_1836)
);

CKINVDCx20_ASAP7_75t_R g1837 ( 
.A(n_1655),
.Y(n_1837)
);

OA21x2_ASAP7_75t_L g1838 ( 
.A1(n_1715),
.A2(n_1706),
.B(n_1730),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1724),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1722),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1716),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1741),
.B(n_1765),
.Y(n_1842)
);

BUFx2_ASAP7_75t_L g1843 ( 
.A(n_1673),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_SL g1844 ( 
.A(n_1695),
.B(n_1703),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1647),
.B(n_1770),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1697),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1801),
.A2(n_1669),
.B1(n_1675),
.B2(n_1754),
.C(n_1654),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1783),
.B(n_1725),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1822),
.B(n_1718),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1783),
.B(n_1701),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1783),
.B(n_1701),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1800),
.B(n_1647),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1823),
.A2(n_1770),
.B1(n_1670),
.B2(n_1721),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1788),
.A2(n_1709),
.B(n_1687),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1796),
.B(n_1727),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1835),
.B(n_1706),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1774),
.B(n_1780),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1835),
.B(n_1843),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1780),
.B(n_1794),
.Y(n_1859)
);

AOI21xp33_ASAP7_75t_L g1860 ( 
.A1(n_1808),
.A2(n_1809),
.B(n_1828),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1782),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1773),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1788),
.A2(n_1810),
.B1(n_1826),
.B2(n_1777),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1831),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1775),
.Y(n_1865)
);

INVx4_ASAP7_75t_L g1866 ( 
.A(n_1787),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1843),
.B(n_1708),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1790),
.B(n_1699),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1798),
.B(n_1759),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1810),
.A2(n_1705),
.B1(n_1658),
.B2(n_1759),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1790),
.B(n_1838),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1810),
.A2(n_1678),
.B1(n_1744),
.B2(n_1763),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1813),
.B(n_1651),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1784),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1784),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1790),
.B(n_1678),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1825),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1825),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1792),
.Y(n_1879)
);

AOI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1832),
.A2(n_1766),
.B(n_1662),
.Y(n_1880)
);

NAND2x1p5_ASAP7_75t_L g1881 ( 
.A(n_1824),
.B(n_1662),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1877),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1867),
.B(n_1781),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1864),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1860),
.A2(n_1810),
.B1(n_1863),
.B2(n_1852),
.Y(n_1885)
);

NAND3xp33_ASAP7_75t_L g1886 ( 
.A(n_1860),
.B(n_1840),
.C(n_1841),
.Y(n_1886)
);

AND2x6_ASAP7_75t_SL g1887 ( 
.A(n_1855),
.B(n_1779),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1863),
.A2(n_1787),
.B(n_1852),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1862),
.Y(n_1889)
);

NAND4xp25_ASAP7_75t_L g1890 ( 
.A(n_1847),
.B(n_1836),
.C(n_1814),
.D(n_1776),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1855),
.B(n_1804),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_R g1892 ( 
.A(n_1853),
.B(n_1837),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1867),
.B(n_1815),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1854),
.B(n_1789),
.Y(n_1894)
);

OAI211xp5_ASAP7_75t_L g1895 ( 
.A1(n_1847),
.A2(n_1791),
.B(n_1786),
.C(n_1834),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1864),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1868),
.B(n_1815),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1859),
.B(n_1802),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1853),
.A2(n_1833),
.B1(n_1795),
.B2(n_1839),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1865),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1868),
.B(n_1857),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1873),
.A2(n_1778),
.B(n_1849),
.C(n_1870),
.Y(n_1902)
);

OAI33xp33_ASAP7_75t_L g1903 ( 
.A1(n_1873),
.A2(n_1812),
.A3(n_1805),
.B1(n_1807),
.B2(n_1803),
.B3(n_1816),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1870),
.A2(n_1795),
.B1(n_1833),
.B2(n_1837),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1868),
.B(n_1857),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1854),
.A2(n_1833),
.B1(n_1797),
.B2(n_1819),
.Y(n_1906)
);

OAI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1866),
.A2(n_1833),
.B1(n_1827),
.B2(n_1830),
.Y(n_1907)
);

NAND3xp33_ASAP7_75t_SL g1908 ( 
.A(n_1872),
.B(n_1785),
.C(n_1811),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1865),
.Y(n_1909)
);

OAI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1881),
.A2(n_1819),
.B1(n_1824),
.B2(n_1786),
.C(n_1791),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1880),
.A2(n_1820),
.B1(n_1789),
.B2(n_1791),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1879),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1862),
.B(n_1793),
.Y(n_1913)
);

AOI222xp33_ASAP7_75t_L g1914 ( 
.A1(n_1872),
.A2(n_1844),
.B1(n_1851),
.B2(n_1850),
.C1(n_1842),
.C2(n_1829),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1857),
.B(n_1846),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1861),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1869),
.B(n_1806),
.Y(n_1917)
);

AND2x2_ASAP7_75t_SL g1918 ( 
.A(n_1866),
.B(n_1821),
.Y(n_1918)
);

BUFx2_ASAP7_75t_L g1919 ( 
.A(n_1862),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1866),
.A2(n_1845),
.B1(n_1818),
.B2(n_1817),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1862),
.B(n_1793),
.Y(n_1921)
);

NOR2x1p5_ASAP7_75t_L g1922 ( 
.A(n_1908),
.B(n_1797),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1888),
.B(n_1881),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1912),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1917),
.B(n_1849),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1912),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1897),
.B(n_1858),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1884),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1896),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1891),
.B(n_1799),
.Y(n_1930)
);

AOI21x1_ASAP7_75t_L g1931 ( 
.A1(n_1889),
.A2(n_1877),
.B(n_1878),
.Y(n_1931)
);

OA21x2_ASAP7_75t_L g1932 ( 
.A1(n_1910),
.A2(n_1871),
.B(n_1848),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1895),
.A2(n_1848),
.B(n_1851),
.Y(n_1933)
);

INVxp67_ASAP7_75t_SL g1934 ( 
.A(n_1900),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1906),
.B(n_1881),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1919),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1916),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1909),
.Y(n_1938)
);

NAND3xp33_ASAP7_75t_L g1939 ( 
.A(n_1886),
.B(n_1851),
.C(n_1876),
.Y(n_1939)
);

INVx4_ASAP7_75t_SL g1940 ( 
.A(n_1913),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1909),
.Y(n_1941)
);

INVx4_ASAP7_75t_L g1942 ( 
.A(n_1887),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1913),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1919),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1913),
.B(n_1921),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1914),
.B(n_1866),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1901),
.B(n_1874),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1915),
.B(n_1875),
.Y(n_1948)
);

OR2x6_ASAP7_75t_L g1949 ( 
.A(n_1904),
.B(n_1881),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1882),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1915),
.B(n_1875),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1901),
.B(n_1856),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1932),
.B(n_1905),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1932),
.B(n_1905),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1932),
.B(n_1918),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1936),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1932),
.B(n_1918),
.Y(n_1957)
);

INVx1_ASAP7_75t_SL g1958 ( 
.A(n_1936),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1928),
.B(n_1898),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1924),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1952),
.B(n_1893),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1952),
.B(n_1893),
.Y(n_1962)
);

INVx4_ASAP7_75t_L g1963 ( 
.A(n_1942),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1933),
.B(n_1940),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1941),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1924),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1950),
.Y(n_1967)
);

NAND2xp33_ASAP7_75t_SL g1968 ( 
.A(n_1942),
.B(n_1922),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1926),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1934),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1926),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1931),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1940),
.B(n_1883),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1940),
.B(n_1927),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1938),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1944),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1937),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1939),
.A2(n_1885),
.B(n_1903),
.Y(n_1978)
);

AOI33xp33_ASAP7_75t_L g1979 ( 
.A1(n_1939),
.A2(n_1911),
.A3(n_1899),
.B1(n_1907),
.B2(n_1876),
.B3(n_1920),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1942),
.A2(n_1890),
.B1(n_1892),
.B2(n_1902),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1923),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1937),
.B(n_1929),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1968),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1960),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1974),
.B(n_1943),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1960),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1966),
.Y(n_1987)
);

OAI21xp33_ASAP7_75t_L g1988 ( 
.A1(n_1979),
.A2(n_1980),
.B(n_1978),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1980),
.B(n_1942),
.Y(n_1989)
);

INVx4_ASAP7_75t_L g1990 ( 
.A(n_1963),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1966),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1969),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1969),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1971),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1961),
.Y(n_1995)
);

AOI322xp5_ASAP7_75t_L g1996 ( 
.A1(n_1955),
.A2(n_1946),
.A3(n_1894),
.B1(n_1925),
.B2(n_1947),
.C1(n_1944),
.C2(n_1930),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1971),
.Y(n_1997)
);

INVx2_ASAP7_75t_SL g1998 ( 
.A(n_1974),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1974),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1977),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1973),
.B(n_1943),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1961),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1963),
.B(n_1943),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1975),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1968),
.A2(n_1922),
.B1(n_1923),
.B2(n_1949),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1979),
.B(n_1947),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1967),
.B(n_1970),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1977),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1963),
.B(n_1945),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1961),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1982),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1967),
.Y(n_2012)
);

NOR2x1_ASAP7_75t_L g2013 ( 
.A(n_1963),
.B(n_1938),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1982),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1962),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1962),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1956),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1978),
.B(n_1948),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1962),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1970),
.B(n_1951),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1959),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1973),
.B(n_1945),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1956),
.B(n_1945),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1988),
.B(n_1963),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2012),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1990),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_2022),
.B(n_1973),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1995),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1989),
.A2(n_1949),
.B1(n_1935),
.B2(n_1923),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2017),
.B(n_1958),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_2013),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2007),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_2007),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1984),
.Y(n_2034)
);

NAND2x1_ASAP7_75t_L g2035 ( 
.A(n_2013),
.B(n_1964),
.Y(n_2035)
);

AND3x2_ASAP7_75t_L g2036 ( 
.A(n_2003),
.B(n_1981),
.C(n_1976),
.Y(n_2036)
);

INVx5_ASAP7_75t_L g2037 ( 
.A(n_1990),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1995),
.B(n_1958),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_2006),
.A2(n_1949),
.B1(n_1935),
.B2(n_1923),
.Y(n_2039)
);

BUFx3_ASAP7_75t_L g2040 ( 
.A(n_2004),
.Y(n_2040)
);

INVx1_ASAP7_75t_SL g2041 ( 
.A(n_1983),
.Y(n_2041)
);

INVxp67_ASAP7_75t_SL g2042 ( 
.A(n_1998),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2018),
.B(n_1965),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1984),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_2004),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_1998),
.Y(n_2046)
);

BUFx2_ASAP7_75t_L g2047 ( 
.A(n_1999),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1986),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1986),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1987),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_1999),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_2022),
.A2(n_1949),
.B1(n_1935),
.B2(n_1923),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2002),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2027),
.B(n_1985),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2041),
.B(n_2033),
.Y(n_2055)
);

AOI211xp5_ASAP7_75t_L g2056 ( 
.A1(n_2024),
.A2(n_2009),
.B(n_2005),
.C(n_1955),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_2041),
.B(n_1990),
.Y(n_2057)
);

OAI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2035),
.A2(n_1949),
.B1(n_1935),
.B2(n_1981),
.Y(n_2058)
);

AOI21xp33_ASAP7_75t_L g2059 ( 
.A1(n_2030),
.A2(n_2042),
.B(n_2035),
.Y(n_2059)
);

NOR2xp67_ASAP7_75t_SL g2060 ( 
.A(n_2037),
.B(n_1975),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2047),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2047),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2032),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_2043),
.B(n_1996),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_SL g2065 ( 
.A1(n_2039),
.A2(n_1957),
.B1(n_1955),
.B2(n_1964),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_2045),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2032),
.Y(n_2067)
);

NOR4xp25_ASAP7_75t_L g2068 ( 
.A(n_2025),
.B(n_2051),
.C(n_2046),
.D(n_2031),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2027),
.B(n_1985),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2034),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2034),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2025),
.A2(n_1957),
.B(n_1964),
.C(n_2023),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2044),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_2046),
.Y(n_2074)
);

NAND2x1_ASAP7_75t_L g2075 ( 
.A(n_2031),
.B(n_2001),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2040),
.B(n_2001),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2061),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2074),
.B(n_2051),
.Y(n_2078)
);

OAI21xp5_ASAP7_75t_SL g2079 ( 
.A1(n_2064),
.A2(n_2036),
.B(n_2029),
.Y(n_2079)
);

OAI221xp5_ASAP7_75t_L g2080 ( 
.A1(n_2064),
.A2(n_2052),
.B1(n_2038),
.B2(n_1981),
.C(n_2040),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2062),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_2068),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2055),
.B(n_2038),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2066),
.B(n_2040),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2054),
.Y(n_2085)
);

NAND2xp33_ASAP7_75t_SL g2086 ( 
.A(n_2060),
.B(n_2075),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2063),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2067),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2070),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2071),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2054),
.B(n_2020),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_2057),
.B(n_2037),
.Y(n_2092)
);

NOR3x1_ASAP7_75t_L g2093 ( 
.A(n_2079),
.B(n_2073),
.C(n_2048),
.Y(n_2093)
);

NAND3xp33_ASAP7_75t_SL g2094 ( 
.A(n_2082),
.B(n_2056),
.C(n_2072),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2085),
.B(n_2076),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_2083),
.B(n_2057),
.Y(n_2096)
);

NOR3xp33_ASAP7_75t_L g2097 ( 
.A(n_2080),
.B(n_2059),
.C(n_2026),
.Y(n_2097)
);

O2A1O1Ixp33_ASAP7_75t_L g2098 ( 
.A1(n_2082),
.A2(n_2058),
.B(n_2026),
.C(n_1972),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2078),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2086),
.A2(n_2069),
.B1(n_2076),
.B2(n_2065),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2086),
.A2(n_2069),
.B1(n_2060),
.B2(n_1957),
.Y(n_2101)
);

AOI211xp5_ASAP7_75t_L g2102 ( 
.A1(n_2084),
.A2(n_2026),
.B(n_2050),
.C(n_2049),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2077),
.B(n_2026),
.Y(n_2103)
);

OAI221xp5_ASAP7_75t_L g2104 ( 
.A1(n_2092),
.A2(n_2037),
.B1(n_2028),
.B2(n_2053),
.C(n_1972),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2081),
.B(n_2002),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2094),
.A2(n_2097),
.B1(n_2096),
.B2(n_2100),
.Y(n_2106)
);

AOI21xp33_ASAP7_75t_L g2107 ( 
.A1(n_2098),
.A2(n_2092),
.B(n_2091),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2095),
.Y(n_2108)
);

AOI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_2101),
.A2(n_2088),
.B(n_2087),
.Y(n_2109)
);

O2A1O1Ixp33_ASAP7_75t_L g2110 ( 
.A1(n_2104),
.A2(n_2090),
.B(n_2089),
.C(n_2049),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2105),
.Y(n_2111)
);

OAI21xp33_ASAP7_75t_SL g2112 ( 
.A1(n_2103),
.A2(n_2053),
.B(n_2028),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2108),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2112),
.Y(n_2114)
);

OAI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_2106),
.A2(n_2099),
.B(n_2102),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_L g2116 ( 
.A(n_2107),
.B(n_2037),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2110),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2111),
.B(n_2093),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2109),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2118),
.Y(n_2120)
);

OAI221xp5_ASAP7_75t_L g2121 ( 
.A1(n_2115),
.A2(n_2037),
.B1(n_2053),
.B2(n_2028),
.C(n_2044),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2114),
.Y(n_2122)
);

A2O1A1Ixp33_ASAP7_75t_L g2123 ( 
.A1(n_2116),
.A2(n_2037),
.B(n_2048),
.C(n_2050),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_L g2124 ( 
.A(n_2119),
.B(n_1975),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2113),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2120),
.Y(n_2126)
);

NAND4xp75_ASAP7_75t_L g2127 ( 
.A(n_2122),
.B(n_2116),
.C(n_2117),
.D(n_2021),
.Y(n_2127)
);

AOI211x1_ASAP7_75t_L g2128 ( 
.A1(n_2121),
.A2(n_2021),
.B(n_2014),
.C(n_2011),
.Y(n_2128)
);

XOR2x2_ASAP7_75t_L g2129 ( 
.A(n_2127),
.B(n_2124),
.Y(n_2129)
);

AOI322xp5_ASAP7_75t_L g2130 ( 
.A1(n_2129),
.A2(n_2126),
.A3(n_2125),
.B1(n_2123),
.B2(n_2128),
.C1(n_1953),
.C2(n_1954),
.Y(n_2130)
);

OR3x1_ASAP7_75t_L g2131 ( 
.A(n_2130),
.B(n_2014),
.C(n_2011),
.Y(n_2131)
);

OA21x2_ASAP7_75t_L g2132 ( 
.A1(n_2130),
.A2(n_2008),
.B(n_2000),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2132),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_2132),
.B(n_2010),
.Y(n_2134)
);

OAI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_2134),
.A2(n_2131),
.B(n_2008),
.Y(n_2135)
);

OAI22x1_ASAP7_75t_SL g2136 ( 
.A1(n_2133),
.A2(n_2019),
.B1(n_2016),
.B2(n_2015),
.Y(n_2136)
);

AOI221xp5_ASAP7_75t_L g2137 ( 
.A1(n_2136),
.A2(n_2000),
.B1(n_1991),
.B2(n_1994),
.C(n_1992),
.Y(n_2137)
);

CKINVDCx20_ASAP7_75t_R g2138 ( 
.A(n_2137),
.Y(n_2138)
);

AOI21xp33_ASAP7_75t_L g2139 ( 
.A1(n_2138),
.A2(n_2135),
.B(n_1991),
.Y(n_2139)
);

AOI22x1_ASAP7_75t_L g2140 ( 
.A1(n_2139),
.A2(n_1987),
.B1(n_1992),
.B2(n_1993),
.Y(n_2140)
);

AOI22xp5_ASAP7_75t_L g2141 ( 
.A1(n_2140),
.A2(n_2019),
.B1(n_2016),
.B2(n_2015),
.Y(n_2141)
);

AOI211xp5_ASAP7_75t_L g2142 ( 
.A1(n_2141),
.A2(n_1997),
.B(n_1994),
.C(n_1993),
.Y(n_2142)
);


endmodule