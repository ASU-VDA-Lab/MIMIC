module fake_jpeg_13565_n_426 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_50),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_15),
.C(n_14),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_79),
.C(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_0),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_59),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_18),
.B(n_33),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_60),
.B(n_26),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_65),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_70),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_66),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_13),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_16),
.B(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_76),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_21),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_91),
.B(n_68),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_30),
.B1(n_40),
.B2(n_36),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_101),
.B1(n_103),
.B2(n_107),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_95),
.A2(n_96),
.B1(n_111),
.B2(n_128),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_42),
.B1(n_40),
.B2(n_36),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_30),
.B1(n_40),
.B2(n_36),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_109),
.A2(n_122),
.B1(n_83),
.B2(n_80),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_42),
.B1(n_31),
.B2(n_26),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_32),
.B1(n_27),
.B2(n_24),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_72),
.C(n_87),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_26),
.B1(n_17),
.B2(n_23),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_52),
.A2(n_17),
.B1(n_23),
.B2(n_22),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_129),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_47),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_50),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_58),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_141),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_86),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_142),
.B(n_154),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_69),
.C(n_78),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_143),
.B(n_147),
.C(n_163),
.Y(n_221)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_89),
.A2(n_49),
.B(n_48),
.C(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_146),
.B(n_160),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_94),
.B(n_77),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

BUFx4f_ASAP7_75t_SL g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_61),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_151),
.B(n_161),
.Y(n_218)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_153),
.B(n_158),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_71),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_57),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_155),
.B(n_156),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_104),
.B(n_131),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_12),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_159),
.B(n_162),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_46),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_126),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_102),
.B(n_11),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_164),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_172),
.B1(n_186),
.B2(n_189),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_187),
.B1(n_191),
.B2(n_140),
.Y(n_212)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_93),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_93),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_68),
.B(n_125),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_10),
.Y(n_182)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_118),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_184),
.B(n_188),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_98),
.B(n_74),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_4),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_100),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_53),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_116),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_202),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_147),
.B1(n_151),
.B2(n_143),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_203),
.A2(n_228),
.B(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_150),
.A2(n_130),
.B1(n_117),
.B2(n_110),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_222),
.B1(n_185),
.B2(n_175),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_176),
.A2(n_63),
.B1(n_54),
.B2(n_45),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_210),
.B1(n_215),
.B2(n_219),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_44),
.B1(n_62),
.B2(n_117),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_212),
.B(n_157),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_119),
.B1(n_133),
.B2(n_140),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_171),
.A2(n_119),
.B1(n_116),
.B2(n_123),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_147),
.A2(n_123),
.B1(n_59),
.B2(n_67),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_188),
.C(n_189),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_146),
.A2(n_187),
.B1(n_163),
.B2(n_160),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_215),
.B1(n_221),
.B2(n_194),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_125),
.B(n_6),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_184),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_196),
.B(n_149),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_236),
.B(n_244),
.Y(n_282)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_240),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_152),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_247),
.C(n_269),
.Y(n_277)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_241),
.B(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_202),
.Y(n_243)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_243),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_149),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_253),
.B1(n_257),
.B2(n_270),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_195),
.A2(n_173),
.B1(n_148),
.B2(n_145),
.Y(n_246)
);

OAI22x1_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_256),
.B1(n_213),
.B2(n_201),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_166),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_186),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_248),
.B(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_251),
.A2(n_267),
.B1(n_193),
.B2(n_269),
.Y(n_303)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_203),
.A2(n_144),
.B1(n_167),
.B2(n_169),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_168),
.B(n_178),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_255),
.A2(n_193),
.B(n_238),
.Y(n_308)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_205),
.A2(n_174),
.B1(n_179),
.B2(n_9),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_7),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_206),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_264),
.Y(n_304)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_7),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_202),
.A2(n_8),
.B(n_228),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_271),
.B(n_273),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_230),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_206),
.Y(n_268)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_223),
.B(n_216),
.C(n_219),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_199),
.A2(n_222),
.B1(n_207),
.B2(n_210),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_SL g271 ( 
.A(n_198),
.B(n_233),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_272),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_234),
.A2(n_227),
.B(n_199),
.C(n_232),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_217),
.C(n_214),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_217),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_275),
.B(n_285),
.Y(n_310)
);

CKINVDCx6p67_ASAP7_75t_R g328 ( 
.A(n_280),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_287),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_254),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_300),
.B1(n_303),
.B2(n_308),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_295),
.B(n_296),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_214),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_238),
.A2(n_198),
.B(n_209),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_297),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_213),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_302),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_254),
.A2(n_208),
.B1(n_211),
.B2(n_224),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_224),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_288),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_312),
.Y(n_341)
);

OAI32xp33_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_273),
.A3(n_243),
.B1(n_255),
.B2(n_253),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_270),
.B1(n_249),
.B2(n_257),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_315),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_291),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_276),
.A2(n_249),
.B1(n_271),
.B2(n_274),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_320),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_282),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_292),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_193),
.B1(n_272),
.B2(n_306),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_323),
.A2(n_326),
.B1(n_335),
.B2(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_302),
.B1(n_283),
.B2(n_304),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_287),
.B(n_304),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_307),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_330),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_298),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_331),
.Y(n_340)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_278),
.B(n_283),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_334),
.A2(n_277),
.B(n_278),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_297),
.B1(n_285),
.B2(n_289),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_337),
.B(n_358),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_324),
.A2(n_277),
.B(n_280),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_328),
.B(n_333),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_275),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_349),
.C(n_355),
.Y(n_371)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_324),
.A2(n_296),
.B(n_286),
.Y(n_346)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

OAI21xp33_ASAP7_75t_L g348 ( 
.A1(n_320),
.A2(n_313),
.B(n_316),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_323),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_305),
.C(n_290),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_319),
.B(n_290),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_352),
.B(n_318),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_326),
.A2(n_316),
.B(n_322),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_353),
.A2(n_322),
.B(n_329),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_354),
.A2(n_312),
.B1(n_328),
.B2(n_332),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_335),
.C(n_329),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_356),
.Y(n_359)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_327),
.Y(n_357)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_345),
.A2(n_328),
.B1(n_334),
.B2(n_314),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_363),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_341),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_373),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_341),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_366),
.B(n_372),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_354),
.A2(n_321),
.B1(n_315),
.B2(n_309),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_SL g382 ( 
.A1(n_369),
.A2(n_370),
.B(n_344),
.C(n_336),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_328),
.B(n_353),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_358),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_355),
.C(n_352),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_350),
.B(n_340),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_377),
.Y(n_385)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_376),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_369),
.C(n_362),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_367),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_384),
.B(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_359),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_388),
.B(n_392),
.Y(n_401)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_365),
.Y(n_395)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_374),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_371),
.C(n_373),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_402),
.C(n_340),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_371),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_396),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_379),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_377),
.C(n_360),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_400),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_349),
.B(n_339),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_398),
.A2(n_403),
.B(n_397),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_364),
.C(n_345),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_387),
.A2(n_370),
.B(n_368),
.C(n_376),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_402),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_394),
.A2(n_391),
.B(n_378),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_409),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_406),
.B(n_408),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_391),
.C(n_390),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_403),
.A2(n_336),
.B(n_382),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_411),
.B(n_342),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_414),
.B(n_415),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_407),
.A2(n_399),
.B1(n_351),
.B2(n_401),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_416),
.A2(n_411),
.B(n_407),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_418),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_351),
.B1(n_347),
.B2(n_338),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_SL g421 ( 
.A1(n_419),
.A2(n_382),
.B(n_413),
.C(n_356),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_421),
.A2(n_417),
.B(n_412),
.Y(n_422)
);

AO21x1_ASAP7_75t_L g423 ( 
.A1(n_422),
.A2(n_420),
.B(n_410),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_382),
.B(n_347),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_338),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_357),
.Y(n_426)
);


endmodule