module fake_jpeg_721_n_190 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_0),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_2),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_63),
.B1(n_59),
.B2(n_56),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_45),
.B1(n_50),
.B2(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_92),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_63),
.B1(n_59),
.B2(n_56),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_58),
.B1(n_52),
.B2(n_62),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_61),
.C(n_44),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_53),
.C(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_61),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_65),
.B1(n_62),
.B2(n_52),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_72),
.B1(n_57),
.B2(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_57),
.B1(n_65),
.B2(n_64),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_97),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_119),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_108),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_72),
.B1(n_45),
.B2(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_45),
.B(n_75),
.C(n_49),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_3),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_72),
.B1(n_49),
.B2(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_72),
.B1(n_41),
.B2(n_39),
.Y(n_130)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_91),
.Y(n_121)
);

XOR2x1_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_5),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_131),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_84),
.B(n_85),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_7),
.B(n_9),
.Y(n_153)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_90),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_129),
.Y(n_146)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_5),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_2),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_3),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_38),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_115),
.C(n_6),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_115),
.B1(n_107),
.B2(n_6),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_151),
.B1(n_144),
.B2(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_157),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_145),
.C(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_154),
.B1(n_14),
.B2(n_15),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_37),
.C(n_36),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_130),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_153),
.A2(n_10),
.B(n_13),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_164),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_159),
.B(n_152),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_137),
.C(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_161),
.C(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_120),
.C(n_23),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_163),
.B(n_153),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_134),
.B(n_125),
.C(n_25),
.D(n_27),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_34),
.C(n_32),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_140),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_134),
.B1(n_15),
.B2(n_17),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_148),
.B1(n_152),
.B2(n_18),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_159),
.Y(n_177)
);

AOI321xp33_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_149),
.A3(n_143),
.B1(n_155),
.B2(n_142),
.C(n_145),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_174),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_26),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_179),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_173),
.A2(n_163),
.B1(n_167),
.B2(n_169),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_170),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_183),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_182),
.B(n_179),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_186),
.B(n_178),
.CI(n_17),
.CON(n_187),
.SN(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_187),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_187),
.C(n_20),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_20),
.Y(n_190)
);


endmodule