module real_jpeg_4649_n_31 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_29, n_10, n_186, n_9, n_12, n_24, n_189, n_187, n_6, n_190, n_28, n_183, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_26, n_27, n_20, n_19, n_182, n_184, n_30, n_16, n_15, n_13, n_31);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_29;
input n_10;
input n_186;
input n_9;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_28;
input n_183;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_182;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_173;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_0),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_0),
.B(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_0),
.B(n_48),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_0),
.A2(n_45),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_1),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_2),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_3),
.B(n_67),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_4),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_6),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_6),
.B(n_64),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_8),
.B(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_10),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_11),
.Y(n_177)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_12),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_13),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_13),
.B(n_81),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_15),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_15),
.B(n_55),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_16),
.B(n_105),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_17),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_18),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_21),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_78),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_22),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_23),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_27),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_27),
.B(n_163),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_29),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_29),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_174),
.Y(n_31)
);

AO21x1_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_41),
.B(n_172),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_35),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_65),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_37),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_37),
.B(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_40),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_171),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_43),
.B(n_45),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_45),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_170),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_158),
.B(n_167),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_133),
.B(n_152),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_72),
.B(n_120),
.C(n_129),
.Y(n_52)
);

NOR4xp25_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.C(n_63),
.D(n_66),
.Y(n_53)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_112),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_63),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_79),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_101),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_115),
.B(n_119),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_110),
.B(n_114),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B(n_83),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_94),
.B(n_109),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_93),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_104),
.B(n_108),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B(n_103),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_113),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B(n_126),
.C(n_127),
.D(n_128),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.C(n_148),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_148),
.B(n_153),
.C(n_156),
.D(n_157),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_181),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_182),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_183),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_184),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_185),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_186),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_187),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_188),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_189),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_190),
.Y(n_117)
);


endmodule