module fake_jpeg_25255_n_81 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_56),
.B(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_65),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_15),
.C(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_69),
.C(n_64),
.Y(n_72)
);

BUFx12f_ASAP7_75t_SL g74 ( 
.A(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_73),
.B1(n_58),
.B2(n_54),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_57),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);


endmodule