module real_jpeg_33417_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_11;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_0),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_0),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_2),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_2),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_3),
.A2(n_53),
.B1(n_90),
.B2(n_93),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_3),
.A2(n_53),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_4),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_5),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_7),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

OAI22x1_ASAP7_75t_SL g41 ( 
.A1(n_8),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_46),
.B1(n_60),
.B2(n_64),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_46),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

INVx2_ASAP7_75t_R g142 ( 
.A(n_8),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_8),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_8),
.B(n_56),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_88),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_189),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_187),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_149),
.Y(n_11)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_12),
.B(n_149),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_57),
.C(n_96),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_15),
.A2(n_58),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_40),
.B1(n_49),
.B2(n_55),
.Y(n_15)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_16),
.A2(n_40),
.B1(n_49),
.B2(n_55),
.Y(n_151)
);

NAND2x1p5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_30),
.Y(n_16)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

AOI22x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_34),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

OAI211xp5_ASAP7_75t_SL g120 ( 
.A1(n_46),
.A2(n_121),
.B(n_124),
.C(n_127),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_46),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_46),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_58),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_58),
.A2(n_194),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AO22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_67),
.B1(n_88),
.B2(n_89),
.Y(n_58)
);

AO22x2_ASAP7_75t_L g184 ( 
.A1(n_59),
.A2(n_67),
.B1(n_88),
.B2(n_89),
.Y(n_184)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_60),
.Y(n_221)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

AOI21x1_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_74),
.B(n_81),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_68),
.A2(n_213),
.B1(n_218),
.B2(n_222),
.Y(n_212)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_85),
.Y(n_224)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_97),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_147),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_120),
.C(n_132),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_133),
.B(n_148),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_100),
.A2(n_133),
.B(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_101),
.A2(n_200),
.B1(n_201),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_102),
.B(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_102),
.B(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_111),
.Y(n_200)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_113),
.B(n_142),
.Y(n_230)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_182),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_181),
.Y(n_150)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_166),
.B2(n_167),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AO22x2_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_161),
.B2(n_163),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_166),
.B(n_210),
.Y(n_238)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_R g245 ( 
.A(n_171),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_184),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_197),
.C(n_206),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_207),
.B(n_247),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_192),
.B(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_211),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B(n_202),
.Y(n_199)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_243),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_239),
.B(n_246),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_225),
.B(n_238),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_228),
.B(n_237),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);


endmodule