module fake_jpeg_30094_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_0),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_64),
.A2(n_55),
.B1(n_54),
.B2(n_48),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_1),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_45),
.B1(n_52),
.B2(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_26),
.B1(n_37),
.B2(n_36),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_52),
.B1(n_53),
.B2(n_50),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_6),
.C(n_7),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_42),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_20),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_1),
.CI(n_2),
.CON(n_83),
.SN(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_49),
.B1(n_55),
.B2(n_51),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_16),
.B1(n_39),
.B2(n_38),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_90),
.B1(n_76),
.B2(n_9),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_14),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_3),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_8),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_91),
.B(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_99),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_76),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_10),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_75),
.C(n_27),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.C(n_83),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_21),
.C(n_34),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_113),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_114),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_86),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_118),
.C(n_107),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_106),
.B1(n_100),
.B2(n_29),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_118)
);

NOR4xp25_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_101),
.C(n_93),
.D(n_96),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_116),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_123),
.B(n_119),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_125),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_115),
.B1(n_110),
.B2(n_108),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_126),
.B(n_111),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_124),
.A3(n_28),
.B1(n_30),
.B2(n_31),
.C1(n_40),
.C2(n_18),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_117),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule