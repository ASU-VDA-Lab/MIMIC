module fake_netlist_6_161_n_1915 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1915);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1915;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_175),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_165),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_56),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_30),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_25),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_28),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_105),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_117),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_85),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_23),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_25),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_53),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_106),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_8),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_125),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_51),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_31),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_53),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_87),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_29),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_107),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_55),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_52),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_98),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_68),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_76),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_133),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_16),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_35),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_69),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_32),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_31),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_35),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_32),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_1),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_10),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_88),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_91),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_36),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_54),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_118),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_81),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_120),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_54),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_139),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_84),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_100),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_48),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_22),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_75),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_65),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_40),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_27),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_52),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_57),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_18),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_90),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_24),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_160),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_78),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_140),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_162),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_29),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_108),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_59),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_93),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_8),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_34),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_143),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_171),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_11),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_176),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_166),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_137),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_13),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_122),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_161),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_66),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_46),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_40),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_169),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_50),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_47),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_28),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_163),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_154),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_62),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_24),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_70),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_72),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_2),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_22),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_111),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_128),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_38),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_15),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_48),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_77),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_156),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_71),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_145),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_157),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_151),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_67),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_132),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_55),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_43),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_101),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_38),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_64),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_73),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_89),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_7),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_41),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_11),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_135),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_95),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_99),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_136),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_17),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_62),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_82),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_50),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_147),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_129),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_116),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_63),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_5),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_115),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_142),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_4),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_26),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_152),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_14),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_57),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_13),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_18),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_4),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_42),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_37),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_180),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_179),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_184),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_209),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_297),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_226),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_205),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_275),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_217),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_217),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_186),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_185),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_195),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_287),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_188),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_187),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_218),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_190),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_193),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_287),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_302),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_322),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_195),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_342),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_199),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_200),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_186),
.B(n_6),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_192),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_6),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_192),
.B(n_7),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_205),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_194),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_226),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_207),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_219),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_273),
.B(n_12),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_273),
.B(n_12),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_194),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_197),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_181),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_202),
.B(n_14),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_220),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_245),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_208),
.B(n_16),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_197),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_201),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_247),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_226),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_201),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_204),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_204),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_251),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_255),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_182),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_215),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_340),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_240),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_215),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_240),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_228),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_256),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_228),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_183),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_235),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_196),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_235),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_237),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_264),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_237),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_270),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_293),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_253),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_293),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_253),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_271),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_198),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_446),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_426),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_446),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_446),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_363),
.B(n_272),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_446),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_446),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_363),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_363),
.B(n_198),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_198),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_359),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_362),
.B(n_379),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

NOR2x1_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_241),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_361),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_400),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_366),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_357),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_362),
.B(n_223),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_404),
.B(n_198),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_277),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_366),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_428),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_360),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_396),
.B(n_241),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_377),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_198),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_371),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_399),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_379),
.B(n_394),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_378),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_378),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_280),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_198),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_405),
.B(n_189),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_381),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_383),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_364),
.B(n_304),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_364),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_385),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_385),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_364),
.B(n_281),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_409),
.B(n_283),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_392),
.B(n_304),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_335),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_387),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_390),
.Y(n_508)
);

AND2x4_ASAP7_75t_SL g509 ( 
.A(n_408),
.B(n_223),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_390),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_391),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_435),
.B(n_335),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_369),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_397),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_412),
.B(n_223),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_370),
.B(n_351),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_406),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_392),
.B(n_211),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_382),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_477),
.B(n_384),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_491),
.B(n_373),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_477),
.B(n_365),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_470),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_497),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_497),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_497),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_491),
.B(n_375),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_449),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_465),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_465),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_519),
.A2(n_489),
.B1(n_469),
.B2(n_502),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_497),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_452),
.B(n_471),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_258),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_504),
.B(n_211),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_456),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_509),
.B(n_376),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_502),
.B(n_432),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_517),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_514),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_452),
.B(n_388),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_518),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_449),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_202),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_505),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_518),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_518),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_471),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_467),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_468),
.B(n_395),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_519),
.A2(n_395),
.B1(n_401),
.B2(n_260),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_469),
.A2(n_260),
.B1(n_282),
.B2(n_258),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_456),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_500),
.B(n_389),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_487),
.B(n_402),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_467),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_504),
.B(n_210),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_505),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_520),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_403),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_504),
.B(n_211),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_479),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_509),
.B(n_410),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_455),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_509),
.A2(n_441),
.B1(n_443),
.B2(n_356),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_475),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_509),
.B(n_411),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_454),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_522),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_416),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_461),
.B(n_421),
.Y(n_602)
);

NOR2x1p5_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_282),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_468),
.B(n_422),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_463),
.B(n_434),
.C(n_423),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_496),
.B(n_407),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_483),
.B(n_203),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_455),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_461),
.B(n_430),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_463),
.B(n_440),
.C(n_438),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_475),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_516),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_457),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_516),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_512),
.B(n_445),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_484),
.B(n_443),
.C(n_441),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_466),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_252),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_516),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_496),
.B(n_211),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_475),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_516),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_466),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_516),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_521),
.B(n_429),
.C(n_368),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_496),
.B(n_318),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_466),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_515),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_466),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_489),
.B(n_320),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_479),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_521),
.B(n_211),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_481),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_457),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_515),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_484),
.B(n_372),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_454),
.Y(n_641)
);

OR2x2_ASAP7_75t_SL g642 ( 
.A(n_481),
.B(n_285),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_521),
.A2(n_310),
.B1(n_323),
.B2(n_330),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_515),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_472),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_512),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_524),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_472),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_524),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_512),
.B(n_447),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_447),
.B(n_334),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_472),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_472),
.Y(n_653)
);

INVxp33_ASAP7_75t_SL g654 ( 
.A(n_483),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_524),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_523),
.B(n_223),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_447),
.B(n_286),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_508),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_450),
.B(n_288),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_454),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_458),
.B(n_413),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_523),
.B(n_292),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_523),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_458),
.B(n_374),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_458),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_454),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_462),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_450),
.B(n_296),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_462),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_523),
.B(n_368),
.Y(n_671)
);

AOI21x1_ASAP7_75t_L g672 ( 
.A1(n_450),
.A2(n_212),
.B(n_210),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_462),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_523),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_506),
.B(n_300),
.Y(n_675)
);

CKINVDCx6p67_ASAP7_75t_R g676 ( 
.A(n_457),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_464),
.B(n_513),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_569),
.B(n_508),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_661),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_556),
.A2(n_425),
.B1(n_415),
.B2(n_309),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_530),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_549),
.B(n_508),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_566),
.B(n_191),
.Y(n_683)
);

NAND2x1p5_ASAP7_75t_L g684 ( 
.A(n_664),
.B(n_212),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_531),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_538),
.A2(n_310),
.B1(n_307),
.B2(n_303),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_530),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_540),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_661),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_540),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_606),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_541),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_566),
.B(n_305),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_643),
.A2(n_285),
.B1(n_294),
.B2(n_303),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_584),
.B(n_527),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_606),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_547),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_584),
.B(n_308),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_531),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_599),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_658),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_599),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_559),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_541),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_534),
.B(n_646),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_579),
.B(n_508),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_671),
.A2(n_266),
.B1(n_208),
.B2(n_289),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_646),
.B(n_528),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_559),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_552),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_596),
.B(n_429),
.Y(n_713)
);

BUFx8_ASAP7_75t_L g714 ( 
.A(n_585),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_604),
.A2(n_319),
.B1(n_314),
.B2(n_315),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_561),
.B(n_231),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_544),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_589),
.B(n_508),
.Y(n_718)
);

O2A1O1Ixp5_ASAP7_75t_L g719 ( 
.A1(n_563),
.A2(n_508),
.B(n_232),
.C(n_289),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_599),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_563),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_567),
.Y(n_722)
);

NAND2x1_ASAP7_75t_L g723 ( 
.A(n_664),
.B(n_457),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_528),
.B(n_316),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_611),
.B(n_436),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_591),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_580),
.B(n_290),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_635),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_525),
.B(n_317),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_674),
.B(n_451),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_525),
.B(n_321),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_674),
.B(n_650),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_544),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_548),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_601),
.B(n_451),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_548),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_567),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_568),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_526),
.B(n_324),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_526),
.B(n_436),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_573),
.A2(n_327),
.B1(n_328),
.B2(n_338),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_568),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_585),
.B(n_444),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_629),
.B(n_346),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_536),
.B(n_451),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_628),
.B(n_349),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_536),
.B(n_454),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_565),
.A2(n_307),
.B1(n_294),
.B2(n_323),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_537),
.B(n_454),
.Y(n_749)
);

BUFx6f_ASAP7_75t_SL g750 ( 
.A(n_552),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_605),
.B(n_213),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_537),
.B(n_221),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_617),
.B(n_214),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_535),
.B(n_444),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_550),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_550),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_665),
.B(n_293),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_539),
.B(n_221),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_588),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_539),
.B(n_543),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_572),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_573),
.A2(n_269),
.B1(n_222),
.B2(n_225),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_573),
.B(n_216),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_558),
.B(n_464),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_533),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_573),
.B(n_224),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_575),
.B(n_211),
.Y(n_767)
);

HB1xp67_ASAP7_75t_SL g768 ( 
.A(n_570),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_620),
.B(n_301),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_552),
.Y(n_770)
);

INVx8_ASAP7_75t_L g771 ( 
.A(n_671),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_671),
.A2(n_222),
.B1(n_244),
.B2(n_269),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_543),
.B(n_225),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_581),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_597),
.Y(n_775)
);

NOR3xp33_ASAP7_75t_L g776 ( 
.A(n_640),
.B(n_236),
.C(n_229),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_581),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_533),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_588),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_602),
.B(n_227),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_545),
.B(n_229),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_618),
.B(n_301),
.Y(n_782)
);

INVx8_ASAP7_75t_L g783 ( 
.A(n_671),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_586),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_603),
.A2(n_284),
.B1(n_332),
.B2(n_236),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_593),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_603),
.A2(n_333),
.B1(n_326),
.B2(n_244),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_594),
.B(n_555),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_637),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_637),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_570),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_592),
.B(n_301),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_609),
.B(n_642),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_636),
.A2(n_513),
.B(n_464),
.C(n_478),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_545),
.B(n_284),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_546),
.B(n_326),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_546),
.B(n_332),
.Y(n_797)
);

BUFx5_ASAP7_75t_L g798 ( 
.A(n_614),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_542),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_658),
.B(n_301),
.Y(n_800)
);

BUFx5_ASAP7_75t_L g801 ( 
.A(n_614),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_565),
.A2(n_232),
.B(n_266),
.C(n_345),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_593),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_637),
.Y(n_804)
);

OAI22xp33_ASAP7_75t_L g805 ( 
.A1(n_634),
.A2(n_350),
.B1(n_339),
.B2(n_336),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_553),
.B(n_301),
.Y(n_806)
);

BUFx8_ASAP7_75t_L g807 ( 
.A(n_654),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_608),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_642),
.B(n_586),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_598),
.B(n_230),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_598),
.B(n_233),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_654),
.B(n_234),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_600),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_542),
.B(n_333),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_600),
.B(n_238),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_610),
.B(n_343),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_610),
.B(n_343),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_564),
.B(n_293),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_565),
.A2(n_583),
.B1(n_551),
.B2(n_663),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_608),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_558),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_612),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_565),
.B(n_345),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_607),
.B(n_330),
.C(n_339),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_583),
.B(n_448),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_583),
.B(n_301),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_612),
.Y(n_827)
);

OR2x6_ASAP7_75t_SL g828 ( 
.A(n_624),
.B(n_582),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_651),
.B(n_239),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_666),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_583),
.B(n_448),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_676),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_668),
.B(n_242),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_656),
.B(n_313),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_668),
.B(n_243),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_615),
.B(n_313),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_670),
.B(n_448),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_615),
.B(n_313),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_SL g839 ( 
.A(n_624),
.B(n_206),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_670),
.B(n_448),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_673),
.B(n_453),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_551),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_673),
.B(n_246),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_532),
.B(n_248),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_619),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_732),
.A2(n_660),
.B(n_638),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_754),
.B(n_582),
.Y(n_847)
);

OAI21xp33_ASAP7_75t_L g848 ( 
.A1(n_727),
.A2(n_716),
.B(n_683),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_760),
.A2(n_638),
.B(n_615),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_678),
.A2(n_638),
.B(n_657),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_682),
.A2(n_669),
.B(n_659),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_713),
.B(n_677),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_727),
.B(n_616),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_800),
.A2(n_622),
.B(n_529),
.Y(n_854)
);

BUFx4f_ASAP7_75t_L g855 ( 
.A(n_789),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_726),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_697),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_529),
.B(n_675),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_695),
.B(n_597),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_719),
.A2(n_621),
.B(n_616),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_793),
.A2(n_707),
.B1(n_695),
.B2(n_710),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_776),
.A2(n_625),
.B(n_627),
.C(n_623),
.Y(n_862)
);

AO21x1_ASAP7_75t_L g863 ( 
.A1(n_709),
.A2(n_672),
.B(n_623),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_743),
.B(n_413),
.Y(n_864)
);

AOI21xp33_ASAP7_75t_L g865 ( 
.A1(n_780),
.A2(n_577),
.B(n_595),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_718),
.A2(n_529),
.B(n_554),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_829),
.B(n_740),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_726),
.B(n_728),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_728),
.B(n_613),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_714),
.Y(n_870)
);

O2A1O1Ixp5_ASAP7_75t_L g871 ( 
.A1(n_834),
.A2(n_672),
.B(n_621),
.C(n_625),
.Y(n_871)
);

AND2x6_ASAP7_75t_L g872 ( 
.A(n_832),
.B(n_627),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_829),
.B(n_641),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_730),
.A2(n_529),
.B(n_554),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_679),
.B(n_641),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_686),
.A2(n_676),
.B1(n_667),
.B2(n_641),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_818),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_765),
.A2(n_529),
.B(n_560),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_719),
.A2(n_632),
.B(n_631),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_701),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_765),
.A2(n_562),
.B(n_560),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_765),
.A2(n_574),
.B(n_562),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_765),
.A2(n_578),
.B(n_574),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_685),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_691),
.B(n_414),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_809),
.A2(n_667),
.B(n_578),
.C(n_655),
.Y(n_886)
);

OAI321xp33_ASAP7_75t_L g887 ( 
.A1(n_686),
.A2(n_336),
.A3(n_350),
.B1(n_439),
.B2(n_414),
.C(n_418),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_707),
.B(n_667),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_793),
.A2(n_553),
.B1(n_590),
.B2(n_662),
.Y(n_889)
);

O2A1O1Ixp5_ASAP7_75t_L g890 ( 
.A1(n_769),
.A2(n_576),
.B(n_587),
.C(n_571),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_809),
.A2(n_745),
.B(n_747),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_757),
.B(n_312),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_704),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_821),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_689),
.B(n_844),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_821),
.Y(n_896)
);

NAND2x1_ASAP7_75t_L g897 ( 
.A(n_832),
.B(n_571),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_749),
.A2(n_632),
.B(n_631),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_696),
.B(n_418),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_714),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_844),
.B(n_639),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_639),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_776),
.A2(n_647),
.B(n_655),
.C(n_644),
.Y(n_903)
);

OAI321xp33_ASAP7_75t_L g904 ( 
.A1(n_805),
.A2(n_433),
.A3(n_442),
.B1(n_439),
.B2(n_437),
.C(n_419),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_711),
.B(n_644),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_701),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_721),
.B(n_647),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_778),
.A2(n_571),
.B(n_576),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_729),
.A2(n_662),
.B(n_649),
.C(n_652),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_752),
.A2(n_649),
.B(n_576),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_731),
.A2(n_739),
.B(n_724),
.C(n_782),
.Y(n_911)
);

BUFx4f_ASAP7_75t_L g912 ( 
.A(n_790),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_788),
.B(n_278),
.C(n_254),
.Y(n_913)
);

AO21x1_ASAP7_75t_L g914 ( 
.A1(n_684),
.A2(n_653),
.B(n_652),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_778),
.A2(n_587),
.B(n_648),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_778),
.A2(n_587),
.B(n_648),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_722),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_737),
.B(n_619),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_778),
.A2(n_653),
.B(n_645),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_812),
.B(n_274),
.C(n_262),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_819),
.A2(n_331),
.B1(n_311),
.B2(n_329),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_799),
.A2(n_645),
.B(n_633),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_738),
.B(n_626),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_791),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_680),
.B(n_263),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_742),
.B(n_626),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_758),
.A2(n_633),
.B(n_630),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_775),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_764),
.B(n_313),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_683),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_832),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_761),
.B(n_630),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_773),
.A2(n_590),
.B(n_553),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_781),
.A2(n_590),
.B(n_553),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_775),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_799),
.A2(n_453),
.B(n_313),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_702),
.A2(n_313),
.B1(n_341),
.B2(n_257),
.Y(n_937)
);

BUFx4f_ASAP7_75t_L g938 ( 
.A(n_804),
.Y(n_938)
);

NAND2x1_ASAP7_75t_L g939 ( 
.A(n_832),
.B(n_553),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_799),
.A2(n_453),
.B(n_341),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_699),
.B(n_419),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_774),
.B(n_553),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_751),
.A2(n_261),
.B(n_259),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_685),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_799),
.A2(n_453),
.B(n_341),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_735),
.A2(n_341),
.B(n_486),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_777),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_825),
.A2(n_341),
.B(n_486),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_723),
.A2(n_474),
.B(n_473),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_784),
.B(n_553),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_702),
.B(n_341),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_748),
.A2(n_249),
.B1(n_267),
.B2(n_268),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_831),
.A2(n_473),
.B(n_485),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_795),
.A2(n_590),
.B(n_480),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_813),
.B(n_590),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_823),
.A2(n_473),
.B(n_485),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_796),
.A2(n_488),
.B(n_513),
.C(n_482),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_839),
.B(n_265),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_685),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_700),
.B(n_478),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_830),
.B(n_590),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_700),
.A2(n_720),
.B(n_703),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_700),
.A2(n_473),
.B(n_511),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_842),
.B(n_420),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_836),
.A2(n_838),
.B(n_797),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_810),
.B(n_590),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_763),
.A2(n_459),
.B1(n_457),
.B2(n_480),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_700),
.A2(n_511),
.B(n_510),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_699),
.B(n_420),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_685),
.Y(n_970)
);

AOI33xp33_ASAP7_75t_L g971 ( 
.A1(n_694),
.A2(n_442),
.A3(n_437),
.B1(n_424),
.B2(n_433),
.B3(n_427),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_810),
.B(n_511),
.Y(n_972)
);

BUFx8_ASAP7_75t_L g973 ( 
.A(n_750),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_703),
.B(n_478),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_703),
.A2(n_511),
.B(n_510),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_842),
.B(n_424),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_766),
.B(n_276),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_751),
.A2(n_279),
.B(n_291),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_794),
.A2(n_459),
.B(n_480),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_753),
.B(n_295),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_811),
.B(n_474),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_681),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_703),
.A2(n_510),
.B(n_507),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_720),
.A2(n_510),
.B(n_507),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_837),
.A2(n_507),
.B(n_474),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_811),
.B(n_507),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_720),
.A2(n_493),
.B(n_485),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_687),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_720),
.B(n_482),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_815),
.B(n_833),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_840),
.A2(n_493),
.B(n_485),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_771),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_688),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_841),
.A2(n_494),
.B(n_486),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_794),
.A2(n_817),
.B(n_816),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_690),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_780),
.A2(n_482),
.B(n_503),
.C(n_488),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_806),
.A2(n_493),
.B(n_486),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_815),
.B(n_474),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_833),
.B(n_490),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_814),
.A2(n_490),
.B(n_493),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_835),
.B(n_490),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_684),
.A2(n_783),
.B1(n_771),
.B2(n_772),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_826),
.A2(n_494),
.B(n_490),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_692),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_712),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_835),
.B(n_494),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_753),
.B(n_299),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_771),
.A2(n_306),
.B1(n_354),
.B2(n_353),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_783),
.A2(n_337),
.B1(n_352),
.B2(n_355),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_706),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_725),
.B(n_427),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_SL g1013 ( 
.A1(n_802),
.A2(n_503),
.B(n_498),
.C(n_495),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_717),
.A2(n_494),
.B(n_499),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_733),
.A2(n_501),
.B(n_499),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_694),
.A2(n_431),
.B(n_503),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_767),
.A2(n_495),
.B(n_488),
.C(n_492),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_734),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_783),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_736),
.A2(n_756),
.B(n_755),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_843),
.B(n_501),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_748),
.A2(n_431),
.B1(n_498),
.B2(n_495),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_843),
.B(n_501),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_693),
.A2(n_501),
.B(n_499),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_698),
.A2(n_499),
.B(n_498),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_741),
.B(n_492),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_805),
.A2(n_492),
.B(n_312),
.C(n_20),
.Y(n_1027)
);

AO21x1_ASAP7_75t_L g1028 ( 
.A1(n_762),
.A2(n_17),
.B(n_19),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_798),
.B(n_506),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_750),
.B(n_312),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_798),
.B(n_506),
.Y(n_1031)
);

BUFx4f_ASAP7_75t_L g1032 ( 
.A(n_768),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_792),
.A2(n_20),
.B(n_21),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_798),
.B(n_506),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_807),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_857),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_990),
.A2(n_715),
.B1(n_744),
.B2(n_787),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_848),
.B(n_768),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_867),
.B(n_770),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_930),
.B(n_746),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_980),
.A2(n_824),
.B(n_785),
.C(n_827),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_SL g1042 ( 
.A(n_931),
.B(n_845),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_849),
.A2(n_850),
.B(n_873),
.Y(n_1043)
);

OAI22x1_ASAP7_75t_L g1044 ( 
.A1(n_925),
.A2(n_824),
.B1(n_828),
.B2(n_807),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_SL g1045 ( 
.A(n_992),
.B(n_822),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_895),
.B(n_798),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_877),
.B(n_312),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_877),
.B(n_820),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_1008),
.B(n_801),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_861),
.B(n_853),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_868),
.B(n_801),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_894),
.B(n_808),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_893),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_865),
.A2(n_803),
.B(n_786),
.C(n_779),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_921),
.B(n_856),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_977),
.A2(n_759),
.B(n_26),
.C(n_27),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_892),
.B(n_506),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_SL g1058 ( 
.A(n_896),
.B(n_801),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_917),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_924),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_869),
.B(n_801),
.Y(n_1061)
);

AO21x1_ASAP7_75t_L g1062 ( 
.A1(n_911),
.A2(n_801),
.B(n_798),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_931),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_947),
.B(n_801),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_851),
.A2(n_798),
.B(n_506),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_901),
.A2(n_506),
.B1(n_94),
.B2(n_96),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_852),
.A2(n_21),
.B(n_30),
.C(n_33),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_SL g1068 ( 
.A(n_992),
.B(n_506),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1019),
.B(n_97),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_931),
.B(n_506),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_966),
.A2(n_92),
.B1(n_178),
.B2(n_177),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_988),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_846),
.A2(n_480),
.B(n_459),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_858),
.A2(n_480),
.B(n_459),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_1006),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_931),
.A2(n_480),
.B(n_459),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1029),
.A2(n_480),
.B(n_459),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_891),
.B(n_480),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_988),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_958),
.B(n_33),
.C(n_34),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_884),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1031),
.A2(n_480),
.B(n_459),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_891),
.A2(n_103),
.B1(n_172),
.B2(n_170),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1034),
.A2(n_459),
.B(n_457),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_864),
.B(n_36),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_885),
.B(n_480),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_884),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_972),
.A2(n_457),
.B(n_459),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_847),
.B(n_83),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1019),
.B(n_86),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_981),
.A2(n_999),
.B(n_986),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_884),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1000),
.A2(n_80),
.B1(n_167),
.B2(n_153),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_941),
.B(n_79),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_970),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_899),
.B(n_459),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_976),
.B(n_39),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1002),
.A2(n_1021),
.B(n_1007),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_964),
.B(n_39),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_970),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_875),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_1032),
.B(n_74),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1023),
.A2(n_457),
.B(n_109),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1012),
.B(n_457),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_993),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_L g1106 ( 
.A1(n_995),
.A2(n_863),
.B(n_914),
.C(n_997),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_970),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1028),
.A2(n_457),
.B1(n_43),
.B2(n_44),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_910),
.A2(n_457),
.B(n_114),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_910),
.A2(n_149),
.B(n_146),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_976),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_R g1112 ( 
.A(n_1032),
.B(n_144),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1011),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_996),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1012),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_943),
.B(n_42),
.Y(n_1116)
);

BUFx4f_ASAP7_75t_L g1117 ( 
.A(n_870),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_918),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_L g1119 ( 
.A1(n_995),
.A2(n_141),
.B(n_138),
.C(n_127),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_923),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_L g1121 ( 
.A(n_944),
.B(n_126),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_941),
.B(n_44),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_854),
.A2(n_119),
.B(n_46),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_969),
.B(n_913),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_969),
.B(n_45),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_920),
.B(n_45),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_L g1127 ( 
.A(n_978),
.B(n_49),
.C(n_56),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1026),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_926),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_944),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1027),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_962),
.A2(n_58),
.B(n_60),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1003),
.A2(n_61),
.B1(n_876),
.B2(n_889),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_886),
.A2(n_61),
.B(n_952),
.C(n_859),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_866),
.A2(n_888),
.B(n_878),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1033),
.A2(n_1016),
.B1(n_952),
.B2(n_1022),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_985),
.A2(n_881),
.B(n_882),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_959),
.B(n_880),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_855),
.B(n_912),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_959),
.B(n_906),
.Y(n_1140)
);

AO21x1_ASAP7_75t_L g1141 ( 
.A1(n_929),
.A2(n_951),
.B(n_903),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_898),
.A2(n_908),
.B(n_874),
.Y(n_1142)
);

CKINVDCx10_ASAP7_75t_R g1143 ( 
.A(n_1035),
.Y(n_1143)
);

AND2x2_ASAP7_75t_SL g1144 ( 
.A(n_1030),
.B(n_855),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_898),
.A2(n_883),
.B(n_933),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_933),
.A2(n_934),
.B(n_916),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_928),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_912),
.B(n_938),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_932),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_934),
.A2(n_915),
.B(n_960),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_SL g1151 ( 
.A(n_1030),
.B(n_971),
.C(n_957),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_935),
.A2(n_907),
.B1(n_905),
.B2(n_902),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_900),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_974),
.A2(n_989),
.B(n_939),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_938),
.B(n_1009),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_982),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_942),
.A2(n_950),
.B1(n_955),
.B2(n_961),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_887),
.B(n_904),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_897),
.A2(n_922),
.B(n_919),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_879),
.A2(n_954),
.B(n_860),
.C(n_979),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1010),
.B(n_1018),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_973),
.B(n_996),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1005),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_871),
.A2(n_862),
.B(n_860),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1005),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_R g1166 ( 
.A(n_973),
.B(n_872),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_937),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1017),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_887),
.B(n_904),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_909),
.B(n_1025),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_872),
.B(n_1022),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_965),
.B(n_927),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1020),
.Y(n_1173)
);

OAI21xp33_ASAP7_75t_SL g1174 ( 
.A1(n_954),
.A2(n_879),
.B(n_979),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_953),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_872),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_890),
.A2(n_927),
.B(n_975),
.Y(n_1177)
);

O2A1O1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1013),
.A2(n_948),
.B(n_1024),
.C(n_946),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_963),
.A2(n_984),
.B(n_987),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_SL g1180 ( 
.A1(n_967),
.A2(n_872),
.B1(n_949),
.B2(n_1001),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_936),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_940),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_968),
.B(n_983),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_956),
.B(n_991),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_994),
.A2(n_998),
.B(n_945),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1004),
.B(n_1014),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1015),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_867),
.B(n_990),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_849),
.A2(n_674),
.B(n_664),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_R g1190 ( 
.A(n_894),
.B(n_558),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_931),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_931),
.Y(n_1192)
);

NAND4xp25_ASAP7_75t_L g1193 ( 
.A(n_1055),
.B(n_1099),
.C(n_1116),
.D(n_1111),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1038),
.B(n_1055),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_1037),
.A2(n_1061),
.B(n_1116),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1085),
.B(n_1047),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1049),
.A2(n_1040),
.B(n_1134),
.C(n_1128),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1127),
.A2(n_1188),
.B1(n_1099),
.B2(n_1128),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1049),
.A2(n_1189),
.B(n_1142),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1065),
.A2(n_1050),
.B(n_1145),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1106),
.A2(n_1164),
.B(n_1172),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1172),
.A2(n_1062),
.A3(n_1177),
.B(n_1141),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1051),
.A2(n_1046),
.B1(n_1040),
.B2(n_1136),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1036),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1051),
.A2(n_1041),
.B(n_1110),
.C(n_1174),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1106),
.A2(n_1146),
.B(n_1119),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1048),
.B(n_1097),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1185),
.A2(n_1179),
.B(n_1150),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1124),
.A2(n_1127),
.B(n_1133),
.C(n_1056),
.Y(n_1211)
);

AOI221x1_ASAP7_75t_L g1212 ( 
.A1(n_1083),
.A2(n_1109),
.B1(n_1066),
.B2(n_1080),
.C(n_1123),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1160),
.A2(n_1170),
.B(n_1152),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1053),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1118),
.B(n_1120),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1108),
.A2(n_1131),
.B(n_1136),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1063),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1063),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1126),
.A2(n_1039),
.B(n_1125),
.C(n_1067),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1115),
.B(n_1139),
.Y(n_1220)
);

AO32x2_ASAP7_75t_L g1221 ( 
.A1(n_1180),
.A2(n_1157),
.A3(n_1071),
.B1(n_1093),
.B2(n_1092),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1075),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1183),
.A2(n_1173),
.B(n_1184),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1060),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1178),
.A2(n_1175),
.B(n_1154),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1148),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1129),
.B(n_1149),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1144),
.B(n_1058),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1119),
.A2(n_1168),
.B(n_1171),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1054),
.A2(n_1073),
.B(n_1186),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1155),
.A2(n_1158),
.B1(n_1169),
.B2(n_1059),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1147),
.B(n_1156),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1064),
.A2(n_1057),
.B(n_1068),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1078),
.A2(n_1045),
.B(n_1101),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1167),
.A2(n_1161),
.B(n_1151),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_1089),
.B(n_1103),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1144),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1122),
.A2(n_1151),
.B(n_1094),
.C(n_1132),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1063),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1074),
.A2(n_1088),
.A3(n_1084),
.B(n_1082),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1077),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1107),
.Y(n_1242)
);

INVx8_ASAP7_75t_L g1243 ( 
.A(n_1063),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1070),
.A2(n_1121),
.B(n_1105),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1113),
.A2(n_1076),
.B(n_1081),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1107),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1108),
.A2(n_1044),
.B1(n_1153),
.B2(n_1156),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1191),
.A2(n_1192),
.B(n_1182),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1191),
.A2(n_1192),
.B(n_1181),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1072),
.B(n_1114),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1079),
.B(n_1052),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1163),
.A2(n_1165),
.A3(n_1104),
.B(n_1130),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1069),
.A2(n_1090),
.B1(n_1086),
.B2(n_1096),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1191),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1176),
.A2(n_1090),
.B(n_1069),
.C(n_1190),
.Y(n_1255)
);

AOI221xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1176),
.A2(n_1087),
.B1(n_1095),
.B2(n_1100),
.C(n_1192),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1191),
.A2(n_1192),
.B(n_1042),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1087),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1087),
.A2(n_1095),
.B(n_1100),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1087),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1095),
.Y(n_1261)
);

AOI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1117),
.A2(n_1092),
.B(n_1095),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1100),
.A2(n_1117),
.B1(n_1112),
.B2(n_1102),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1100),
.A2(n_1166),
.B(n_1162),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1143),
.B(n_848),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1063),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1050),
.A2(n_990),
.B(n_848),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1116),
.A2(n_848),
.B1(n_990),
.B2(n_980),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1038),
.B(n_848),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1188),
.B(n_864),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1145),
.A2(n_1177),
.B(n_1065),
.Y(n_1275)
);

OAI211xp5_ASAP7_75t_L g1276 ( 
.A1(n_1055),
.A2(n_848),
.B(n_594),
.C(n_925),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1036),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1188),
.B(n_848),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1188),
.B(n_848),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1172),
.A2(n_1062),
.A3(n_914),
.B(n_1177),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1049),
.A2(n_848),
.B(n_990),
.C(n_980),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1188),
.B(n_864),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1063),
.B(n_931),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1049),
.A2(n_848),
.B(n_990),
.C(n_980),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1049),
.A2(n_848),
.B(n_990),
.C(n_980),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1128),
.B(n_861),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1060),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1172),
.A2(n_1062),
.A3(n_914),
.B(n_1177),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1036),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1050),
.A2(n_990),
.B(n_848),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1036),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_1038),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_864),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1075),
.Y(n_1299)
);

AO21x1_ASAP7_75t_L g1300 ( 
.A1(n_1049),
.A2(n_990),
.B(n_1133),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1036),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1075),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1128),
.B(n_861),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1188),
.A2(n_848),
.B(n_1008),
.C(n_980),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1063),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1060),
.Y(n_1311)
);

AOI31xp67_ASAP7_75t_L g1312 ( 
.A1(n_1170),
.A2(n_1184),
.A3(n_1188),
.B(n_1050),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1190),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1036),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1049),
.A2(n_848),
.B(n_990),
.C(n_980),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1188),
.B(n_848),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1036),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1036),
.Y(n_1318)
);

O2A1O1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1188),
.A2(n_848),
.B(n_1008),
.C(n_980),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1188),
.B(n_848),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_SL g1322 ( 
.A(n_1144),
.B(n_1032),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1188),
.B(n_848),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1060),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1049),
.A2(n_848),
.B(n_990),
.C(n_980),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1172),
.A2(n_1062),
.A3(n_914),
.B(n_1177),
.Y(n_1326)
);

INVx5_ASAP7_75t_L g1327 ( 
.A(n_1063),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1172),
.A2(n_1062),
.A3(n_914),
.B(n_1177),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1036),
.Y(n_1329)
);

OAI22x1_ASAP7_75t_L g1330 ( 
.A1(n_1055),
.A2(n_925),
.B1(n_788),
.B2(n_1116),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1049),
.A2(n_848),
.B(n_990),
.C(n_980),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1116),
.A2(n_848),
.B1(n_1008),
.B2(n_980),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1036),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1060),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1060),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1036),
.Y(n_1338)
);

AOI31xp67_ASAP7_75t_L g1339 ( 
.A1(n_1170),
.A2(n_1184),
.A3(n_1188),
.B(n_1050),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_1159),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1188),
.B(n_848),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1172),
.A2(n_1062),
.A3(n_914),
.B(n_1177),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1091),
.A2(n_1098),
.B(n_1043),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1188),
.A2(n_848),
.B(n_1008),
.C(n_980),
.Y(n_1345)
);

OAI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1271),
.A2(n_1193),
.B1(n_1228),
.B2(n_1216),
.Y(n_1346)
);

BUFx8_ASAP7_75t_L g1347 ( 
.A(n_1324),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1311),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1332),
.A2(n_1194),
.B1(n_1271),
.B2(n_1272),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1276),
.A2(n_1216),
.B(n_1193),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1330),
.A2(n_1195),
.B1(n_1270),
.B2(n_1294),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1247),
.A2(n_1300),
.B1(n_1199),
.B2(n_1288),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1243),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1247),
.A2(n_1199),
.B1(n_1304),
.B2(n_1288),
.Y(n_1354)
);

BUFx8_ASAP7_75t_L g1355 ( 
.A(n_1222),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1304),
.A2(n_1205),
.B1(n_1235),
.B2(n_1341),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1313),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1224),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1299),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1279),
.A2(n_1321),
.B1(n_1323),
.B2(n_1316),
.Y(n_1360)
);

BUFx8_ASAP7_75t_SL g1361 ( 
.A(n_1265),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1224),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1303),
.Y(n_1363)
);

BUFx12f_ASAP7_75t_L g1364 ( 
.A(n_1226),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1336),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1215),
.B(n_1227),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1280),
.A2(n_1274),
.B1(n_1284),
.B2(n_1298),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1214),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1243),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1296),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1327),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1253),
.A2(n_1325),
.B1(n_1283),
.B2(n_1286),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1228),
.A2(n_1231),
.B1(n_1322),
.B2(n_1197),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1327),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1209),
.B(n_1232),
.Y(n_1375)
);

INVx6_ASAP7_75t_L g1376 ( 
.A(n_1327),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1226),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1322),
.A2(n_1237),
.B1(n_1296),
.B2(n_1203),
.Y(n_1378)
);

BUFx4f_ASAP7_75t_SL g1379 ( 
.A(n_1220),
.Y(n_1379)
);

CKINVDCx6p67_ASAP7_75t_R g1380 ( 
.A(n_1243),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1290),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1237),
.A2(n_1203),
.B1(n_1338),
.B2(n_1278),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_1254),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1254),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1293),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1254),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1295),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1301),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_SL g1389 ( 
.A(n_1260),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1309),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_1263),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1314),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1246),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1309),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1317),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1251),
.A2(n_1236),
.B1(n_1318),
.B2(n_1329),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1253),
.A2(n_1287),
.B1(n_1315),
.B2(n_1331),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1260),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_L g1399 ( 
.A(n_1285),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1260),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1335),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1242),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1213),
.A2(n_1208),
.B1(n_1229),
.B2(n_1202),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1250),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1259),
.B(n_1248),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1258),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1312),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1337),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1262),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1252),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1217),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1339),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1261),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1212),
.A2(n_1264),
.B1(n_1249),
.B2(n_1208),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1217),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1211),
.B(n_1198),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1308),
.A2(n_1345),
.B1(n_1319),
.B2(n_1229),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1218),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1255),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1252),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1218),
.A2(n_1239),
.B1(n_1268),
.B2(n_1257),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1252),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1201),
.A2(n_1234),
.B1(n_1223),
.B2(n_1233),
.Y(n_1423)
);

INVx6_ASAP7_75t_L g1424 ( 
.A(n_1239),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1268),
.Y(n_1425)
);

BUFx8_ASAP7_75t_L g1426 ( 
.A(n_1221),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1219),
.A2(n_1238),
.B(n_1207),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1245),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1240),
.Y(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1256),
.Y(n_1430)
);

BUFx2_ASAP7_75t_SL g1431 ( 
.A(n_1196),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1267),
.A2(n_1289),
.B1(n_1343),
.B2(n_1334),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1282),
.A2(n_1344),
.B1(n_1291),
.B2(n_1333),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1240),
.Y(n_1434)
);

BUFx8_ASAP7_75t_SL g1435 ( 
.A(n_1275),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1244),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1302),
.A2(n_1320),
.B1(n_1307),
.B2(n_1305),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1241),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1306),
.Y(n_1439)
);

CKINVDCx11_ASAP7_75t_R g1440 ( 
.A(n_1256),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1221),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1240),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1225),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1221),
.A2(n_1230),
.B1(n_1210),
.B2(n_1277),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1200),
.A2(n_1273),
.B1(n_1266),
.B2(n_1269),
.Y(n_1445)
);

CKINVDCx6p67_ASAP7_75t_R g1446 ( 
.A(n_1281),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1281),
.Y(n_1447)
);

BUFx12f_ASAP7_75t_L g1448 ( 
.A(n_1292),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1204),
.B(n_1292),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1297),
.A2(n_1310),
.B1(n_1340),
.B2(n_1204),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1204),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1326),
.A2(n_1271),
.B1(n_990),
.B2(n_1193),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1342),
.B(n_1326),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1328),
.A2(n_1276),
.B1(n_1194),
.B2(n_925),
.Y(n_1454)
);

INVx8_ASAP7_75t_L g1455 ( 
.A(n_1342),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1342),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1332),
.A2(n_848),
.B1(n_1330),
.B2(n_1194),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1324),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1209),
.B(n_1197),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1276),
.A2(n_1194),
.B1(n_925),
.B2(n_604),
.Y(n_1460)
);

BUFx8_ASAP7_75t_L g1461 ( 
.A(n_1324),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1243),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1332),
.A2(n_1194),
.B1(n_1271),
.B2(n_990),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1324),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1332),
.A2(n_1194),
.B1(n_1271),
.B2(n_990),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1222),
.Y(n_1466)
);

INVx6_ASAP7_75t_L g1467 ( 
.A(n_1327),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1327),
.Y(n_1468)
);

BUFx2_ASAP7_75t_SL g1469 ( 
.A(n_1313),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1194),
.A2(n_1330),
.B1(n_980),
.B2(n_1008),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1332),
.A2(n_848),
.B1(n_1330),
.B2(n_1194),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1332),
.A2(n_1194),
.B1(n_1271),
.B2(n_990),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1206),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1196),
.A2(n_1282),
.B(n_1267),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1324),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1222),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1327),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1332),
.A2(n_848),
.B1(n_1330),
.B2(n_1194),
.Y(n_1478)
);

BUFx10_ASAP7_75t_L g1479 ( 
.A(n_1222),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1410),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1420),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1393),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1453),
.B(n_1449),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1422),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1447),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1441),
.B(n_1416),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1445),
.A2(n_1450),
.B(n_1432),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1442),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1429),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1439),
.B(n_1436),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1460),
.A2(n_1349),
.B1(n_1463),
.B2(n_1465),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1351),
.B(n_1368),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1438),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1448),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1456),
.B(n_1434),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1427),
.A2(n_1354),
.B(n_1350),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1387),
.B(n_1392),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1351),
.B(n_1387),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1402),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1435),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1348),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1445),
.A2(n_1450),
.B(n_1403),
.Y(n_1502)
);

AOI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1443),
.A2(n_1428),
.B(n_1407),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1395),
.B(n_1356),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1403),
.A2(n_1437),
.B(n_1412),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1446),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1448),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1356),
.B(n_1451),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1455),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1431),
.B(n_1372),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1430),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1459),
.B(n_1375),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1357),
.Y(n_1513)
);

NAND2x1_ASAP7_75t_L g1514 ( 
.A(n_1423),
.B(n_1438),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1397),
.B(n_1405),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1382),
.B(n_1367),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1382),
.B(n_1367),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1385),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1433),
.A2(n_1414),
.B(n_1452),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1388),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1426),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1413),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1401),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1366),
.B(n_1360),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1381),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1472),
.A2(n_1454),
.B1(n_1346),
.B2(n_1478),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1358),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1437),
.A2(n_1423),
.B(n_1474),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1473),
.B(n_1360),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1470),
.B(n_1457),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1430),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1362),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1430),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1430),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1474),
.Y(n_1535)
);

INVx4_ASAP7_75t_SL g1536 ( 
.A(n_1374),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1474),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1426),
.Y(n_1538)
);

AO21x1_ASAP7_75t_SL g1539 ( 
.A1(n_1352),
.A2(n_1373),
.B(n_1354),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1457),
.A2(n_1478),
.B1(n_1471),
.B2(n_1409),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1425),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1433),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1471),
.A2(n_1417),
.B(n_1396),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1404),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1374),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1414),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1418),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1444),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1452),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1374),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1440),
.Y(n_1551)
);

AO21x1_ASAP7_75t_SL g1552 ( 
.A1(n_1378),
.A2(n_1346),
.B(n_1419),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1347),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1406),
.B(n_1421),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1347),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1365),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1379),
.A2(n_1391),
.B1(n_1370),
.B2(n_1458),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1415),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1458),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1411),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1491),
.A2(n_1408),
.B(n_1399),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1486),
.A2(n_1379),
.B1(n_1464),
.B2(n_1475),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1483),
.B(n_1475),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1490),
.B(n_1377),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1490),
.B(n_1363),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1507),
.B(n_1390),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_SL g1567 ( 
.A1(n_1540),
.A2(n_1466),
.B(n_1462),
.C(n_1371),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1536),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1483),
.B(n_1469),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1492),
.B(n_1390),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1530),
.B(n_1364),
.Y(n_1571)
);

AOI211xp5_ASAP7_75t_L g1572 ( 
.A1(n_1543),
.A2(n_1369),
.B(n_1468),
.C(n_1477),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_SL g1573 ( 
.A1(n_1551),
.A2(n_1524),
.B(n_1513),
.C(n_1558),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1510),
.B(n_1467),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1510),
.A2(n_1514),
.B(n_1519),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1492),
.B(n_1477),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1526),
.A2(n_1399),
.B(n_1369),
.C(n_1468),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1502),
.A2(n_1398),
.B(n_1376),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1512),
.B(n_1361),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1525),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1497),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1487),
.A2(n_1462),
.B(n_1376),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1490),
.B(n_1384),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_SL g1584 ( 
.A(n_1510),
.B(n_1477),
.Y(n_1584)
);

NAND4xp25_ASAP7_75t_L g1585 ( 
.A(n_1546),
.B(n_1461),
.C(n_1476),
.D(n_1359),
.Y(n_1585)
);

CKINVDCx11_ASAP7_75t_R g1586 ( 
.A(n_1527),
.Y(n_1586)
);

AO21x2_ASAP7_75t_L g1587 ( 
.A1(n_1535),
.A2(n_1467),
.B(n_1398),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1559),
.B(n_1400),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1502),
.A2(n_1424),
.B(n_1383),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1498),
.B(n_1477),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1551),
.A2(n_1364),
.B1(n_1461),
.B2(n_1359),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1522),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1480),
.Y(n_1593)
);

OR2x6_ASAP7_75t_L g1594 ( 
.A(n_1510),
.B(n_1476),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1559),
.Y(n_1595)
);

OAI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1549),
.A2(n_1353),
.B(n_1479),
.Y(n_1596)
);

OAI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1549),
.A2(n_1386),
.B1(n_1353),
.B2(n_1355),
.C(n_1479),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1516),
.B(n_1380),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1546),
.A2(n_1353),
.B(n_1394),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1486),
.A2(n_1353),
.B(n_1389),
.C(n_1355),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1553),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1551),
.A2(n_1386),
.B(n_1508),
.C(n_1500),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1528),
.A2(n_1537),
.B(n_1542),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1496),
.A2(n_1386),
.B(n_1499),
.C(n_1501),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1521),
.A2(n_1538),
.B1(n_1508),
.B2(n_1500),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1514),
.A2(n_1519),
.B(n_1528),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1500),
.A2(n_1515),
.B1(n_1557),
.B2(n_1504),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1518),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1515),
.A2(n_1504),
.B1(n_1554),
.B2(n_1494),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1542),
.A2(n_1516),
.B(n_1517),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1547),
.B(n_1538),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1509),
.B(n_1506),
.Y(n_1613)
);

OA21x2_ASAP7_75t_L g1614 ( 
.A1(n_1537),
.A2(n_1531),
.B(n_1533),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1517),
.A2(n_1515),
.B(n_1498),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1520),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1533),
.A2(n_1534),
.B(n_1503),
.Y(n_1617)
);

AOI211xp5_ASAP7_75t_L g1618 ( 
.A1(n_1554),
.A2(n_1548),
.B(n_1506),
.C(n_1556),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1529),
.B(n_1544),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1560),
.Y(n_1620)
);

AO21x1_ASAP7_75t_L g1621 ( 
.A1(n_1558),
.A2(n_1534),
.B(n_1523),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1515),
.B(n_1511),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1603),
.B(n_1519),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1619),
.B(n_1480),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1614),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1578),
.B(n_1505),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1614),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1578),
.B(n_1505),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1589),
.B(n_1505),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1619),
.B(n_1548),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1609),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1607),
.B(n_1481),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1581),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1615),
.B(n_1489),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1616),
.B(n_1575),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1615),
.B(n_1489),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1622),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1561),
.A2(n_1496),
.B1(n_1539),
.B2(n_1552),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1587),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1572),
.A2(n_1515),
.B1(n_1482),
.B2(n_1539),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1616),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1611),
.B(n_1484),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1598),
.B(n_1485),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1621),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1587),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1582),
.B(n_1493),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1592),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1484),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1622),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1570),
.B(n_1495),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1626),
.B(n_1620),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1606),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1570),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1645),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1651),
.B(n_1488),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1642),
.A2(n_1552),
.B1(n_1561),
.B2(n_1594),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1650),
.B(n_1574),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1632),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1650),
.B(n_1612),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

INVx5_ASAP7_75t_SL g1665 ( 
.A(n_1649),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1626),
.B(n_1610),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

AOI21xp33_ASAP7_75t_L g1668 ( 
.A1(n_1647),
.A2(n_1604),
.B(n_1618),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1650),
.B(n_1595),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1630),
.B(n_1563),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

INVx5_ASAP7_75t_L g1674 ( 
.A(n_1641),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1627),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1630),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1634),
.B(n_1565),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1625),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1640),
.A2(n_1642),
.B1(n_1608),
.B2(n_1562),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1630),
.B(n_1576),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1625),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1630),
.B(n_1576),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1647),
.A2(n_1605),
.B1(n_1584),
.B2(n_1562),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1634),
.B(n_1636),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1646),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1590),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1646),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1639),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1647),
.A2(n_1574),
.B(n_1567),
.Y(n_1689)
);

OA332x1_ASAP7_75t_L g1690 ( 
.A1(n_1637),
.A2(n_1605),
.A3(n_1571),
.B1(n_1586),
.B2(n_1585),
.B3(n_1573),
.C1(n_1602),
.C2(n_1604),
.Y(n_1690)
);

AO21x2_ASAP7_75t_L g1691 ( 
.A1(n_1646),
.A2(n_1596),
.B(n_1599),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1627),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1634),
.B(n_1613),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1685),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1684),
.B(n_1626),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1671),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1684),
.B(n_1628),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1676),
.B(n_1637),
.Y(n_1698)
);

NAND2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1674),
.B(n_1648),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1643),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1665),
.B(n_1655),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1678),
.B(n_1637),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1678),
.B(n_1637),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1665),
.B(n_1628),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1665),
.B(n_1655),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1671),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1665),
.B(n_1628),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1655),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1662),
.B(n_1643),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1662),
.B(n_1624),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1681),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1685),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1666),
.B(n_1628),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1681),
.B(n_1633),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1666),
.B(n_1629),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1687),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1666),
.B(n_1629),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1656),
.B(n_1629),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1664),
.B(n_1624),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1687),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1656),
.B(n_1663),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1664),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1669),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1674),
.B(n_1641),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1674),
.B(n_1641),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1675),
.B(n_1633),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1656),
.B(n_1663),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1688),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1669),
.Y(n_1730)
);

AND2x4_ASAP7_75t_SL g1731 ( 
.A(n_1661),
.B(n_1594),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1667),
.B(n_1644),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1675),
.B(n_1629),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1723),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1729),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1729),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1723),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_R g1738 ( 
.A(n_1701),
.B(n_1658),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1731),
.A2(n_1660),
.B1(n_1683),
.B2(n_1668),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1711),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1729),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1698),
.B(n_1680),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_R g1743 ( 
.A(n_1729),
.B(n_1527),
.Y(n_1743)
);

NAND2x1_ASAP7_75t_L g1744 ( 
.A(n_1725),
.B(n_1661),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1724),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1722),
.B(n_1693),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1668),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1698),
.B(n_1680),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

OAI322xp33_ASAP7_75t_L g1750 ( 
.A1(n_1698),
.A2(n_1657),
.A3(n_1679),
.B1(n_1652),
.B2(n_1682),
.C1(n_1672),
.C2(n_1659),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1722),
.B(n_1693),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1730),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1709),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1731),
.B(n_1683),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1709),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1694),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_SL g1757 ( 
.A(n_1730),
.B(n_1532),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1694),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1702),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1699),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1696),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1712),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1712),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1732),
.B(n_1682),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1701),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1696),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1731),
.B(n_1532),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1702),
.B(n_1672),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1717),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1702),
.B(n_1686),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1717),
.Y(n_1771)
);

AOI222xp33_ASAP7_75t_L g1772 ( 
.A1(n_1731),
.A2(n_1640),
.B1(n_1623),
.B2(n_1644),
.C1(n_1636),
.C2(n_1638),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1722),
.B(n_1688),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1710),
.B(n_1657),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1688),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1728),
.B(n_1677),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1750),
.A2(n_1754),
.B1(n_1739),
.B2(n_1747),
.C(n_1736),
.Y(n_1777)
);

NOR2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1744),
.B(n_1553),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1763),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1735),
.B(n_1728),
.Y(n_1780)
);

NOR2x1p5_ASAP7_75t_SL g1781 ( 
.A(n_1761),
.B(n_1696),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1734),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1741),
.B(n_1553),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1737),
.Y(n_1784)
);

AND2x4_ASAP7_75t_SL g1785 ( 
.A(n_1741),
.B(n_1583),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1757),
.B(n_1679),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1701),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1767),
.B(n_1555),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1738),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1756),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1758),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1773),
.B(n_1705),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1752),
.B(n_1686),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1745),
.B(n_1710),
.Y(n_1794)
);

AND3x1_ASAP7_75t_L g1795 ( 
.A(n_1765),
.B(n_1591),
.C(n_1600),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1765),
.B(n_1705),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1746),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1773),
.B(n_1705),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1762),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1754),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1775),
.B(n_1708),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1775),
.B(n_1708),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1774),
.B(n_1720),
.Y(n_1803)
);

NAND4xp25_ASAP7_75t_L g1804 ( 
.A(n_1772),
.B(n_1571),
.C(n_1689),
.D(n_1585),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1740),
.B(n_1720),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1769),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1776),
.B(n_1708),
.Y(n_1807)
);

OAI211xp5_ASAP7_75t_L g1808 ( 
.A1(n_1743),
.A2(n_1744),
.B(n_1749),
.C(n_1689),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_SL g1809 ( 
.A1(n_1771),
.A2(n_1555),
.B(n_1577),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1776),
.B(n_1753),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1755),
.B(n_1715),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1760),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1777),
.A2(n_1760),
.B(n_1699),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1800),
.B(n_1779),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1789),
.B(n_1746),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1796),
.Y(n_1816)
);

OAI22x1_ASAP7_75t_L g1817 ( 
.A1(n_1786),
.A2(n_1760),
.B1(n_1699),
.B2(n_1601),
.Y(n_1817)
);

AOI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1808),
.A2(n_1759),
.B1(n_1768),
.B2(n_1742),
.C(n_1748),
.Y(n_1818)
);

OAI31xp33_ASAP7_75t_L g1819 ( 
.A1(n_1786),
.A2(n_1699),
.A3(n_1690),
.B(n_1704),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1795),
.A2(n_1691),
.B1(n_1704),
.B2(n_1707),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1785),
.B(n_1751),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1783),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1804),
.A2(n_1785),
.B1(n_1780),
.B2(n_1788),
.Y(n_1823)
);

INVxp33_ASAP7_75t_L g1824 ( 
.A(n_1788),
.Y(n_1824)
);

OAI21xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1778),
.A2(n_1801),
.B(n_1798),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1782),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1784),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1790),
.Y(n_1828)
);

AOI21xp33_ASAP7_75t_L g1829 ( 
.A1(n_1787),
.A2(n_1759),
.B(n_1768),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1798),
.B(n_1751),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1791),
.Y(n_1831)
);

OAI32xp33_ASAP7_75t_L g1832 ( 
.A1(n_1794),
.A2(n_1770),
.A3(n_1703),
.B1(n_1742),
.B2(n_1748),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_SL g1833 ( 
.A(n_1787),
.B(n_1568),
.Y(n_1833)
);

AOI322xp5_ASAP7_75t_L g1834 ( 
.A1(n_1797),
.A2(n_1718),
.A3(n_1715),
.B1(n_1713),
.B2(n_1719),
.C1(n_1695),
.C2(n_1697),
.Y(n_1834)
);

AOI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1787),
.A2(n_1770),
.B(n_1764),
.Y(n_1835)
);

OAI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1810),
.A2(n_1764),
.B(n_1645),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1801),
.A2(n_1691),
.B1(n_1707),
.B2(n_1704),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1799),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1816),
.Y(n_1839)
);

AOI21xp33_ASAP7_75t_L g1840 ( 
.A1(n_1824),
.A2(n_1812),
.B(n_1806),
.Y(n_1840)
);

NOR2xp67_ASAP7_75t_L g1841 ( 
.A(n_1822),
.B(n_1796),
.Y(n_1841)
);

NAND2xp33_ASAP7_75t_SL g1842 ( 
.A(n_1816),
.B(n_1792),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1821),
.B(n_1802),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1826),
.Y(n_1844)
);

OAI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1813),
.A2(n_1797),
.B1(n_1793),
.B2(n_1812),
.Y(n_1845)
);

AOI32xp33_ASAP7_75t_L g1846 ( 
.A1(n_1823),
.A2(n_1796),
.A3(n_1807),
.B1(n_1805),
.B2(n_1811),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1832),
.A2(n_1809),
.B1(n_1803),
.B2(n_1807),
.C(n_1761),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1827),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1825),
.A2(n_1807),
.B1(n_1707),
.B2(n_1691),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1819),
.A2(n_1809),
.B(n_1579),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1828),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1833),
.A2(n_1691),
.B1(n_1623),
.B2(n_1661),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1831),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1815),
.A2(n_1580),
.B(n_1703),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1822),
.A2(n_1623),
.B1(n_1639),
.B2(n_1653),
.Y(n_1855)
);

OAI21xp33_ASAP7_75t_L g1856 ( 
.A1(n_1823),
.A2(n_1781),
.B(n_1623),
.Y(n_1856)
);

AO32x1_ASAP7_75t_L g1857 ( 
.A1(n_1838),
.A2(n_1721),
.A3(n_1766),
.B1(n_1814),
.B2(n_1818),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1820),
.A2(n_1703),
.B(n_1725),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1839),
.B(n_1830),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1850),
.A2(n_1847),
.B(n_1845),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1841),
.Y(n_1861)
);

OAI321xp33_ASAP7_75t_L g1862 ( 
.A1(n_1846),
.A2(n_1837),
.A3(n_1836),
.B1(n_1829),
.B2(n_1817),
.C(n_1835),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1843),
.B(n_1834),
.Y(n_1863)
);

NAND2x1_ASAP7_75t_L g1864 ( 
.A(n_1849),
.B(n_1721),
.Y(n_1864)
);

OA21x2_ASAP7_75t_SL g1865 ( 
.A1(n_1842),
.A2(n_1726),
.B(n_1725),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1844),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1840),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1848),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1851),
.Y(n_1869)
);

XOR2x2_ASAP7_75t_L g1870 ( 
.A(n_1854),
.B(n_1555),
.Y(n_1870)
);

NAND4xp25_ASAP7_75t_L g1871 ( 
.A(n_1860),
.B(n_1856),
.C(n_1853),
.D(n_1855),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1861),
.B(n_1858),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1867),
.A2(n_1852),
.B1(n_1857),
.B2(n_1726),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1859),
.Y(n_1874)
);

OAI211xp5_ASAP7_75t_L g1875 ( 
.A1(n_1867),
.A2(n_1857),
.B(n_1588),
.C(n_1597),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1862),
.B(n_1857),
.Y(n_1876)
);

AOI222xp33_ASAP7_75t_L g1877 ( 
.A1(n_1862),
.A2(n_1718),
.B1(n_1715),
.B2(n_1713),
.C1(n_1726),
.C2(n_1725),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1863),
.B(n_1718),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1866),
.B(n_1766),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1868),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1870),
.B(n_1869),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1864),
.B(n_1713),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1881),
.B(n_1865),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1876),
.A2(n_1594),
.B1(n_1639),
.B2(n_1653),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1871),
.A2(n_1726),
.B1(n_1725),
.B2(n_1597),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1874),
.Y(n_1886)
);

AOI311xp33_ASAP7_75t_L g1887 ( 
.A1(n_1875),
.A2(n_1670),
.A3(n_1667),
.B(n_1700),
.C(n_1673),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1872),
.A2(n_1726),
.B1(n_1714),
.B2(n_1706),
.C(n_1716),
.Y(n_1888)
);

AOI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1884),
.A2(n_1873),
.B1(n_1878),
.B2(n_1880),
.C(n_1882),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1886),
.B(n_1879),
.Y(n_1890)
);

O2A1O1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1883),
.A2(n_1877),
.B(n_1714),
.C(n_1700),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1888),
.A2(n_1706),
.B(n_1696),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1885),
.Y(n_1893)
);

AND3x2_ASAP7_75t_L g1894 ( 
.A(n_1887),
.B(n_1564),
.C(n_1648),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1889),
.B(n_1733),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1893),
.Y(n_1896)
);

XNOR2xp5_ASAP7_75t_L g1897 ( 
.A(n_1894),
.B(n_1566),
.Y(n_1897)
);

XOR2xp5_ASAP7_75t_L g1898 ( 
.A(n_1891),
.B(n_1569),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1890),
.Y(n_1899)
);

NAND4xp75_ASAP7_75t_L g1900 ( 
.A(n_1899),
.B(n_1892),
.C(n_1550),
.D(n_1545),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1896),
.B(n_1895),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1898),
.B(n_1714),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1900),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1897),
.B1(n_1902),
.B2(n_1901),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1904),
.Y(n_1905)
);

AOI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1904),
.A2(n_1733),
.B1(n_1706),
.B2(n_1716),
.Y(n_1906)
);

OAI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1716),
.B(n_1706),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1905),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1907),
.B1(n_1716),
.B2(n_1674),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1908),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1910),
.A2(n_1674),
.B1(n_1733),
.B2(n_1670),
.Y(n_1911)
);

OAI32xp33_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1909),
.A3(n_1727),
.B1(n_1692),
.B2(n_1675),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1912),
.Y(n_1913)
);

OAI221xp5_ASAP7_75t_R g1914 ( 
.A1(n_1913),
.A2(n_1674),
.B1(n_1727),
.B2(n_1697),
.C(n_1695),
.Y(n_1914)
);

AOI211xp5_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1545),
.B(n_1550),
.C(n_1599),
.Y(n_1915)
);


endmodule