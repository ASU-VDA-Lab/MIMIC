module fake_jpeg_20006_n_237 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_27),
.Y(n_67)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_54),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_70),
.B1(n_73),
.B2(n_53),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_30),
.Y(n_104)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_25),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_66),
.A3(n_45),
.B1(n_34),
.B2(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_27),
.B(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_25),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_22),
.C(n_17),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_30),
.C(n_29),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_19),
.B1(n_22),
.B2(n_17),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_43),
.B1(n_45),
.B2(n_34),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_38),
.A2(n_19),
.B1(n_33),
.B2(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_32),
.B1(n_31),
.B2(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_78),
.B(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_94),
.B1(n_69),
.B2(n_53),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_100),
.B1(n_61),
.B2(n_57),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_34),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_92),
.Y(n_114)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_21),
.B1(n_29),
.B2(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_14),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_3),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_107),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_24),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_52),
.B1(n_62),
.B2(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_68),
.B1(n_53),
.B2(n_52),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_131),
.B1(n_102),
.B2(n_83),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_49),
.B1(n_75),
.B2(n_60),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_120),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_59),
.A3(n_51),
.B1(n_30),
.B2(n_29),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_75),
.B1(n_51),
.B2(n_48),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_127),
.B(n_79),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_99),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_24),
.A3(n_20),
.B1(n_75),
.B2(n_7),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_4),
.B(n_5),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_80),
.B(n_95),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_8),
.B(n_9),
.Y(n_129)
);

NAND2xp67_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_10),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_8),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_123),
.C(n_110),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_128),
.B1(n_126),
.B2(n_125),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_84),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_84),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_80),
.B(n_86),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_127),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_86),
.B1(n_101),
.B2(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_124),
.B1(n_126),
.B2(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_89),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_89),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_106),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_165),
.C(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_141),
.B1(n_134),
.B2(n_136),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_111),
.C(n_117),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_116),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_175),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_120),
.B1(n_133),
.B2(n_131),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_143),
.B1(n_145),
.B2(n_151),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_121),
.C(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_11),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_12),
.C(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_147),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_146),
.B(n_142),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_185),
.B(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_154),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_188),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_187),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_142),
.B(n_137),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_149),
.B(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_140),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_173),
.B1(n_176),
.B2(n_159),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_193),
.B1(n_164),
.B2(n_179),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_143),
.B1(n_139),
.B2(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_192),
.B1(n_182),
.B2(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_173),
.A3(n_165),
.B1(n_163),
.B2(n_177),
.C1(n_158),
.C2(n_176),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_187),
.B(n_190),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_174),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_205),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_191),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_153),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_214),
.C(n_194),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_188),
.B(n_185),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_210),
.B(n_215),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_178),
.B(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_178),
.C(n_12),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_12),
.C(n_13),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_201),
.B(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_219),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_222),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_196),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_197),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_196),
.Y(n_222)
);

OAI21x1_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_197),
.B(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_226),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_212),
.C(n_214),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_224),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_229),
.B(n_227),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_218),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_236),
.B(n_235),
.Y(n_237)
);


endmodule