module fake_jpeg_15455_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_16),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_1),
.C(n_2),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_8),
.C(n_13),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_20),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.C(n_10),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_7),
.B1(n_21),
.B2(n_10),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_33),
.C(n_34),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_7),
.B1(n_9),
.B2(n_27),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_34),
.B(n_30),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.C(n_29),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_33),
.Y(n_40)
);

OAI321xp33_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_37),
.A3(n_32),
.B1(n_26),
.B2(n_23),
.C(n_7),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_9),
.B1(n_32),
.B2(n_30),
.Y(n_43)
);


endmodule