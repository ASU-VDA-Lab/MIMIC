module real_aes_9008_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_756;
wire n_713;
wire n_728;
wire n_598;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_162;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_1), .A2(n_139), .B(n_143), .C(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_2), .A2(n_173), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g516 ( .A(n_3), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_4), .B(n_240), .Y(n_259) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_5), .A2(n_173), .B(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_L g139 ( .A(n_6), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g214 ( .A(n_7), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_8), .B(n_41), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_8), .B(n_41), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_9), .A2(n_172), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_10), .B(n_151), .Y(n_226) );
INVx1_ASAP7_75t_L g486 ( .A(n_11), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_12), .B(n_254), .Y(n_541) );
INVx1_ASAP7_75t_L g159 ( .A(n_13), .Y(n_159) );
INVx1_ASAP7_75t_L g553 ( .A(n_14), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_15), .A2(n_149), .B(n_236), .C(n_238), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_16), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_17), .B(n_504), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_18), .B(n_173), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_19), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_20), .A2(n_254), .B(n_269), .C(n_271), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_21), .B(n_240), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_22), .B(n_151), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_23), .A2(n_181), .B(n_238), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_24), .B(n_151), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_25), .Y(n_190) );
INVx1_ASAP7_75t_L g147 ( .A(n_26), .Y(n_147) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_27), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_28), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_29), .B(n_151), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_30), .A2(n_31), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_30), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_31), .Y(n_751) );
INVx1_ASAP7_75t_L g179 ( .A(n_32), .Y(n_179) );
INVx1_ASAP7_75t_L g495 ( .A(n_33), .Y(n_495) );
INVx2_ASAP7_75t_L g137 ( .A(n_34), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_35), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_36), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
INVxp67_ASAP7_75t_L g180 ( .A(n_37), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_38), .A2(n_143), .B(n_146), .C(n_154), .Y(n_142) );
CKINVDCx14_ASAP7_75t_R g252 ( .A(n_39), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_40), .A2(n_139), .B(n_143), .C(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g494 ( .A(n_42), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_43), .A2(n_198), .B(n_212), .C(n_213), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_44), .B(n_151), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_45), .A2(n_749), .B1(n_750), .B2(n_753), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_45), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_46), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_47), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_48), .A2(n_104), .B1(n_117), .B2(n_762), .Y(n_103) );
INVx1_ASAP7_75t_L g267 ( .A(n_49), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_50), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_51), .B(n_173), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_52), .B(n_462), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_53), .A2(n_143), .B1(n_271), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_54), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_55), .Y(n_513) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_56), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_57), .A2(n_212), .B(n_257), .C(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_58), .Y(n_569) );
INVx1_ASAP7_75t_L g483 ( .A(n_59), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_60), .A2(n_89), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_60), .Y(n_454) );
INVx1_ASAP7_75t_L g140 ( .A(n_61), .Y(n_140) );
INVx1_ASAP7_75t_L g158 ( .A(n_62), .Y(n_158) );
INVx1_ASAP7_75t_SL g256 ( .A(n_63), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_64), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_65), .B(n_240), .Y(n_273) );
INVx1_ASAP7_75t_L g193 ( .A(n_66), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_SL g503 ( .A1(n_67), .A2(n_257), .B(n_504), .C(n_505), .Y(n_503) );
INVxp67_ASAP7_75t_L g506 ( .A(n_68), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_69), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_69), .Y(n_124) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_71), .A2(n_173), .B(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_72), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_73), .A2(n_173), .B(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_74), .Y(n_498) );
INVx1_ASAP7_75t_L g563 ( .A(n_75), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_76), .A2(n_172), .B(n_174), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_77), .Y(n_141) );
INVx1_ASAP7_75t_L g234 ( .A(n_78), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_79), .A2(n_139), .B(n_143), .C(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_80), .A2(n_173), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g237 ( .A(n_81), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_82), .B(n_148), .Y(n_529) );
INVx2_ASAP7_75t_L g156 ( .A(n_83), .Y(n_156) );
INVx1_ASAP7_75t_L g225 ( .A(n_84), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_85), .B(n_504), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_86), .A2(n_139), .B(n_143), .C(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g457 ( .A(n_87), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g469 ( .A(n_87), .B(n_459), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_88), .A2(n_143), .B(n_192), .C(n_200), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_89), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_90), .B(n_155), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_91), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_92), .A2(n_139), .B(n_143), .C(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_93), .Y(n_545) );
INVx1_ASAP7_75t_L g502 ( .A(n_94), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_95), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_96), .B(n_148), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_97), .B(n_163), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_98), .B(n_163), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_99), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g270 ( .A(n_100), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_101), .A2(n_173), .B(n_501), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_102), .A2(n_466), .B1(n_747), .B2(n_748), .C1(n_754), .C2(n_757), .Y(n_465) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g762 ( .A(n_106), .Y(n_762) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g459 ( .A(n_112), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g472 ( .A(n_113), .B(n_459), .Y(n_472) );
NOR2x2_ASAP7_75t_L g759 ( .A(n_113), .B(n_458), .Y(n_759) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_464), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g761 ( .A(n_120), .Y(n_761) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_455), .B(n_461), .Y(n_122) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
XOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_452), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_127), .A2(n_467), .B1(n_470), .B2(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g755 ( .A(n_127), .Y(n_755) );
OR4x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_342), .C(n_389), .D(n_429), .Y(n_127) );
NAND3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_288), .C(n_317), .Y(n_128) );
AOI211xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_203), .B(n_241), .C(n_281), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_130), .A2(n_301), .B(n_318), .C(n_322), .Y(n_317) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_165), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_132), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_SL g284 ( .A(n_132), .Y(n_284) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_132), .Y(n_296) );
AND2x4_ASAP7_75t_L g300 ( .A(n_132), .B(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g311 ( .A(n_132), .B(n_188), .Y(n_311) );
OR2x2_ASAP7_75t_L g335 ( .A(n_132), .B(n_244), .Y(n_335) );
AND2x2_ASAP7_75t_L g348 ( .A(n_132), .B(n_249), .Y(n_348) );
AND2x2_ASAP7_75t_L g388 ( .A(n_132), .B(n_374), .Y(n_388) );
AND2x2_ASAP7_75t_L g395 ( .A(n_132), .B(n_358), .Y(n_395) );
AND2x2_ASAP7_75t_L g425 ( .A(n_132), .B(n_166), .Y(n_425) );
OR2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_160), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_142), .C(n_155), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_134), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_134), .A2(n_222), .B(n_223), .Y(n_221) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_134), .A2(n_183), .B1(n_492), .B2(n_496), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_134), .A2(n_513), .B(n_514), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_134), .A2(n_563), .B(n_564), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
AND2x4_ASAP7_75t_L g173 ( .A(n_135), .B(n_139), .Y(n_173) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
INVx1_ASAP7_75t_L g272 ( .A(n_137), .Y(n_272) );
INVx1_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx3_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_138), .Y(n_151) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
INVx1_ASAP7_75t_L g504 ( .A(n_138), .Y(n_504) );
BUFx3_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx4_ASAP7_75t_SL g183 ( .A(n_139), .Y(n_183) );
INVx5_ASAP7_75t_L g176 ( .A(n_143), .Y(n_176) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g199 ( .A(n_144), .Y(n_199) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_144), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .C(n_152), .Y(n_146) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_148), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_148), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_149), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_149), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_149), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx4_ASAP7_75t_L g254 ( .A(n_151), .Y(n_254) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_153), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_155), .A2(n_208), .B(n_215), .Y(n_207) );
INVx1_ASAP7_75t_L g220 ( .A(n_155), .Y(n_220) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_155), .A2(n_548), .B(n_554), .Y(n_547) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g164 ( .A(n_156), .B(n_157), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_189), .B(n_201), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_162), .B(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g240 ( .A(n_162), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g531 ( .A(n_162), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_163), .Y(n_231) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_163), .A2(n_500), .B(n_507), .Y(n_499) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_165), .B(n_352), .Y(n_364) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_187), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_166), .B(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g302 ( .A(n_166), .B(n_187), .Y(n_302) );
BUFx3_ASAP7_75t_L g310 ( .A(n_166), .Y(n_310) );
OR2x2_ASAP7_75t_L g331 ( .A(n_166), .B(n_206), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_166), .B(n_352), .Y(n_442) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_184), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_168), .A2(n_245), .B(n_246), .Y(n_244) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_168), .A2(n_562), .B(n_568), .Y(n_561) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_169), .A2(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_170), .A2(n_491), .B(n_497), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_170), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_170), .A2(n_512), .B(n_519), .Y(n_511) );
INVx1_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g209 ( .A1(n_176), .A2(n_183), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g233 ( .A1(n_176), .A2(n_183), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_176), .A2(n_183), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_176), .A2(n_183), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_176), .A2(n_183), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_176), .A2(n_183), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_176), .A2(n_183), .B(n_550), .C(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_181), .B(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_181), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_181), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_182), .A2(n_195), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
INVx1_ASAP7_75t_L g246 ( .A(n_184), .Y(n_246) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_186), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_186), .A2(n_537), .B(n_544), .Y(n_536) );
AND2x2_ASAP7_75t_L g247 ( .A(n_187), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g295 ( .A(n_187), .Y(n_295) );
AND2x2_ASAP7_75t_L g358 ( .A(n_187), .B(n_249), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_187), .A2(n_361), .B1(n_363), .B2(n_365), .C(n_366), .Y(n_360) );
AND2x2_ASAP7_75t_L g374 ( .A(n_187), .B(n_244), .Y(n_374) );
AND2x2_ASAP7_75t_L g400 ( .A(n_187), .B(n_284), .Y(n_400) );
INVx2_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g280 ( .A(n_188), .B(n_249), .Y(n_280) );
BUFx2_ASAP7_75t_L g414 ( .A(n_188), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_194), .A2(n_197), .B(n_225), .C(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_197), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_197), .A2(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OAI32xp33_ASAP7_75t_L g380 ( .A1(n_204), .A2(n_341), .A3(n_355), .B1(n_381), .B2(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_216), .Y(n_204) );
AND2x2_ASAP7_75t_L g321 ( .A(n_205), .B(n_263), .Y(n_321) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g303 ( .A(n_206), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_206), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g375 ( .A(n_206), .B(n_263), .Y(n_375) );
AND2x2_ASAP7_75t_L g386 ( .A(n_206), .B(n_278), .Y(n_386) );
BUFx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g287 ( .A(n_207), .B(n_264), .Y(n_287) );
AND2x2_ASAP7_75t_L g291 ( .A(n_207), .B(n_264), .Y(n_291) );
AND2x2_ASAP7_75t_L g326 ( .A(n_207), .B(n_277), .Y(n_326) );
AND2x2_ASAP7_75t_L g333 ( .A(n_207), .B(n_229), .Y(n_333) );
OAI211xp5_ASAP7_75t_L g338 ( .A1(n_207), .A2(n_284), .B(n_295), .C(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g392 ( .A(n_207), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_207), .B(n_218), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_216), .B(n_275), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_216), .B(n_291), .Y(n_381) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g286 ( .A(n_217), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_229), .Y(n_217) );
AND2x2_ASAP7_75t_L g278 ( .A(n_218), .B(n_230), .Y(n_278) );
OR2x2_ASAP7_75t_L g293 ( .A(n_218), .B(n_230), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_218), .B(n_277), .Y(n_316) );
INVx1_ASAP7_75t_L g320 ( .A(n_218), .Y(n_320) );
AND2x2_ASAP7_75t_L g339 ( .A(n_218), .B(n_276), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_218), .A2(n_304), .B1(n_350), .B2(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_218), .B(n_392), .Y(n_416) );
AND2x2_ASAP7_75t_L g431 ( .A(n_218), .B(n_291), .Y(n_431) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx3_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
AND2x2_ASAP7_75t_L g305 ( .A(n_219), .B(n_230), .Y(n_305) );
AND2x2_ASAP7_75t_L g307 ( .A(n_219), .B(n_263), .Y(n_307) );
AND3x2_ASAP7_75t_L g369 ( .A(n_219), .B(n_333), .C(n_370), .Y(n_369) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_227), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_220), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_220), .B(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_220), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g404 ( .A(n_229), .B(n_276), .Y(n_404) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g263 ( .A(n_230), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_230), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_230), .B(n_275), .Y(n_337) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_230), .B(n_316), .C(n_392), .Y(n_444) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_239), .Y(n_230) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_231), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_231), .A2(n_265), .B(n_273), .Y(n_264) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_240), .A2(n_481), .B(n_487), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_260), .B1(n_274), .B2(n_279), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_244), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g356 ( .A(n_244), .Y(n_356) );
OAI31xp33_ASAP7_75t_L g372 ( .A1(n_247), .A2(n_373), .A3(n_374), .B(n_375), .Y(n_372) );
AND2x2_ASAP7_75t_L g397 ( .A(n_247), .B(n_284), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_247), .B(n_310), .Y(n_443) );
AND2x2_ASAP7_75t_L g352 ( .A(n_248), .B(n_284), .Y(n_352) );
AND2x2_ASAP7_75t_L g413 ( .A(n_248), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g283 ( .A(n_249), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g341 ( .A(n_249), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_258), .Y(n_542) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_261), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_262), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AOI221x1_ASAP7_75t_SL g329 ( .A1(n_263), .A2(n_330), .B1(n_332), .B2(n_334), .C(n_336), .Y(n_329) );
INVx2_ASAP7_75t_L g277 ( .A(n_264), .Y(n_277) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_264), .Y(n_371) );
INVx2_ASAP7_75t_L g518 ( .A(n_271), .Y(n_518) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g359 ( .A(n_274), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_275), .B(n_292), .Y(n_384) );
INVx1_ASAP7_75t_SL g447 ( .A(n_275), .Y(n_447) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g365 ( .A(n_278), .B(n_291), .Y(n_365) );
INVx1_ASAP7_75t_L g433 ( .A(n_279), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_279), .B(n_362), .Y(n_446) );
INVx2_ASAP7_75t_SL g285 ( .A(n_280), .Y(n_285) );
AND2x2_ASAP7_75t_L g328 ( .A(n_280), .B(n_284), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_280), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_280), .B(n_355), .Y(n_382) );
AOI21xp33_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_285), .B(n_286), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_283), .B(n_355), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_283), .B(n_310), .Y(n_451) );
OR2x2_ASAP7_75t_L g323 ( .A(n_284), .B(n_302), .Y(n_323) );
AND2x2_ASAP7_75t_L g422 ( .A(n_284), .B(n_413), .Y(n_422) );
OAI22xp5_ASAP7_75t_SL g297 ( .A1(n_285), .A2(n_298), .B1(n_303), .B2(n_306), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_285), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g345 ( .A(n_287), .B(n_293), .Y(n_345) );
INVx1_ASAP7_75t_L g409 ( .A(n_287), .Y(n_409) );
AOI311xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_294), .A3(n_296), .B(n_297), .C(n_308), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_292), .A2(n_424), .B1(n_436), .B2(n_439), .C(n_441), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_292), .B(n_447), .Y(n_449) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_295), .A2(n_337), .B(n_338), .C(n_340), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_SL g405 ( .A1(n_299), .A2(n_301), .B(n_406), .C(n_407), .Y(n_405) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_300), .B(n_374), .Y(n_440) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_303), .A2(n_323), .B1(n_324), .B2(n_327), .C(n_329), .Y(n_322) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g325 ( .A(n_305), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g408 ( .A(n_305), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_309), .A2(n_367), .B(n_368), .C(n_372), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_310), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_310), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_316), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_320), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g434 ( .A(n_323), .Y(n_434) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_326), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_326), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g438 ( .A(n_326), .Y(n_438) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g379 ( .A(n_328), .B(n_355), .Y(n_379) );
INVx1_ASAP7_75t_SL g373 ( .A(n_335), .Y(n_373) );
INVx1_ASAP7_75t_L g350 ( .A(n_341), .Y(n_350) );
NAND3xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_360), .C(n_376), .Y(n_342) );
AOI322xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .A3(n_347), .B1(n_349), .B2(n_353), .C1(n_357), .C2(n_359), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g396 ( .A1(n_344), .A2(n_397), .B(n_398), .C(n_405), .Y(n_396) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_347), .A2(n_368), .B1(n_399), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g357 ( .A(n_355), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_355), .B(n_395), .Y(n_394) );
AOI32xp33_ASAP7_75t_L g445 ( .A1(n_355), .A2(n_446), .A3(n_447), .B1(n_448), .B2(n_450), .Y(n_445) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g367 ( .A(n_358), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_358), .A2(n_411), .B1(n_415), .B2(n_417), .C(n_420), .Y(n_410) );
AND2x2_ASAP7_75t_L g424 ( .A(n_358), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g427 ( .A(n_362), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g437 ( .A(n_362), .B(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g428 ( .A(n_371), .B(n_392), .Y(n_428) );
AOI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_380), .C(n_383), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_393), .B(n_396), .C(n_410), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_404), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_416), .Y(n_419) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_426), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI211xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_432), .B(n_435), .C(n_445), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_457), .Y(n_463) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_461), .A2(n_465), .B(n_760), .Y(n_464) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22x1_ASAP7_75t_L g754 ( .A1(n_467), .A2(n_470), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g756 ( .A(n_474), .Y(n_756) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND3x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_669), .C(n_714), .Y(n_475) );
NOR4xp25_ASAP7_75t_L g476 ( .A(n_477), .B(n_592), .C(n_633), .D(n_650), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_508), .B(n_522), .C(n_555), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_479), .B(n_509), .Y(n_508) );
NOR4xp25_ASAP7_75t_L g616 ( .A(n_479), .B(n_610), .C(n_617), .D(n_623), .Y(n_616) );
AND2x2_ASAP7_75t_L g689 ( .A(n_479), .B(n_578), .Y(n_689) );
AND2x2_ASAP7_75t_L g708 ( .A(n_479), .B(n_654), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_479), .B(n_703), .Y(n_717) );
AND2x2_ASAP7_75t_L g730 ( .A(n_479), .B(n_521), .Y(n_730) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g575 ( .A(n_480), .Y(n_575) );
AND2x2_ASAP7_75t_L g582 ( .A(n_480), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g632 ( .A(n_480), .B(n_489), .Y(n_632) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_480), .B(n_578), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_480), .B(n_489), .Y(n_647) );
AND2x2_ASAP7_75t_L g656 ( .A(n_480), .B(n_581), .Y(n_656) );
BUFx2_ASAP7_75t_L g679 ( .A(n_480), .Y(n_679) );
AND2x2_ASAP7_75t_L g683 ( .A(n_480), .B(n_499), .Y(n_683) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_499), .Y(n_488) );
AND2x2_ASAP7_75t_L g521 ( .A(n_489), .B(n_499), .Y(n_521) );
BUFx2_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_489), .A2(n_618), .B1(n_620), .B2(n_621), .Y(n_617) );
OR2x2_ASAP7_75t_L g639 ( .A(n_489), .B(n_511), .Y(n_639) );
AND2x2_ASAP7_75t_L g703 ( .A(n_489), .B(n_581), .Y(n_703) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g571 ( .A(n_490), .B(n_511), .Y(n_571) );
AND2x2_ASAP7_75t_L g578 ( .A(n_490), .B(n_499), .Y(n_578) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_490), .Y(n_620) );
OR2x2_ASAP7_75t_L g655 ( .A(n_490), .B(n_510), .Y(n_655) );
INVx1_ASAP7_75t_L g574 ( .A(n_499), .Y(n_574) );
INVx3_ASAP7_75t_L g583 ( .A(n_499), .Y(n_583) );
BUFx2_ASAP7_75t_L g607 ( .A(n_499), .Y(n_607) );
AND2x2_ASAP7_75t_L g640 ( .A(n_499), .B(n_575), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_508), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_510), .B(n_583), .Y(n_587) );
INVx1_ASAP7_75t_L g615 ( .A(n_510), .Y(n_615) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
INVx1_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
NAND2x1_ASAP7_75t_SL g522 ( .A(n_523), .B(n_533), .Y(n_522) );
AND2x2_ASAP7_75t_L g591 ( .A(n_523), .B(n_546), .Y(n_591) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_523), .Y(n_665) );
AND2x2_ASAP7_75t_L g692 ( .A(n_523), .B(n_612), .Y(n_692) );
AND2x2_ASAP7_75t_L g700 ( .A(n_523), .B(n_662), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_523), .B(n_558), .Y(n_727) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g559 ( .A(n_524), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g576 ( .A(n_524), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g597 ( .A(n_524), .Y(n_597) );
INVx1_ASAP7_75t_L g603 ( .A(n_524), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_524), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g636 ( .A(n_524), .B(n_561), .Y(n_636) );
OR2x2_ASAP7_75t_L g674 ( .A(n_524), .B(n_629), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g686 ( .A1(n_524), .A2(n_687), .A3(n_690), .B1(n_691), .B2(n_692), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_524), .B(n_662), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_524), .B(n_622), .Y(n_737) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g648 ( .A(n_534), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_546), .Y(n_534) );
INVx1_ASAP7_75t_L g610 ( .A(n_535), .Y(n_610) );
AND2x2_ASAP7_75t_L g612 ( .A(n_535), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_535), .B(n_560), .Y(n_629) );
AND2x2_ASAP7_75t_L g662 ( .A(n_535), .B(n_638), .Y(n_662) );
AND2x2_ASAP7_75t_L g699 ( .A(n_535), .B(n_561), .Y(n_699) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g558 ( .A(n_536), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_536), .B(n_560), .Y(n_589) );
AND2x2_ASAP7_75t_L g596 ( .A(n_536), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g637 ( .A(n_536), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_542), .Y(n_539) );
INVx2_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_546), .B(n_560), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_546), .B(n_604), .Y(n_685) );
INVx1_ASAP7_75t_L g707 ( .A(n_546), .Y(n_707) );
INVx1_ASAP7_75t_L g724 ( .A(n_546), .Y(n_724) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g577 ( .A(n_547), .B(n_560), .Y(n_577) );
AND2x2_ASAP7_75t_L g599 ( .A(n_547), .B(n_561), .Y(n_599) );
INVx1_ASAP7_75t_L g638 ( .A(n_547), .Y(n_638) );
AOI221x1_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_570), .B1(n_576), .B2(n_578), .C(n_579), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_556), .A2(n_643), .B1(n_710), .B2(n_711), .Y(n_709) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND2x2_ASAP7_75t_L g601 ( .A(n_557), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g696 ( .A(n_557), .B(n_576), .Y(n_696) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g652 ( .A(n_558), .B(n_577), .Y(n_652) );
INVx1_ASAP7_75t_L g664 ( .A(n_559), .Y(n_664) );
AND2x2_ASAP7_75t_L g675 ( .A(n_559), .B(n_662), .Y(n_675) );
AND2x2_ASAP7_75t_L g742 ( .A(n_559), .B(n_637), .Y(n_742) );
INVx2_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_571), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g694 ( .A(n_571), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_572), .B(n_655), .Y(n_658) );
INVx3_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_573), .A2(n_694), .B(n_739), .Y(n_738) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NOR2xp33_ASAP7_75t_SL g716 ( .A(n_576), .B(n_602), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_577), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g668 ( .A(n_577), .B(n_596), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_577), .B(n_603), .Y(n_745) );
AND2x2_ASAP7_75t_L g614 ( .A(n_578), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g681 ( .A(n_578), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B(n_588), .Y(n_579) );
NAND2x1_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_581), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g630 ( .A(n_581), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g642 ( .A(n_581), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_581), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g666 ( .A(n_582), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_582), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_582), .B(n_585), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_585), .A2(n_624), .B(n_654), .C(n_656), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_585), .A2(n_672), .B1(n_675), .B2(n_676), .C(n_680), .Y(n_671) );
AND2x2_ASAP7_75t_L g667 ( .A(n_586), .B(n_620), .Y(n_667) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g627 ( .A(n_591), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g698 ( .A(n_591), .B(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_600), .C(n_625), .Y(n_592) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_593), .B(n_712), .C(n_713), .Y(n_711) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
OR2x2_ASAP7_75t_L g684 ( .A(n_595), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B1(n_608), .B2(n_614), .C(n_616), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_602), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g624 ( .A(n_607), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_607), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_663) );
OR2x2_ASAP7_75t_L g744 ( .A(n_607), .B(n_655), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVxp67_ASAP7_75t_L g718 ( .A(n_610), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_612), .B(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_L g619 ( .A(n_613), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_615), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_615), .B(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_615), .B(n_682), .Y(n_721) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_619), .Y(n_645) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g735 ( .A(n_624), .B(n_655), .Y(n_735) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g713 ( .A(n_630), .Y(n_713) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI322xp33_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_639), .A3(n_640), .B1(n_641), .B2(n_644), .C1(n_646), .C2(n_648), .Y(n_633) );
OAI322xp33_ASAP7_75t_L g715 ( .A1(n_634), .A2(n_716), .A3(n_717), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_722), .Y(n_715) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx4_ASAP7_75t_L g649 ( .A(n_636), .Y(n_649) );
AND2x2_ASAP7_75t_L g710 ( .A(n_636), .B(n_662), .Y(n_710) );
AND2x2_ASAP7_75t_L g723 ( .A(n_636), .B(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_639), .Y(n_734) );
INVx1_ASAP7_75t_L g712 ( .A(n_640), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OR2x2_ASAP7_75t_L g646 ( .A(n_642), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g729 ( .A(n_642), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_642), .B(n_683), .Y(n_740) );
OR2x2_ASAP7_75t_L g673 ( .A(n_645), .B(n_674), .Y(n_673) );
INVxp33_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
OAI221xp5_ASAP7_75t_SL g650 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_657), .C(n_659), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g706 ( .A(n_649), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g733 ( .A(n_649), .Y(n_733) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx3_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_656), .A2(n_681), .A3(n_698), .B1(n_700), .B2(n_701), .C1(n_704), .C2(n_708), .Y(n_697) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_667), .B2(n_668), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_693), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_686), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_674), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
NAND2xp33_ASAP7_75t_SL g691 ( .A(n_677), .B(n_688), .Y(n_691) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
OAI322xp33_ASAP7_75t_L g731 ( .A1(n_679), .A2(n_732), .A3(n_734), .B1(n_735), .B2(n_736), .C1(n_738), .C2(n_741), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_689), .B(n_737), .Y(n_746) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_695), .B(n_697), .C(n_709), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR4xp25_ASAP7_75t_L g714 ( .A(n_715), .B(n_725), .C(n_731), .D(n_743), .Y(n_714) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx14_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g743 ( .A1(n_744), .A2(n_745), .B(n_746), .Y(n_743) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule