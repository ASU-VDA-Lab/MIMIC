module real_aes_6401_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g268 ( .A1(n_0), .A2(n_269), .B(n_270), .C(n_273), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_1), .B(n_210), .Y(n_274) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_3), .B(n_180), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_4), .A2(n_150), .B(n_153), .C(n_478), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_5), .A2(n_170), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_6), .A2(n_170), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_7), .B(n_210), .Y(n_524) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_8), .A2(n_137), .B(n_190), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_9), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_9), .Y(n_744) );
AND2x6_ASAP7_75t_L g150 ( .A(n_10), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_11), .A2(n_150), .B(n_153), .C(n_156), .Y(n_152) );
INVx1_ASAP7_75t_L g494 ( .A(n_12), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_13), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_13), .B(n_41), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_14), .A2(n_45), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_14), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_15), .B(n_160), .Y(n_480) );
INVx1_ASAP7_75t_L g142 ( .A(n_16), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_17), .B(n_180), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_18), .A2(n_158), .B(n_502), .C(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_19), .B(n_210), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_20), .B(n_234), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_21), .A2(n_153), .B(n_197), .C(n_230), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_22), .A2(n_162), .B(n_272), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_23), .B(n_160), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_24), .B(n_160), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_25), .Y(n_552) );
INVx1_ASAP7_75t_L g544 ( .A(n_26), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_27), .A2(n_153), .B(n_193), .C(n_197), .Y(n_192) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_29), .Y(n_476) );
INVx1_ASAP7_75t_L g535 ( .A(n_30), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_31), .A2(n_170), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g148 ( .A(n_32), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_33), .A2(n_172), .B(n_183), .C(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_34), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_35), .A2(n_272), .B(n_521), .C(n_523), .Y(n_520) );
INVxp67_ASAP7_75t_L g536 ( .A(n_36), .Y(n_536) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_37), .A2(n_78), .B1(n_451), .B2(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_37), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_38), .B(n_195), .Y(n_194) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_39), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_40), .A2(n_153), .B(n_197), .C(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_42), .A2(n_273), .B(n_492), .C(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_43), .B(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_44), .Y(n_165) );
INVx1_ASAP7_75t_L g742 ( .A(n_45), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_46), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_47), .B(n_170), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_48), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_49), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_50), .A2(n_172), .B(n_174), .C(n_183), .Y(n_171) );
INVx1_ASAP7_75t_L g271 ( .A(n_51), .Y(n_271) );
INVx1_ASAP7_75t_L g175 ( .A(n_52), .Y(n_175) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_53), .A2(n_462), .B1(n_735), .B2(n_736), .C1(n_745), .C2(n_748), .Y(n_461) );
INVx1_ASAP7_75t_L g509 ( .A(n_54), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_55), .B(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_56), .A2(n_59), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_56), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_57), .Y(n_237) );
CKINVDCx14_ASAP7_75t_R g490 ( .A(n_58), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_59), .Y(n_125) );
INVx1_ASAP7_75t_L g151 ( .A(n_60), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_61), .B(n_170), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_62), .B(n_210), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_63), .A2(n_204), .B(n_206), .C(n_208), .Y(n_203) );
INVx1_ASAP7_75t_L g141 ( .A(n_64), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_65), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g522 ( .A(n_66), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_68), .B(n_180), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_69), .B(n_210), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_70), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g555 ( .A(n_71), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_72), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_73), .B(n_177), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_74), .A2(n_153), .B(n_183), .C(n_244), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_75), .Y(n_202) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_77), .A2(n_170), .B(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_78), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_79), .A2(n_170), .B(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_80), .A2(n_228), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g500 ( .A(n_81), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_82), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_83), .B(n_176), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_84), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_85), .A2(n_170), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g503 ( .A(n_86), .Y(n_503) );
INVx2_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g479 ( .A(n_88), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_89), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_90), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g109 ( .A(n_91), .Y(n_109) );
OR2x2_ASAP7_75t_L g446 ( .A(n_91), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g465 ( .A(n_91), .B(n_448), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_92), .A2(n_153), .B(n_183), .C(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_93), .B(n_170), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_94), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_94), .Y(n_737) );
INVx1_ASAP7_75t_L g219 ( .A(n_95), .Y(n_219) );
INVxp67_ASAP7_75t_L g207 ( .A(n_96), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_97), .B(n_137), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
INVx1_ASAP7_75t_L g245 ( .A(n_100), .Y(n_245) );
INVx2_ASAP7_75t_L g512 ( .A(n_101), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_102), .A2(n_105), .B1(n_115), .B2(n_753), .Y(n_104) );
AND2x2_ASAP7_75t_L g186 ( .A(n_103), .B(n_185), .Y(n_186) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g754 ( .A(n_106), .Y(n_754) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g448 ( .A(n_108), .B(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g734 ( .A(n_109), .B(n_448), .Y(n_734) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_109), .B(n_447), .Y(n_750) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_460), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g752 ( .A(n_119), .Y(n_752) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_444), .A3(n_450), .B1(n_453), .B2(n_454), .C(n_457), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_122), .B(n_455), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_127), .B2(n_128), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22x1_ASAP7_75t_SL g462 ( .A1(n_127), .A2(n_463), .B1(n_466), .B2(n_732), .Y(n_462) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_128), .A2(n_467), .B1(n_746), .B2(n_747), .Y(n_745) );
OR3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_342), .C(n_407), .Y(n_128) );
NAND4xp25_ASAP7_75t_SL g129 ( .A(n_130), .B(n_283), .C(n_309), .D(n_332), .Y(n_129) );
AOI221xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_211), .B1(n_252), .B2(n_259), .C(n_275), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_132), .A2(n_276), .B1(n_300), .B2(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_187), .Y(n_132) );
INVx1_ASAP7_75t_SL g336 ( .A(n_133), .Y(n_336) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_167), .Y(n_133) );
OR2x2_ASAP7_75t_L g257 ( .A(n_134), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g278 ( .A(n_134), .B(n_188), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_134), .B(n_198), .Y(n_291) );
AND2x2_ASAP7_75t_L g308 ( .A(n_134), .B(n_167), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_134), .B(n_255), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_134), .B(n_307), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_134), .B(n_187), .Y(n_429) );
AOI211xp5_ASAP7_75t_SL g440 ( .A1(n_134), .A2(n_346), .B(n_441), .C(n_442), .Y(n_440) );
INVx5_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_135), .B(n_188), .Y(n_312) );
AND2x2_ASAP7_75t_L g315 ( .A(n_135), .B(n_189), .Y(n_315) );
OR2x2_ASAP7_75t_L g360 ( .A(n_135), .B(n_188), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_135), .B(n_198), .Y(n_369) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_164), .Y(n_135) );
INVx3_ASAP7_75t_L g210 ( .A(n_136), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_136), .B(n_222), .Y(n_221) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_136), .A2(n_242), .B(n_250), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_136), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_136), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_136), .B(n_547), .Y(n_546) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_136), .A2(n_551), .B(n_557), .Y(n_550) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_137), .A2(n_191), .B(n_192), .Y(n_190) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_139), .B(n_140), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_152), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g475 ( .A1(n_145), .A2(n_476), .B(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_145), .A2(n_185), .B(n_541), .C(n_542), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_145), .A2(n_552), .B(n_553), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
AND2x4_ASAP7_75t_L g170 ( .A(n_146), .B(n_150), .Y(n_170) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx3_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx1_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
INVx4_ASAP7_75t_SL g184 ( .A(n_150), .Y(n_184) );
BUFx3_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
INVx5_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_154), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_161), .Y(n_156) );
INVx5_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_158), .B(n_494), .Y(n_493) );
INVx4_ASAP7_75t_L g272 ( .A(n_160), .Y(n_272) );
INVx2_ASAP7_75t_L g492 ( .A(n_160), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_161), .A2(n_194), .B(n_196), .Y(n_193) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx2_ASAP7_75t_L g529 ( .A(n_166), .Y(n_529) );
INVx5_ASAP7_75t_SL g258 ( .A(n_167), .Y(n_258) );
AND2x2_ASAP7_75t_L g277 ( .A(n_167), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_167), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g363 ( .A(n_167), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g395 ( .A(n_167), .B(n_198), .Y(n_395) );
OR2x2_ASAP7_75t_L g401 ( .A(n_167), .B(n_291), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_167), .B(n_351), .Y(n_410) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_186), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_185), .Y(n_168) );
BUFx2_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_173), .A2(n_184), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_173), .A2(n_184), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_173), .A2(n_184), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_173), .A2(n_184), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_173), .A2(n_184), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_173), .A2(n_184), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_173), .A2(n_184), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_179), .C(n_181), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_176), .A2(n_181), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp5_ASAP7_75t_L g478 ( .A1(n_176), .A2(n_479), .B(n_480), .C(n_481), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_176), .A2(n_481), .B(n_555), .C(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx4_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_180), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g269 ( .A(n_180), .Y(n_269) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_180), .A2(n_205), .B1(n_535), .B2(n_536), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_180), .A2(n_233), .B(n_544), .C(n_545), .Y(n_543) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g273 ( .A(n_182), .Y(n_273) );
INVx1_ASAP7_75t_L g504 ( .A(n_182), .Y(n_504) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_185), .A2(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g238 ( .A(n_185), .Y(n_238) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_185), .A2(n_488), .B(n_495), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_198), .Y(n_187) );
AND2x2_ASAP7_75t_L g292 ( .A(n_188), .B(n_258), .Y(n_292) );
INVx1_ASAP7_75t_SL g305 ( .A(n_188), .Y(n_305) );
OR2x2_ASAP7_75t_L g340 ( .A(n_188), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g346 ( .A(n_188), .B(n_198), .Y(n_346) );
AND2x2_ASAP7_75t_L g404 ( .A(n_188), .B(n_255), .Y(n_404) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_189), .B(n_258), .Y(n_331) );
INVx3_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
OR2x2_ASAP7_75t_L g297 ( .A(n_198), .B(n_258), .Y(n_297) );
AND2x2_ASAP7_75t_L g307 ( .A(n_198), .B(n_305), .Y(n_307) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_198), .Y(n_355) );
AND2x2_ASAP7_75t_L g364 ( .A(n_198), .B(n_278), .Y(n_364) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_209), .Y(n_198) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_199), .A2(n_498), .B(n_505), .Y(n_497) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_199), .A2(n_507), .B(n_513), .Y(n_506) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_199), .A2(n_517), .B(n_524), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_204), .A2(n_245), .B(n_246), .C(n_247), .Y(n_244) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_205), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_205), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g233 ( .A(n_208), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_208), .B(n_534), .Y(n_533) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_210), .A2(n_265), .B(n_274), .Y(n_264) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_211), .A2(n_381), .B1(n_383), .B2(n_385), .C(n_388), .Y(n_380) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AND2x2_ASAP7_75t_L g354 ( .A(n_213), .B(n_335), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_213), .B(n_413), .Y(n_417) );
OR2x2_ASAP7_75t_L g438 ( .A(n_213), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_213), .B(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx5_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
AND2x2_ASAP7_75t_L g362 ( .A(n_214), .B(n_225), .Y(n_362) );
AND2x2_ASAP7_75t_L g423 ( .A(n_214), .B(n_302), .Y(n_423) );
AND2x2_ASAP7_75t_L g436 ( .A(n_214), .B(n_255), .Y(n_436) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_239), .Y(n_223) );
AND2x4_ASAP7_75t_L g262 ( .A(n_224), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g281 ( .A(n_224), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
AND2x2_ASAP7_75t_L g357 ( .A(n_224), .B(n_335), .Y(n_357) );
AND2x2_ASAP7_75t_L g367 ( .A(n_224), .B(n_285), .Y(n_367) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_224), .Y(n_375) );
AND2x2_ASAP7_75t_L g387 ( .A(n_224), .B(n_264), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_224), .B(n_319), .Y(n_391) );
AND2x2_ASAP7_75t_L g428 ( .A(n_224), .B(n_423), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_224), .B(n_302), .Y(n_439) );
OR2x2_ASAP7_75t_L g441 ( .A(n_224), .B(n_377), .Y(n_441) );
INVx5_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g327 ( .A(n_225), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_225), .B(n_282), .Y(n_337) );
AND2x2_ASAP7_75t_L g349 ( .A(n_225), .B(n_264), .Y(n_349) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_225), .Y(n_379) );
AND2x4_ASAP7_75t_L g413 ( .A(n_225), .B(n_263), .Y(n_413) );
OR2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_236), .Y(n_225) );
AOI21xp5_ASAP7_75t_SL g226 ( .A1(n_227), .A2(n_229), .B(n_234), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_235), .B(n_452), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_238), .A2(n_475), .B(n_482), .Y(n_474) );
BUFx2_ASAP7_75t_L g261 ( .A(n_239), .Y(n_261) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g302 ( .A(n_240), .Y(n_302) );
AND2x2_ASAP7_75t_L g335 ( .A(n_240), .B(n_264), .Y(n_335) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g282 ( .A(n_241), .B(n_264), .Y(n_282) );
BUFx2_ASAP7_75t_L g328 ( .A(n_241), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_249), .Y(n_242) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx3_ASAP7_75t_L g523 ( .A(n_248), .Y(n_523) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_254), .B(n_336), .Y(n_415) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_255), .B(n_278), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_255), .B(n_258), .Y(n_317) );
AND2x2_ASAP7_75t_L g372 ( .A(n_255), .B(n_308), .Y(n_372) );
AOI221xp5_ASAP7_75t_SL g309 ( .A1(n_256), .A2(n_310), .B1(n_318), .B2(n_320), .C(n_324), .Y(n_309) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g304 ( .A(n_257), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g345 ( .A(n_257), .B(n_346), .Y(n_345) );
OAI321xp33_ASAP7_75t_L g352 ( .A1(n_257), .A2(n_311), .A3(n_353), .B1(n_355), .B2(n_356), .C(n_358), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_258), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_261), .B(n_413), .Y(n_431) );
AND2x2_ASAP7_75t_L g318 ( .A(n_262), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_262), .B(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_263), .Y(n_294) );
AND2x2_ASAP7_75t_L g301 ( .A(n_263), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_263), .B(n_376), .Y(n_406) );
INVx1_ASAP7_75t_L g443 ( .A(n_263), .Y(n_443) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_272), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g481 ( .A(n_273), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_280), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_277), .A2(n_387), .B(n_436), .C(n_437), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_278), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_278), .B(n_316), .Y(n_382) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_282), .B(n_285), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_282), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_282), .B(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .B1(n_298), .B2(n_303), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g299 ( .A(n_285), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g334 ( .A(n_285), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_285), .B(n_328), .Y(n_370) );
OR2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_302), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_285), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g427 ( .A(n_285), .B(n_413), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B1(n_293), .B2(n_295), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g333 ( .A(n_288), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_291), .A2(n_306), .B1(n_374), .B2(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g421 ( .A(n_292), .Y(n_421) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_296), .A2(n_333), .B1(n_336), .B2(n_337), .C(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g311 ( .A(n_297), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_301), .B(n_367), .Y(n_399) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g341 ( .A(n_308), .Y(n_341) );
AND2x2_ASAP7_75t_L g350 ( .A(n_308), .B(n_351), .Y(n_350) );
NAND2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g394 ( .A(n_315), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_318), .A2(n_344), .B1(n_347), .B2(n_350), .C(n_352), .Y(n_343) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_322), .B(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B(n_329), .Y(n_324) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_329), .Y(n_426) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
OR2x2_ASAP7_75t_L g368 ( .A(n_331), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g389 ( .A(n_334), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_334), .B(n_394), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_337), .B(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_361), .C(n_380), .D(n_393), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g351 ( .A(n_346), .Y(n_351) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g384 ( .A(n_355), .B(n_360), .Y(n_384) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B(n_365), .C(n_373), .Y(n_361) );
AOI211xp5_ASAP7_75t_L g432 ( .A1(n_363), .A2(n_405), .B(n_433), .C(n_440), .Y(n_432) );
INVx1_ASAP7_75t_SL g392 ( .A(n_364), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_370), .B2(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g396 ( .A(n_370), .Y(n_396) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_376), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_376), .B(n_387), .Y(n_420) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g397 ( .A(n_387), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_392), .Y(n_388) );
INVxp33_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI322xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .A3(n_397), .B1(n_398), .B2(n_400), .C1(n_402), .C2(n_405), .Y(n_393) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_425), .C(n_432), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B1(n_414), .B2(n_416), .C(n_418), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g424 ( .A(n_413), .Y(n_424) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_428), .B2(n_429), .C(n_430), .Y(n_425) );
NAND2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g456 ( .A(n_446), .Y(n_456) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_446), .Y(n_459) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g453 ( .A(n_450), .Y(n_453) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_457), .B(n_461), .C(n_751), .Y(n_460) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g746 ( .A(n_464), .Y(n_746) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_SL g467 ( .A(n_468), .B(n_687), .Y(n_467) );
NAND5xp2_ASAP7_75t_L g468 ( .A(n_469), .B(n_599), .C(n_637), .D(n_658), .E(n_675), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_571), .C(n_592), .Y(n_469) );
OAI221xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_514), .B1(n_538), .B2(n_558), .C(n_562), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_484), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_473), .B(n_560), .Y(n_579) );
OR2x2_ASAP7_75t_L g606 ( .A(n_473), .B(n_497), .Y(n_606) );
AND2x2_ASAP7_75t_L g620 ( .A(n_473), .B(n_497), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_473), .B(n_487), .Y(n_634) );
AND2x2_ASAP7_75t_L g672 ( .A(n_473), .B(n_636), .Y(n_672) );
AND2x2_ASAP7_75t_L g701 ( .A(n_473), .B(n_611), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_473), .B(n_583), .Y(n_718) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g598 ( .A(n_474), .B(n_496), .Y(n_598) );
BUFx3_ASAP7_75t_L g623 ( .A(n_474), .Y(n_623) );
AND2x2_ASAP7_75t_L g652 ( .A(n_474), .B(n_497), .Y(n_652) );
AND3x2_ASAP7_75t_L g665 ( .A(n_474), .B(n_666), .C(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g588 ( .A(n_484), .Y(n_588) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_496), .Y(n_484) );
AOI32xp33_ASAP7_75t_L g643 ( .A1(n_485), .A2(n_595), .A3(n_644), .B1(n_647), .B2(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g570 ( .A(n_486), .B(n_496), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_486), .B(n_598), .Y(n_641) );
AND2x2_ASAP7_75t_L g648 ( .A(n_486), .B(n_620), .Y(n_648) );
OR2x2_ASAP7_75t_L g654 ( .A(n_486), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_486), .B(n_609), .Y(n_679) );
OR2x2_ASAP7_75t_L g697 ( .A(n_486), .B(n_526), .Y(n_697) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g561 ( .A(n_487), .B(n_506), .Y(n_561) );
INVx2_ASAP7_75t_L g583 ( .A(n_487), .Y(n_583) );
OR2x2_ASAP7_75t_L g605 ( .A(n_487), .B(n_506), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_487), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_487), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g666 ( .A(n_487), .B(n_560), .Y(n_666) );
INVx1_ASAP7_75t_SL g717 ( .A(n_496), .Y(n_717) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
INVx1_ASAP7_75t_SL g560 ( .A(n_497), .Y(n_560) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_497), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_497), .B(n_646), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_497), .B(n_583), .C(n_701), .Y(n_712) );
INVx2_ASAP7_75t_L g611 ( .A(n_506), .Y(n_611) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_506), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_525), .Y(n_514) );
INVx1_ASAP7_75t_L g647 ( .A(n_515), .Y(n_647) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g565 ( .A(n_516), .B(n_549), .Y(n_565) );
INVx2_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
AND2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_550), .Y(n_587) );
AND2x2_ASAP7_75t_L g602 ( .A(n_516), .B(n_539), .Y(n_602) );
AND2x2_ASAP7_75t_L g614 ( .A(n_516), .B(n_586), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_525), .B(n_630), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_525), .B(n_587), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_525), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_525), .B(n_581), .Y(n_709) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g548 ( .A(n_526), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_526), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g591 ( .A(n_526), .B(n_539), .Y(n_591) );
AND2x2_ASAP7_75t_L g617 ( .A(n_526), .B(n_549), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_526), .B(n_657), .Y(n_656) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_530), .B(n_537), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_528), .A2(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_537), .Y(n_577) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_548), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_539), .B(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g581 ( .A(n_539), .B(n_582), .Y(n_581) );
INVx3_ASAP7_75t_SL g586 ( .A(n_539), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_539), .B(n_573), .Y(n_639) );
OR2x2_ASAP7_75t_L g649 ( .A(n_539), .B(n_575), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_539), .B(n_617), .Y(n_677) );
OR2x2_ASAP7_75t_L g707 ( .A(n_539), .B(n_549), .Y(n_707) );
AND2x2_ASAP7_75t_L g711 ( .A(n_539), .B(n_550), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_539), .B(n_587), .Y(n_724) );
AND2x2_ASAP7_75t_L g731 ( .A(n_539), .B(n_613), .Y(n_731) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
INVx1_ASAP7_75t_SL g674 ( .A(n_548), .Y(n_674) );
AND2x2_ASAP7_75t_L g613 ( .A(n_549), .B(n_575), .Y(n_613) );
AND2x2_ASAP7_75t_L g627 ( .A(n_549), .B(n_582), .Y(n_627) );
AND2x2_ASAP7_75t_L g630 ( .A(n_549), .B(n_586), .Y(n_630) );
INVx1_ASAP7_75t_L g657 ( .A(n_549), .Y(n_657) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g569 ( .A(n_550), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_559), .A2(n_605), .B(n_729), .C(n_730), .Y(n_728) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g635 ( .A(n_560), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_561), .B(n_578), .Y(n_593) );
AND2x2_ASAP7_75t_L g619 ( .A(n_561), .B(n_620), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_566), .B(n_570), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_564), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g590 ( .A(n_565), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_565), .B(n_586), .Y(n_631) );
AND2x2_ASAP7_75t_L g722 ( .A(n_565), .B(n_573), .Y(n_722) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g595 ( .A(n_569), .B(n_582), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_569), .B(n_580), .Y(n_596) );
OAI322xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_579), .A3(n_580), .B1(n_583), .B2(n_584), .C1(n_588), .C2(n_589), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
AND2x2_ASAP7_75t_L g683 ( .A(n_573), .B(n_595), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_573), .B(n_647), .Y(n_729) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g626 ( .A(n_575), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g692 ( .A(n_579), .B(n_605), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_580), .B(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_581), .B(n_613), .Y(n_670) );
AND2x2_ASAP7_75t_L g616 ( .A(n_582), .B(n_586), .Y(n_616) );
AND2x2_ASAP7_75t_L g624 ( .A(n_583), .B(n_625), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g721 ( .A1(n_583), .A2(n_662), .B(n_722), .C(n_723), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_584), .A2(n_597), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_586), .B(n_613), .Y(n_653) );
AND2x2_ASAP7_75t_L g659 ( .A(n_586), .B(n_627), .Y(n_659) );
AND2x2_ASAP7_75t_L g693 ( .A(n_586), .B(n_595), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_587), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g703 ( .A(n_587), .Y(n_703) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_591), .A2(n_619), .B1(n_621), .B2(n_626), .Y(n_618) );
OAI22xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_596), .B2(n_597), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_593), .A2(n_629), .B1(n_631), .B2(n_632), .Y(n_628) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_598), .A2(n_700), .B1(n_702), .B2(n_704), .C(n_708), .Y(n_699) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B(n_607), .C(n_628), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OR2x2_ASAP7_75t_L g669 ( .A(n_605), .B(n_622), .Y(n_669) );
INVx1_ASAP7_75t_L g720 ( .A(n_605), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_606), .A2(n_608), .B1(n_612), .B2(n_615), .C(n_618), .Y(n_607) );
INVx2_ASAP7_75t_SL g662 ( .A(n_606), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g727 ( .A(n_609), .Y(n_727) );
AND2x2_ASAP7_75t_L g651 ( .A(n_610), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g636 ( .A(n_611), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g698 ( .A(n_614), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_622), .B(n_724), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g622 ( .A(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g667 ( .A(n_625), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_626), .A2(n_638), .B(n_640), .C(n_642), .Y(n_637) );
INVx1_ASAP7_75t_L g715 ( .A(n_629), .Y(n_715) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_633), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g646 ( .A(n_636), .Y(n_646) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_649), .B1(n_650), .B2(n_653), .C1(n_654), .C2(n_656), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g682 ( .A(n_646), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_649), .B(n_703), .Y(n_702) );
NAND2xp33_ASAP7_75t_SL g680 ( .A(n_650), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g655 ( .A(n_652), .Y(n_655) );
AND2x2_ASAP7_75t_L g719 ( .A(n_652), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g685 ( .A(n_655), .B(n_682), .Y(n_685) );
INVx1_ASAP7_75t_L g714 ( .A(n_656), .Y(n_714) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_663), .C(n_668), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_662), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g713 ( .A1(n_665), .A2(n_693), .A3(n_698), .B1(n_714), .B2(n_715), .C1(n_716), .C2(n_719), .Y(n_713) );
AND2x2_ASAP7_75t_L g700 ( .A(n_666), .B(n_701), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_671), .B2(n_673), .Y(n_668) );
INVxp33_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B1(n_680), .B2(n_683), .C(n_684), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND5xp2_ASAP7_75t_L g687 ( .A(n_688), .B(n_699), .C(n_713), .D(n_721), .E(n_725), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_693), .B(n_694), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp33_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_701), .A2(n_726), .B(n_727), .C(n_728), .Y(n_725) );
AOI31xp33_ASAP7_75t_L g708 ( .A1(n_703), .A2(n_709), .A3(n_710), .B(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g726 ( .A(n_724), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g747 ( .A(n_733), .Y(n_747) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_740), .Y(n_743) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
endmodule