module fake_netlist_6_2557_n_1126 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1126);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1126;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_886;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_852;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_901;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_1060;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_816;
wire n_743;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_46),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_6),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_144),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_59),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_93),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_58),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_113),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_44),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_130),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_140),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_47),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_30),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_23),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_71),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_87),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_173),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_5),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_38),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_194),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_35),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_204),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_111),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_68),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_5),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_165),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_2),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_105),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_167),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_21),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_170),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_99),
.Y(n_260)
);

BUFx8_ASAP7_75t_SL g261 ( 
.A(n_52),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_158),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_106),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_27),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_23),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_122),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_16),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_4),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_70),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_129),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_120),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_123),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_41),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_159),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_79),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_25),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_69),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_107),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_53),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_202),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_49),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_231),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_271),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_269),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_231),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_218),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_228),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_266),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_272),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_270),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_235),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_239),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_215),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_261),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_261),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_217),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_220),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_221),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_232),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_225),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_248),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_299),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_226),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_314),
.Y(n_340)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_233),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_227),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_229),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_276),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_288),
.A2(n_248),
.B1(n_249),
.B2(n_279),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_230),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_295),
.B(n_249),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_298),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_304),
.A2(n_255),
.B1(n_280),
.B2(n_277),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_236),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

AOI22x1_ASAP7_75t_SL g360 ( 
.A1(n_289),
.A2(n_283),
.B1(n_264),
.B2(n_263),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_304),
.A2(n_262),
.B1(n_260),
.B2(n_259),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_298),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_295),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_286),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_328),
.B(n_257),
.Y(n_372)
);

OA21x2_ASAP7_75t_L g373 ( 
.A1(n_290),
.A2(n_243),
.B(n_240),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_294),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_329),
.B(n_244),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_327),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_331),
.B(n_253),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_296),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_302),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_287),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_245),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_284),
.B(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_284),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_375),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_386),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_386),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_383),
.Y(n_396)
);

NAND2x1_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_24),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_R g398 ( 
.A(n_368),
.B(n_325),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_383),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_384),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_383),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_383),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_368),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_380),
.Y(n_410)
);

AO21x2_ASAP7_75t_L g411 ( 
.A1(n_337),
.A2(n_326),
.B(n_308),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_354),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_325),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_387),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_381),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_381),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_336),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_336),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_354),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_385),
.B(n_305),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_350),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_349),
.B(n_305),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_381),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_R g433 ( 
.A(n_389),
.B(n_330),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_381),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_382),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_382),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_382),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_382),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_357),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_361),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_336),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_365),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_R g446 ( 
.A(n_373),
.B(n_308),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_349),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_355),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_372),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_356),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_339),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_359),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_379),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_R g457 ( 
.A(n_378),
.B(n_330),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_377),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_377),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_377),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_378),
.B(n_334),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_359),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_347),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_347),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_347),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_446),
.A2(n_420),
.B1(n_463),
.B2(n_456),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_401),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_449),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_402),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_341),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_398),
.B(n_334),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_419),
.B(n_373),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_425),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_412),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_440),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_373),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_434),
.B(n_353),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_453),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_409),
.B(n_342),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_342),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_353),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

AO21x2_ASAP7_75t_L g494 ( 
.A1(n_418),
.A2(n_342),
.B(n_353),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_429),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_457),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_438),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_424),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_390),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_439),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_399),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_396),
.B(n_358),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_413),
.B(n_416),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_L g513 ( 
.A(n_400),
.B(n_358),
.C(n_370),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_405),
.B(n_358),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_441),
.A2(n_378),
.B1(n_250),
.B2(n_251),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_421),
.B(n_378),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_430),
.B(n_363),
.Y(n_517)
);

INVx8_ASAP7_75t_L g518 ( 
.A(n_458),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_411),
.B(n_370),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_431),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_392),
.B(n_370),
.Y(n_522)
);

BUFx8_ASAP7_75t_SL g523 ( 
.A(n_403),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_457),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_411),
.B(n_289),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_421),
.B(n_363),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_291),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_364),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_454),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_443),
.B(n_378),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_397),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_428),
.A2(n_447),
.B1(n_442),
.B2(n_367),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_427),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_395),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_426),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_461),
.B(n_335),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_406),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_461),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_427),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_398),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_433),
.B(n_291),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_335),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_482),
.B(n_364),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

OR2x6_ASAP7_75t_SL g548 ( 
.A(n_464),
.B(n_366),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_502),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_L g550 ( 
.A(n_513),
.B(n_346),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_468),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_340),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_510),
.B(n_366),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_482),
.B(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_469),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_502),
.B(n_367),
.C(n_369),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_470),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_369),
.Y(n_558)
);

NOR2x1_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_346),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_517),
.Y(n_560)
);

NAND2x1p5_ASAP7_75t_L g561 ( 
.A(n_470),
.B(n_339),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_533),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_514),
.B(n_344),
.Y(n_563)
);

A2O1A1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_513),
.A2(n_345),
.B(n_343),
.C(n_338),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_490),
.B(n_338),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_522),
.B(n_343),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_464),
.B(n_0),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_514),
.B(n_26),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_471),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_545),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_477),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_28),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_465),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_478),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_466),
.B(n_541),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_481),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_537),
.B(n_3),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_483),
.B(n_29),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_512),
.B(n_31),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_495),
.B(n_7),
.Y(n_590)
);

NOR2x1_ASAP7_75t_L g591 ( 
.A(n_483),
.B(n_32),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_473),
.Y(n_593)
);

OAI221xp5_ASAP7_75t_L g594 ( 
.A1(n_487),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_499),
.B(n_8),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_521),
.Y(n_597)
);

NAND2x1p5_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_33),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_542),
.B(n_34),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_519),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_600)
);

NAND2x1p5_ASAP7_75t_L g601 ( 
.A(n_542),
.B(n_36),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_480),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_484),
.Y(n_603)
);

OR2x2_ASAP7_75t_SL g604 ( 
.A(n_544),
.B(n_11),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_480),
.Y(n_605)
);

OAI221xp5_ASAP7_75t_L g606 ( 
.A1(n_487),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_495),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_529),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_512),
.B(n_37),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_505),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_576),
.A2(n_491),
.B(n_505),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_562),
.B(n_542),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_576),
.A2(n_491),
.B(n_485),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_571),
.B(n_525),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_589),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_583),
.B(n_512),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_467),
.Y(n_617)
);

BUFx4f_ASAP7_75t_L g618 ( 
.A(n_586),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_554),
.B(n_499),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_593),
.A2(n_485),
.B(n_477),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_593),
.A2(n_538),
.B(n_532),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_543),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_587),
.A2(n_538),
.B(n_516),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_568),
.A2(n_474),
.B(n_536),
.C(n_515),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_602),
.A2(n_498),
.B1(n_524),
.B2(n_501),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_587),
.A2(n_516),
.B(n_494),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_500),
.Y(n_627)
);

O2A1O1Ixp5_ASAP7_75t_L g628 ( 
.A1(n_609),
.A2(n_531),
.B(n_506),
.C(n_530),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_546),
.B(n_527),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_609),
.A2(n_610),
.B(n_605),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_603),
.B(n_534),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_557),
.Y(n_632)
);

BUFx4f_ASAP7_75t_L g633 ( 
.A(n_586),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_548),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_556),
.A2(n_512),
.B(n_474),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_547),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_565),
.B(n_501),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_566),
.B(n_508),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_561),
.A2(n_494),
.B(n_531),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_551),
.B(n_508),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_557),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_524),
.B1(n_498),
.B2(n_540),
.Y(n_642)
);

O2A1O1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_595),
.A2(n_528),
.B(n_535),
.C(n_539),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_570),
.B(n_528),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_572),
.B(n_492),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_590),
.B(n_507),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_561),
.A2(n_504),
.B(n_497),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_556),
.A2(n_504),
.B(n_497),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_550),
.A2(n_506),
.B(n_526),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_574),
.B(n_526),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_569),
.A2(n_475),
.B1(n_526),
.B2(n_518),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_560),
.A2(n_518),
.B(n_526),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_567),
.B(n_518),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_599),
.A2(n_539),
.B(n_40),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_567),
.A2(n_42),
.B(n_39),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_567),
.A2(n_523),
.B1(n_127),
.B2(n_128),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_577),
.B(n_13),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_578),
.B(n_14),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_592),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_597),
.B(n_15),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_582),
.B(n_16),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_550),
.A2(n_132),
.B(n_212),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_569),
.A2(n_131),
.B(n_211),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_604),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_596),
.Y(n_666)
);

NOR2x1_ASAP7_75t_L g667 ( 
.A(n_591),
.B(n_48),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_553),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_579),
.B(n_17),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_608),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_564),
.A2(n_126),
.B(n_210),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_585),
.B(n_17),
.Y(n_672)
);

OAI21xp33_ASAP7_75t_L g673 ( 
.A1(n_575),
.A2(n_18),
.B(n_19),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_553),
.B(n_18),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_563),
.A2(n_134),
.B(n_209),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_627),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_629),
.A2(n_580),
.B(n_581),
.C(n_584),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_614),
.B(n_558),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_617),
.A2(n_558),
.B1(n_563),
.B2(n_562),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_615),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_622),
.B(n_552),
.Y(n_681)
);

O2A1O1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_624),
.A2(n_643),
.B(n_612),
.C(n_642),
.Y(n_682)
);

BUFx4f_ASAP7_75t_L g683 ( 
.A(n_646),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_660),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_637),
.B(n_559),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_SL g686 ( 
.A(n_634),
.B(n_606),
.C(n_594),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_613),
.A2(n_611),
.B(n_623),
.Y(n_688)
);

AOI21x1_ASAP7_75t_L g689 ( 
.A1(n_639),
.A2(n_549),
.B(n_600),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_645),
.B(n_549),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_638),
.B(n_598),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_632),
.Y(n_692)
);

CKINVDCx6p67_ASAP7_75t_R g693 ( 
.A(n_668),
.Y(n_693)
);

OAI22x1_ASAP7_75t_L g694 ( 
.A1(n_612),
.A2(n_600),
.B1(n_601),
.B2(n_598),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_640),
.B(n_601),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_631),
.B(n_625),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_671),
.A2(n_606),
.B(n_594),
.C(n_21),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_666),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_644),
.B(n_19),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_620),
.A2(n_135),
.B(n_208),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_654),
.B(n_618),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_633),
.B(n_20),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_668),
.B(n_20),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_665),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_633),
.A2(n_22),
.B1(n_50),
.B2(n_51),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_670),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_632),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_651),
.B(n_22),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_619),
.B(n_213),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

NOR3xp33_ASAP7_75t_L g711 ( 
.A(n_673),
.B(n_54),
.C(n_55),
.Y(n_711)
);

AOI21x1_ASAP7_75t_L g712 ( 
.A1(n_626),
.A2(n_56),
.B(n_57),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_641),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_653),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_653),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_672),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_658),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_616),
.B(n_207),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_630),
.A2(n_64),
.B(n_65),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_663),
.A2(n_66),
.B(n_67),
.C(n_72),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_636),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_669),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_674),
.Y(n_723)
);

BUFx8_ASAP7_75t_L g724 ( 
.A(n_657),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_659),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_661),
.B(n_73),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_662),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_650),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_635),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_621),
.A2(n_78),
.B(n_80),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_655),
.B(n_81),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_SL g732 ( 
.A(n_648),
.B(n_82),
.Y(n_732)
);

BUFx6f_ASAP7_75t_SL g733 ( 
.A(n_667),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_664),
.B(n_206),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_652),
.B(n_83),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_675),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_736)
);

BUFx12f_ASAP7_75t_L g737 ( 
.A(n_704),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_676),
.Y(n_738)
);

BUFx8_ASAP7_75t_L g739 ( 
.A(n_680),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_683),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_683),
.Y(n_742)
);

BUFx2_ASAP7_75t_SL g743 ( 
.A(n_687),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_687),
.Y(n_744)
);

INVx5_ASAP7_75t_L g745 ( 
.A(n_687),
.Y(n_745)
);

BUFx2_ASAP7_75t_SL g746 ( 
.A(n_733),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_693),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_728),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_692),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_707),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

INVx5_ASAP7_75t_L g752 ( 
.A(n_728),
.Y(n_752)
);

CKINVDCx11_ASAP7_75t_R g753 ( 
.A(n_710),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_698),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_716),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_715),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_656),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_713),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_728),
.B(n_647),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_714),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_696),
.B(n_649),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_715),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_733),
.Y(n_763)
);

BUFx12f_ASAP7_75t_L g764 ( 
.A(n_724),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_724),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_706),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_721),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_679),
.B(n_88),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_681),
.Y(n_769)
);

INVx6_ASAP7_75t_L g770 ( 
.A(n_726),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_727),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_709),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_723),
.B(n_89),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_722),
.B(n_90),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_725),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_703),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_677),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_689),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_699),
.Y(n_779)
);

NAND2x1p5_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_628),
.Y(n_780)
);

INVx3_ASAP7_75t_SL g781 ( 
.A(n_702),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_735),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_690),
.B(n_91),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_694),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_691),
.B(n_92),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_682),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_712),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_688),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_695),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_701),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_708),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_732),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_686),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_731),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_718),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_700),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_734),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_705),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_719),
.Y(n_799)
);

BUFx12f_ASAP7_75t_L g800 ( 
.A(n_717),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_697),
.B(n_94),
.Y(n_801)
);

BUFx12f_ASAP7_75t_L g802 ( 
.A(n_736),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_787),
.A2(n_730),
.B(n_729),
.Y(n_803)
);

OAI21xp33_ASAP7_75t_L g804 ( 
.A1(n_801),
.A2(n_711),
.B(n_720),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_793),
.B(n_769),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_778),
.A2(n_95),
.B(n_96),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_739),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_778),
.A2(n_97),
.B(n_98),
.Y(n_808)
);

AO21x2_ASAP7_75t_L g809 ( 
.A1(n_788),
.A2(n_100),
.B(n_101),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_764),
.Y(n_810)
);

OA21x2_ASAP7_75t_L g811 ( 
.A1(n_788),
.A2(n_102),
.B(n_104),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_750),
.B(n_108),
.Y(n_812)
);

CKINVDCx6p67_ASAP7_75t_R g813 ( 
.A(n_745),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_801),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_775),
.B(n_114),
.Y(n_815)
);

AO21x1_ASAP7_75t_L g816 ( 
.A1(n_761),
.A2(n_115),
.B(n_116),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_781),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_769),
.B(n_121),
.Y(n_818)
);

AOI221xp5_ASAP7_75t_L g819 ( 
.A1(n_761),
.A2(n_779),
.B1(n_795),
.B2(n_786),
.C(n_783),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_759),
.A2(n_124),
.B(n_125),
.Y(n_820)
);

AND2x2_ASAP7_75t_SL g821 ( 
.A(n_797),
.B(n_136),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_759),
.A2(n_137),
.B(n_139),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_SL g823 ( 
.A1(n_785),
.A2(n_141),
.B(n_143),
.C(n_145),
.Y(n_823)
);

NOR4xp25_ASAP7_75t_L g824 ( 
.A(n_768),
.B(n_146),
.C(n_148),
.D(n_149),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_783),
.A2(n_150),
.B(n_153),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_780),
.A2(n_154),
.B(n_155),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_784),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_780),
.A2(n_156),
.B(n_157),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_799),
.A2(n_160),
.B(n_161),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_741),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_754),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_762),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_789),
.B(n_162),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_798),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_834)
);

AO31x2_ASAP7_75t_L g835 ( 
.A1(n_777),
.A2(n_168),
.A3(n_169),
.B(n_171),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_766),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_762),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_785),
.A2(n_172),
.B(n_174),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_771),
.B(n_175),
.Y(n_839)
);

OAI221xp5_ASAP7_75t_L g840 ( 
.A1(n_776),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.C(n_179),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_775),
.Y(n_841)
);

CKINVDCx6p67_ASAP7_75t_R g842 ( 
.A(n_745),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_767),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_799),
.A2(n_180),
.B(n_181),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_738),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_767),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_774),
.A2(n_182),
.B(n_183),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_769),
.B(n_185),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_774),
.A2(n_186),
.B(n_187),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_781),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_740),
.Y(n_851)
);

A2O1A1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_798),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_749),
.A2(n_195),
.B(n_197),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_749),
.A2(n_198),
.B(n_199),
.Y(n_854)
);

AO21x2_ASAP7_75t_L g855 ( 
.A1(n_757),
.A2(n_201),
.B(n_203),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_782),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_758),
.A2(n_205),
.B(n_773),
.Y(n_857)
);

AOI21x1_ASAP7_75t_SL g858 ( 
.A1(n_800),
.A2(n_746),
.B(n_802),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_782),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_797),
.B(n_794),
.Y(n_860)
);

NAND2x1_ASAP7_75t_L g861 ( 
.A(n_794),
.B(n_797),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_756),
.A2(n_763),
.B(n_796),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_756),
.A2(n_763),
.B(n_796),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_767),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_831),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_810),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_862),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_841),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_856),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_827),
.B(n_772),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_836),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_827),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_856),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_859),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_860),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_803),
.A2(n_792),
.B(n_794),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_830),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_863),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_835),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_864),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_864),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_843),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_819),
.B(n_738),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_861),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_846),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_835),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_845),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_804),
.A2(n_772),
.B1(n_791),
.B2(n_792),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_860),
.B(n_791),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_805),
.B(n_770),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_826),
.A2(n_792),
.B(n_770),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_811),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_811),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_847),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_860),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_860),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_815),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_809),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_832),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_828),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_806),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_808),
.A2(n_792),
.B(n_770),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_849),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_832),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_820),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_838),
.Y(n_906)
);

INVx11_ASAP7_75t_L g907 ( 
.A(n_810),
.Y(n_907)
);

AO21x1_ASAP7_75t_L g908 ( 
.A1(n_825),
.A2(n_751),
.B(n_752),
.Y(n_908)
);

OAI21x1_ASAP7_75t_SL g909 ( 
.A1(n_857),
.A2(n_751),
.B(n_755),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_822),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_853),
.A2(n_748),
.B(n_752),
.Y(n_911)
);

BUFx8_ASAP7_75t_SL g912 ( 
.A(n_866),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_868),
.B(n_807),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_866),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_883),
.A2(n_814),
.B1(n_888),
.B2(n_821),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_872),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_876),
.A2(n_854),
.B(n_858),
.Y(n_917)
);

BUFx4f_ASAP7_75t_SL g918 ( 
.A(n_875),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_887),
.B(n_824),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_908),
.A2(n_816),
.B1(n_840),
.B2(n_848),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_872),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_865),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_865),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_R g924 ( 
.A(n_875),
.B(n_753),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_SL g925 ( 
.A(n_889),
.B(n_818),
.C(n_850),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_907),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_871),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_907),
.Y(n_928)
);

CKINVDCx11_ASAP7_75t_R g929 ( 
.A(n_897),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_SL g930 ( 
.A(n_903),
.B(n_817),
.C(n_852),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_896),
.A2(n_834),
.B1(n_765),
.B2(n_790),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_869),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_890),
.B(n_737),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_890),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_908),
.B(n_876),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_871),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_878),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_881),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_870),
.B(n_837),
.Y(n_939)
);

CKINVDCx16_ASAP7_75t_R g940 ( 
.A(n_870),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_900),
.A2(n_855),
.B1(n_844),
.B2(n_829),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_884),
.B(n_753),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_R g943 ( 
.A(n_884),
.B(n_765),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_877),
.B(n_837),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_874),
.B(n_760),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_877),
.B(n_760),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_940),
.B(n_867),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_929),
.B(n_884),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_916),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_915),
.A2(n_920),
.B1(n_919),
.B2(n_931),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_932),
.B(n_867),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_937),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_921),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_922),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_932),
.B(n_935),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_935),
.B(n_867),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_935),
.B(n_878),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_943),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_923),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_927),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_936),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_938),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_944),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_945),
.Y(n_965)
);

CKINVDCx6p67_ASAP7_75t_R g966 ( 
.A(n_912),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_939),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_946),
.B(n_881),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_913),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_914),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_934),
.B(n_874),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_917),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_965),
.B(n_873),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_873),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_953),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_970),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_954),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_948),
.B(n_933),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_951),
.A2(n_941),
.B(n_823),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_954),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_947),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_955),
.Y(n_982)
);

INVx5_ASAP7_75t_L g983 ( 
.A(n_970),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_948),
.B(n_942),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_972),
.A2(n_893),
.B(n_892),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_955),
.Y(n_986)
);

OAI22xp33_ASAP7_75t_L g987 ( 
.A1(n_959),
.A2(n_918),
.B1(n_898),
.B2(n_903),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_972),
.A2(n_898),
.B(n_909),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_961),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_973),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_959),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_983),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_974),
.B(n_967),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_975),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_983),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_982),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_983),
.B(n_978),
.Y(n_997)
);

AOI221xp5_ASAP7_75t_L g998 ( 
.A1(n_979),
.A2(n_964),
.B1(n_956),
.B2(n_958),
.C(n_969),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_977),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_983),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_980),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_986),
.B(n_964),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_1000),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_991),
.B(n_966),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_997),
.B(n_976),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_997),
.B(n_966),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_992),
.B(n_956),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_996),
.B(n_975),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_992),
.B(n_949),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_979),
.C(n_995),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1003),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1011),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1004),
.B(n_999),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_1005),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1016),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_1007),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_1017),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1018),
.B(n_1006),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1014),
.B(n_1016),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1013),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1012),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1016),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1015),
.B(n_1009),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_1015),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_1021),
.B(n_995),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1020),
.B(n_1008),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_1028),
.B(n_928),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1022),
.B(n_990),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_1025),
.B(n_998),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_993),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1027),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_1024),
.B(n_926),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1030),
.B(n_1019),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1034),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_1031),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1032),
.B(n_1026),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1036),
.B(n_1023),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1033),
.A2(n_1029),
.B1(n_1031),
.B2(n_1023),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1040),
.B(n_1001),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1038),
.B(n_1001),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1042),
.B(n_1002),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1037),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1041),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_1047),
.B(n_1039),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1048),
.B(n_1043),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_1044),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_1045),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1046),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_1048),
.B(n_747),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_L g1055 ( 
.A(n_1054),
.B(n_747),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_1051),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_L g1057 ( 
.A(n_1050),
.B(n_987),
.C(n_790),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1053),
.B(n_981),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_1052),
.B(n_987),
.C(n_833),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1049),
.A2(n_981),
.B1(n_918),
.B2(n_957),
.Y(n_1060)
);

OAI211xp5_ASAP7_75t_SL g1061 ( 
.A1(n_1056),
.A2(n_930),
.B(n_925),
.C(n_839),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1055),
.A2(n_988),
.B(n_930),
.C(n_957),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_1058),
.B(n_739),
.Y(n_1063)
);

NAND5xp2_ASAP7_75t_L g1064 ( 
.A(n_1057),
.B(n_925),
.C(n_924),
.D(n_988),
.E(n_958),
.Y(n_1064)
);

AOI211xp5_ASAP7_75t_L g1065 ( 
.A1(n_1060),
.A2(n_747),
.B(n_812),
.C(n_740),
.Y(n_1065)
);

XNOR2x1_ASAP7_75t_L g1066 ( 
.A(n_1063),
.B(n_812),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1064),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1062),
.A2(n_1059),
.B(n_989),
.Y(n_1069)
);

AO22x2_ASAP7_75t_L g1070 ( 
.A1(n_1061),
.A2(n_743),
.B1(n_953),
.B2(n_947),
.Y(n_1070)
);

NAND4xp25_ASAP7_75t_L g1071 ( 
.A(n_1065),
.B(n_750),
.C(n_971),
.D(n_952),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1063),
.B(n_745),
.Y(n_1072)
);

OAI211xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1065),
.A2(n_968),
.B(n_906),
.C(n_894),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

NAND3x1_ASAP7_75t_SL g1075 ( 
.A(n_1067),
.B(n_971),
.C(n_842),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_1072),
.B(n_744),
.C(n_745),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1069),
.A2(n_952),
.B(n_985),
.C(n_744),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_1066),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1070),
.B(n_882),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1070),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1071),
.B(n_885),
.Y(n_1081)
);

NOR2x1_ASAP7_75t_L g1082 ( 
.A(n_1073),
.B(n_740),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_960),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_L g1084 ( 
.A(n_1080),
.B(n_744),
.C(n_742),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1078),
.B(n_962),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1076),
.B(n_742),
.Y(n_1086)
);

NAND5xp2_ASAP7_75t_L g1087 ( 
.A(n_1077),
.B(n_742),
.C(n_900),
.D(n_813),
.E(n_901),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1081),
.B(n_851),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1079),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1082),
.B(n_950),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_1075),
.B(n_906),
.C(n_894),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1080),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1080),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1078),
.B(n_851),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_1074),
.B(n_851),
.C(n_762),
.Y(n_1095)
);

AND3x1_ASAP7_75t_L g1096 ( 
.A(n_1092),
.B(n_895),
.C(n_961),
.Y(n_1096)
);

NAND4xp25_ASAP7_75t_L g1097 ( 
.A(n_1084),
.B(n_880),
.C(n_905),
.D(n_901),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_1093),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1094),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1089),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1083),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_1085),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_1088),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1086),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1098),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_1102),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_SL g1107 ( 
.A1(n_1100),
.A2(n_1095),
.B1(n_1090),
.B2(n_1091),
.Y(n_1107)
);

XNOR2xp5_ASAP7_75t_L g1108 ( 
.A(n_1103),
.B(n_1101),
.Y(n_1108)
);

AOI22x1_ASAP7_75t_L g1109 ( 
.A1(n_1104),
.A2(n_1087),
.B1(n_909),
.B2(n_895),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1099),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_L g1111 ( 
.A(n_1110),
.B(n_1097),
.C(n_1096),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1105),
.B(n_899),
.Y(n_1112)
);

AO21x2_ASAP7_75t_L g1113 ( 
.A1(n_1108),
.A2(n_911),
.B(n_891),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

XNOR2xp5_ASAP7_75t_L g1115 ( 
.A(n_1114),
.B(n_1106),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1115),
.Y(n_1116)
);

OR3x2_ASAP7_75t_L g1117 ( 
.A(n_1116),
.B(n_1107),
.C(n_1111),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1116),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_1109),
.B1(n_1113),
.B2(n_963),
.Y(n_1119)
);

O2A1O1Ixp5_ASAP7_75t_L g1120 ( 
.A1(n_1118),
.A2(n_963),
.B(n_905),
.C(n_886),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1119),
.A2(n_899),
.B1(n_748),
.B2(n_752),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1120),
.A2(n_905),
.B1(n_910),
.B2(n_886),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_911),
.B(n_891),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_902),
.B(n_904),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1124),
.A2(n_748),
.B(n_752),
.Y(n_1125)
);

AOI211xp5_ASAP7_75t_L g1126 ( 
.A1(n_1125),
.A2(n_1123),
.B(n_902),
.C(n_879),
.Y(n_1126)
);


endmodule