module fake_jpeg_15071_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_33),
.Y(n_58)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_47),
.B1(n_49),
.B2(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_29),
.B1(n_36),
.B2(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_56),
.B1(n_22),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_60),
.A3(n_49),
.B1(n_51),
.B2(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_22),
.B1(n_20),
.B2(n_0),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_30),
.B(n_28),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_63),
.B(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_65),
.B1(n_84),
.B2(n_61),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_29),
.B(n_28),
.C(n_30),
.Y(n_66)
);

FAx1_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_36),
.CI(n_35),
.CON(n_67),
.SN(n_67)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_33),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_37),
.C(n_30),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_71),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_76),
.Y(n_109)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_17),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_58),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_0),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_81),
.Y(n_87)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_46),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_102),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_87),
.B1(n_102),
.B2(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_97),
.Y(n_112)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_58),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_107),
.B1(n_81),
.B2(n_65),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_37),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_71),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_12),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_133),
.B1(n_44),
.B2(n_59),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_118),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_84),
.B(n_79),
.C(n_71),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_109),
.B(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_74),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_81),
.B(n_76),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_125),
.B(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_132),
.B1(n_90),
.B2(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_83),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_71),
.B1(n_66),
.B2(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_68),
.B1(n_82),
.B2(n_75),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_44),
.B1(n_59),
.B2(n_33),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_100),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_146),
.C(n_128),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_107),
.A3(n_96),
.B1(n_91),
.B2(n_109),
.C1(n_101),
.C2(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_152),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_101),
.B1(n_96),
.B2(n_105),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_113),
.B1(n_116),
.B2(n_133),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_149),
.B(n_153),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_37),
.C(n_46),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_147),
.A2(n_112),
.B1(n_116),
.B2(n_127),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_28),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_94),
.B(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_17),
.B(n_97),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_110),
.B1(n_125),
.B2(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_166),
.C(n_170),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_110),
.B1(n_126),
.B2(n_98),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_116),
.B1(n_124),
.B2(n_120),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_116),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_116),
.B1(n_131),
.B2(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_178),
.B1(n_155),
.B2(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_30),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_46),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_28),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_146),
.C(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_98),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_138),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_185),
.B1(n_188),
.B2(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_144),
.C(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_192),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_140),
.B1(n_135),
.B2(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_135),
.C(n_150),
.Y(n_190)
);

OAI21x1_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_178),
.B(n_174),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_141),
.B1(n_151),
.B2(n_6),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_172),
.C(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_164),
.B1(n_171),
.B2(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_198),
.B1(n_209),
.B2(n_201),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_173),
.B1(n_160),
.B2(n_175),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_208),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_213),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_199),
.A2(n_178),
.B1(n_181),
.B2(n_183),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_198),
.B(n_197),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_181),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_186),
.B1(n_192),
.B2(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_5),
.C(n_6),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_6),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_225),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_215),
.B(n_212),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_205),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_206),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_230),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_227),
.B(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_222),
.C(n_224),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_234),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_196),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_203),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_238),
.A3(n_213),
.B1(n_222),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_215),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_235),
.B(n_8),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_14),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_7),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_244),
.B(n_10),
.Y(n_245)
);

AOI32xp33_ASAP7_75t_L g246 ( 
.A1(n_245),
.A2(n_242),
.A3(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_15),
.Y(n_247)
);


endmodule