module fake_jpeg_14839_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_63),
.Y(n_68)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_57),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_71),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_52),
.B(n_57),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_58),
.B(n_44),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_76),
.Y(n_96)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_83),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_65),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_99),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_88),
.B1(n_98),
.B2(n_103),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_5),
.B(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_56),
.B1(n_43),
.B2(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_97),
.Y(n_110)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_1),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_42),
.B1(n_49),
.B2(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_1),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_42),
.B1(n_51),
.B2(n_24),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_103),
.B1(n_98),
.B2(n_89),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_51),
.CI(n_6),
.CON(n_105),
.SN(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_115),
.Y(n_116)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_90),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_25),
.B1(n_37),
.B2(n_36),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_8),
.B1(n_105),
.B2(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_96),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_121),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_7),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_94),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_128),
.B1(n_117),
.B2(n_12),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_111),
.B1(n_108),
.B2(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_113),
.B1(n_13),
.B2(n_16),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_133),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_138),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_134),
.B(n_17),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_135),
.C(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_113),
.C(n_20),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_11),
.C(n_21),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_22),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

OAI311xp33_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_29),
.A3(n_30),
.B1(n_31),
.C1(n_32),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_34),
.B(n_35),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_149),
.Y(n_150)
);


endmodule