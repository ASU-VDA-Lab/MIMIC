module fake_jpeg_24103_n_184 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.C(n_1),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_34),
.B1(n_43),
.B2(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_22),
.B1(n_31),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_34),
.B1(n_30),
.B2(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_23),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_43),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_18),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_41),
.B1(n_40),
.B2(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_71),
.B1(n_79),
.B2(n_81),
.Y(n_95)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_57),
.C(n_54),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_43),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_80),
.B(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_36),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_83),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_42),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_42),
.B1(n_20),
.B2(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_0),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_88),
.B(n_90),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_39),
.Y(n_92)
);

OA21x2_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_102),
.B(n_80),
.Y(n_112)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_9),
.Y(n_124)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_37),
.B(n_53),
.C(n_24),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_81),
.B1(n_82),
.B2(n_66),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_24),
.B(n_2),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_68),
.B(n_80),
.C(n_77),
.D(n_73),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_118),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_79),
.B1(n_78),
.B2(n_71),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_112),
.B(n_92),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_68),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_123),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_0),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_2),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_2),
.C(n_4),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_95),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_94),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_143),
.C(n_116),
.Y(n_148)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_97),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_146),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_117),
.C(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_91),
.B(n_96),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_138),
.B(n_144),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_140),
.C(n_136),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_119),
.C(n_111),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_156),
.C(n_93),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_134),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_121),
.C(n_123),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_139),
.B1(n_142),
.B2(n_133),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_129),
.B1(n_145),
.B2(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_154),
.B(n_152),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_134),
.CI(n_135),
.CON(n_162),
.SN(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_166),
.B1(n_164),
.B2(n_162),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_171),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_156),
.B(n_96),
.Y(n_170)
);

HAxp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_162),
.CON(n_175),
.SN(n_175)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_166),
.B1(n_165),
.B2(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_176),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_6),
.B(n_11),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_176)
);

AOI31xp67_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_170),
.A3(n_172),
.B(n_15),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_179),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_173),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_181),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);


endmodule