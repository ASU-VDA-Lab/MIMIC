module fake_jpeg_27491_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_19),
.B1(n_27),
.B2(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_19),
.B1(n_25),
.B2(n_22),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_18),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_66),
.B1(n_70),
.B2(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_22),
.C(n_29),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_43),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_0),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_26),
.B(n_1),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_16),
.B1(n_28),
.B2(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_2),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_0),
.Y(n_110)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_48),
.A3(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_82)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_54),
.B(n_42),
.C(n_45),
.D(n_46),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_90),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_69),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_68),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_44),
.B(n_46),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_71),
.B(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_46),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_110),
.B(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_105),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_108),
.C(n_95),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_54),
.B1(n_42),
.B2(n_75),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_54),
.B1(n_81),
.B2(n_79),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_75),
.B(n_68),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_109),
.B(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_88),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_45),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_120),
.B(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_98),
.B1(n_84),
.B2(n_103),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_76),
.C(n_79),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_125),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_86),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_100),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_96),
.B1(n_109),
.B2(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_129),
.A2(n_132),
.B1(n_135),
.B2(n_1),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_112),
.C(n_108),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_137),
.C(n_138),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_112),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_97),
.C(n_80),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_46),
.C(n_77),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_101),
.C(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_140),
.C(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_114),
.B1(n_120),
.B2(n_113),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_127),
.C(n_115),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_150),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_122),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_148),
.B(n_149),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_0),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_13),
.B1(n_10),
.B2(n_3),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_141),
.C(n_151),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_131),
.C(n_10),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_2),
.B(n_3),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_142),
.C(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_146),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_6),
.B(n_7),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_2),
.B(n_4),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_161),
.C(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_165),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_167),
.A2(n_158),
.B(n_8),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_8),
.B(n_170),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_172),
.CI(n_161),
.CON(n_173),
.SN(n_173)
);


endmodule