module fake_jpeg_27874_n_401 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_401);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_39),
.B(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_45),
.Y(n_98)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_50),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_53),
.Y(n_89)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_17),
.B(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_56),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_32),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_17),
.B(n_8),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_17),
.B1(n_36),
.B2(n_34),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_20),
.B(n_30),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_87),
.A2(n_33),
.B(n_62),
.C(n_30),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_26),
.B1(n_38),
.B2(n_36),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_102),
.B1(n_110),
.B2(n_55),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_49),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_38),
.B1(n_29),
.B2(n_36),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_71),
.B1(n_65),
.B2(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_67),
.B1(n_51),
.B2(n_56),
.Y(n_120)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_21),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_29),
.B1(n_34),
.B2(n_37),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_111),
.Y(n_142)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_34),
.B1(n_29),
.B2(n_50),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_118),
.B1(n_149),
.B2(n_152),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_117),
.B(n_122),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_48),
.B1(n_72),
.B2(n_54),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_47),
.B1(n_97),
.B2(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_119),
.A2(n_21),
.B1(n_20),
.B2(n_10),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_143),
.B1(n_92),
.B2(n_84),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_23),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_134),
.B(n_62),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_31),
.B1(n_30),
.B2(n_66),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_98),
.B1(n_86),
.B2(n_79),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_138),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_22),
.B1(n_37),
.B2(n_25),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_78),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_146),
.B(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_42),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_139),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_23),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_44),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_145),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_94),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_31),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_30),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_141),
.A2(n_1),
.B(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_22),
.B1(n_37),
.B2(n_25),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_22),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_96),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_155),
.Y(n_183)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_25),
.B1(n_31),
.B2(n_33),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_81),
.B(n_12),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_98),
.A2(n_33),
.B1(n_11),
.B2(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_109),
.B1(n_75),
.B2(n_82),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_96),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_159),
.A2(n_163),
.B1(n_170),
.B2(n_173),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_160),
.A2(n_182),
.B1(n_142),
.B2(n_121),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_101),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_101),
.B1(n_99),
.B2(n_93),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_93),
.B1(n_30),
.B2(n_33),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_189),
.B1(n_142),
.B2(n_121),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_122),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_0),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_0),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_181),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_178),
.Y(n_201)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_0),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_1),
.B(n_2),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_20),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_130),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_121),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

XOR2x1_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_1),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_196),
.A2(n_200),
.B(n_161),
.Y(n_249)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_225),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_184),
.B(n_166),
.C(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_151),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_205),
.B(n_209),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_134),
.B(n_124),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_206),
.A2(n_214),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_146),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_125),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_222),
.Y(n_252)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_142),
.B1(n_144),
.B2(n_135),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_129),
.B1(n_5),
.B2(n_6),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_167),
.A2(n_151),
.B1(n_155),
.B2(n_147),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_219),
.B1(n_227),
.B2(n_192),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_130),
.C(n_137),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_189),
.C(n_161),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_224),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_221),
.B(n_158),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_140),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_158),
.B(n_11),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_140),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_170),
.A2(n_140),
.B1(n_129),
.B2(n_4),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_2),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

INVxp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_245),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_156),
.B(n_176),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_242),
.B(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_157),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_239),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_171),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_202),
.A2(n_176),
.B(n_193),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_251),
.C(n_264),
.Y(n_276)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_253),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_199),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_248),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_196),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_255),
.B(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_196),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_223),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_201),
.A2(n_162),
.B(n_178),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_199),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

OAI22x1_ASAP7_75t_L g259 ( 
.A1(n_214),
.A2(n_129),
.B1(n_190),
.B2(n_188),
.Y(n_259)
);

OAI22x1_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_232),
.B1(n_227),
.B2(n_216),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_162),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_232),
.B(n_206),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_278),
.B(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_288),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_240),
.B1(n_237),
.B2(n_235),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_207),
.C(n_195),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_284),
.C(n_292),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_236),
.Y(n_283)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_195),
.C(n_197),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_234),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_243),
.B(n_197),
.C(n_222),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_209),
.C(n_212),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_251),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_247),
.A2(n_229),
.B1(n_223),
.B2(n_230),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_294),
.A2(n_215),
.B1(n_216),
.B2(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_249),
.B(n_265),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_302),
.B(n_269),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_316),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_274),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_301),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_245),
.B1(n_255),
.B2(n_263),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_279),
.A2(n_258),
.B1(n_233),
.B2(n_242),
.Y(n_303)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_277),
.B(n_261),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_307),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_282),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_317),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_233),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_267),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_265),
.Y(n_315)
);

XOR2x2_ASAP7_75t_SL g316 ( 
.A(n_289),
.B(n_257),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_271),
.A2(n_260),
.B1(n_266),
.B2(n_5),
.Y(n_318)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_296),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_288),
.Y(n_324)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_292),
.C(n_281),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_327),
.C(n_328),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_284),
.C(n_268),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_268),
.C(n_293),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_291),
.Y(n_329)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_270),
.Y(n_330)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_316),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_295),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_272),
.B(n_280),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_306),
.A2(n_286),
.B(n_283),
.Y(n_338)
);

AOI21xp33_ASAP7_75t_L g353 ( 
.A1(n_338),
.A2(n_286),
.B(n_300),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_323),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_340),
.B(n_342),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_322),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_298),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_346),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_345),
.B(n_332),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_275),
.B(n_299),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_329),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_349),
.B(n_331),
.Y(n_366)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_350),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_353),
.A2(n_337),
.B(n_334),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_326),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_354),
.B(n_324),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_357),
.A2(n_360),
.B(n_362),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_334),
.B1(n_320),
.B2(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_359),
.B(n_364),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_352),
.A2(n_338),
.B(n_321),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_333),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_333),
.Y(n_369)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_305),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_315),
.Y(n_365)
);

OAI21x1_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_336),
.B(n_343),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_366),
.B(n_367),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_325),
.C(n_327),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_330),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_371),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_343),
.B(n_357),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_344),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_351),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_377),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_311),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_376),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_303),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_317),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g387 ( 
.A1(n_379),
.A2(n_348),
.B(n_341),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_384),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_362),
.B(n_360),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_382),
.A2(n_347),
.B(n_348),
.Y(n_391)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_312),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_273),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_300),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_388),
.B(n_390),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_367),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_373),
.Y(n_390)
);

AO21x1_ASAP7_75t_L g393 ( 
.A1(n_391),
.A2(n_392),
.B(n_383),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_395),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_389),
.A2(n_379),
.B1(n_380),
.B2(n_310),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_SL g397 ( 
.A1(n_394),
.A2(n_389),
.B(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_397),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_SL g399 ( 
.A1(n_398),
.A2(n_396),
.B(n_318),
.C(n_273),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_399),
.A2(n_266),
.B(n_336),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_400),
.A2(n_369),
.B(n_371),
.Y(n_401)
);


endmodule