module fake_jpeg_22187_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_218;
wire n_63;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_27),
.B1(n_16),
.B2(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_23),
.B1(n_18),
.B2(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_60),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_54),
.B1(n_38),
.B2(n_43),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_67),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_54),
.B1(n_38),
.B2(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_92),
.B1(n_57),
.B2(n_55),
.Y(n_108)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_46),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_55),
.C(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_46),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_66),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_38),
.B1(n_54),
.B2(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_69),
.B1(n_56),
.B2(n_48),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_101),
.B1(n_117),
.B2(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_71),
.B1(n_61),
.B2(n_58),
.Y(n_100)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_100),
.A2(n_24),
.B(n_25),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_49),
.B1(n_45),
.B2(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_109),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_44),
.B(n_68),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_96),
.B(n_82),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_48),
.B1(n_45),
.B2(n_39),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_89),
.B1(n_80),
.B2(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_53),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_128),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_87),
.B(n_93),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_129),
.B(n_138),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_95),
.B1(n_89),
.B2(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_133),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_96),
.B1(n_56),
.B2(n_87),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_96),
.B1(n_97),
.B2(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_124),
.B1(n_125),
.B2(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_105),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_115),
.B1(n_99),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_163),
.B1(n_29),
.B2(n_30),
.Y(n_183)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_103),
.B1(n_116),
.B2(n_102),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_128),
.B1(n_138),
.B2(n_139),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_29),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_103),
.C(n_113),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_160),
.C(n_164),
.Y(n_181)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_120),
.B1(n_141),
.B2(n_28),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_159),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_28),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_0),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_0),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_113),
.B1(n_119),
.B2(n_81),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_119),
.C(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_161),
.B(n_149),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_122),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_176),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_147),
.B1(n_166),
.B2(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_53),
.B1(n_51),
.B2(n_39),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_185),
.B1(n_158),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_14),
.B1(n_26),
.B2(n_21),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_30),
.C(n_53),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_163),
.C(n_160),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_152),
.B1(n_158),
.B2(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_189),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_145),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_144),
.B(n_25),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_25),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_148),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_198),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_148),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_209),
.C(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_206),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_204),
.B1(n_208),
.B2(n_199),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_187),
.B1(n_174),
.B2(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_210),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_161),
.B1(n_154),
.B2(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_178),
.C(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_183),
.Y(n_220)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_215),
.C(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_178),
.C(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_223),
.B(n_230),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_224),
.B1(n_21),
.B2(n_19),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_201),
.C(n_193),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_184),
.C(n_182),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_228),
.C(n_26),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_211),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_172),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_12),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_175),
.B1(n_174),
.B2(n_63),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_227),
.B(n_1),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_63),
.C(n_51),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_220),
.B1(n_219),
.B2(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_198),
.B1(n_194),
.B2(n_196),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_237),
.B(n_238),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_51),
.B1(n_39),
.B2(n_26),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_21),
.B1(n_19),
.B2(n_3),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_5),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_19),
.B1(n_2),
.B2(n_4),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_245),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_11),
.B1(n_2),
.B2(n_4),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_6),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_232),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_250),
.B(n_235),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_214),
.B(n_5),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_1),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_5),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_257),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_6),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_7),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_262),
.B(n_264),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_261),
.B(n_265),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_233),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_243),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_6),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_24),
.B1(n_8),
.B2(n_10),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_269),
.C(n_255),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_7),
.B(n_8),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_276),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_255),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_256),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_279),
.B(n_280),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_24),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_270),
.B(n_277),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_283),
.B1(n_282),
.B2(n_24),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_7),
.B(n_8),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_10),
.B(n_7),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_8),
.C(n_10),
.Y(n_289)
);


endmodule