module fake_jpeg_30853_n_534 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_18),
.B(n_0),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_76),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_2),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx12f_ASAP7_75t_SL g89 ( 
.A(n_44),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g148 ( 
.A(n_89),
.B(n_93),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_101),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_104),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_44),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_44),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_51),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_110),
.B(n_120),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_87),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_128),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_50),
.C(n_47),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_46),
.C(n_43),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_43),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_35),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_42),
.B1(n_20),
.B2(n_17),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_132),
.B1(n_157),
.B2(n_104),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_127),
.A2(n_153),
.B1(n_160),
.B2(n_27),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_30),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_33),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_34),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_20),
.B1(n_17),
.B2(n_42),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_34),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_96),
.A2(n_38),
.B1(n_50),
.B2(n_47),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_86),
.A2(n_17),
.B1(n_42),
.B2(n_20),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_55),
.A2(n_58),
.B1(n_91),
.B2(n_90),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_85),
.B(n_38),
.Y(n_162)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_181),
.Y(n_227)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_174),
.A2(n_184),
.B1(n_166),
.B2(n_25),
.Y(n_225)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_177),
.Y(n_260)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_84),
.Y(n_181)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_191),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_105),
.A2(n_85),
.B1(n_42),
.B2(n_20),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_199),
.B1(n_211),
.B2(n_154),
.Y(n_222)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_190),
.Y(n_264)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_31),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_192),
.B(n_196),
.Y(n_252)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_106),
.B(n_155),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_31),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_118),
.B(n_46),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_198),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_25),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_105),
.A2(n_20),
.B1(n_42),
.B2(n_83),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_148),
.A2(n_52),
.B(n_29),
.C(n_27),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_161),
.Y(n_223)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_206),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_52),
.B(n_29),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_212),
.C(n_159),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_113),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_209),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_137),
.A2(n_68),
.B1(n_66),
.B2(n_64),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_214),
.B1(n_154),
.B2(n_137),
.Y(n_232)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_215),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_133),
.B(n_52),
.C(n_29),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_213),
.A2(n_164),
.B1(n_122),
.B2(n_39),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_132),
.A2(n_157),
.B1(n_119),
.B2(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_27),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_220),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_115),
.A2(n_25),
.B1(n_98),
.B2(n_39),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_121),
.B1(n_149),
.B2(n_125),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_140),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_136),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_234),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_184),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_23),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_232),
.A2(n_233),
.B1(n_262),
.B2(n_263),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_138),
.B1(n_136),
.B2(n_115),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_39),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_170),
.B(n_146),
.C(n_138),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_214),
.C(n_212),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_245),
.A2(n_261),
.B1(n_39),
.B2(n_23),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_185),
.B(n_172),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_190),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_214),
.A2(n_122),
.B1(n_121),
.B2(n_125),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_213),
.A2(n_164),
.B1(n_149),
.B2(n_111),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_265),
.B(n_287),
.Y(n_324)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_271),
.C(n_296),
.Y(n_302)
);

AOI22x1_ASAP7_75t_SL g269 ( 
.A1(n_223),
.A2(n_181),
.B1(n_201),
.B2(n_179),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_243),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_270),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_182),
.Y(n_271)
);

BUFx6f_ASAP7_75t_SL g272 ( 
.A(n_249),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_227),
.A2(n_202),
.B(n_180),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_273),
.A2(n_278),
.B(n_284),
.Y(n_334)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_169),
.B1(n_183),
.B2(n_189),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_275),
.A2(n_277),
.B1(n_295),
.B2(n_228),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_225),
.A2(n_208),
.B1(n_199),
.B2(n_188),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_173),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_216),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_283),
.Y(n_311)
);

AO22x1_ASAP7_75t_SL g282 ( 
.A1(n_232),
.A2(n_220),
.B1(n_211),
.B2(n_178),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_293),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_219),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_227),
.A2(n_176),
.B(n_190),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_39),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_2),
.B(n_3),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_289),
.A2(n_264),
.B(n_238),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_234),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_234),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_249),
.B1(n_226),
.B2(n_238),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_39),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_23),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_245),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_23),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_298),
.B(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_230),
.B(n_2),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_230),
.B(n_4),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_228),
.Y(n_322)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_239),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_303),
.B(n_309),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_281),
.B(n_283),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_308),
.B(n_241),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_243),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_247),
.C(n_235),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_326),
.C(n_284),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_243),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_314),
.B(n_317),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_322),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_268),
.B(n_282),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_316),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_272),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_318),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_319),
.A2(n_327),
.B1(n_333),
.B2(n_285),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_320),
.B(n_241),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_323),
.B(n_253),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_289),
.B1(n_276),
.B2(n_301),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_247),
.C(n_259),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_226),
.B1(n_249),
.B2(n_259),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_279),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_329),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_253),
.B1(n_250),
.B2(n_238),
.Y(n_333)
);

AOI32xp33_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_279),
.A3(n_267),
.B1(n_291),
.B2(n_268),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_339),
.B(n_315),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_340),
.A2(n_344),
.B1(n_350),
.B2(n_327),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_366),
.B1(n_320),
.B2(n_329),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_342),
.A2(n_319),
.B(n_333),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_323),
.A2(n_270),
.B1(n_282),
.B2(n_278),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_331),
.A2(n_270),
.B1(n_278),
.B2(n_273),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_356),
.C(n_302),
.Y(n_372)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_297),
.Y(n_349)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_325),
.A2(n_294),
.B1(n_292),
.B2(n_250),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_360),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_308),
.B(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_299),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_357),
.B(n_326),
.Y(n_376)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_248),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_359),
.B(n_368),
.Y(n_398)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_305),
.Y(n_362)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_313),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_365),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_324),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_364),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_231),
.B1(n_237),
.B2(n_240),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_367),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_248),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_369),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_381),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_351),
.A2(n_328),
.B(n_334),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_371),
.A2(n_345),
.B(n_353),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_377),
.C(n_378),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_374),
.A2(n_340),
.B1(n_350),
.B2(n_364),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_375),
.A2(n_387),
.B1(n_388),
.B2(n_396),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_352),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_321),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_310),
.C(n_321),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_SL g380 ( 
.A1(n_338),
.A2(n_316),
.B(n_315),
.C(n_335),
.Y(n_380)
);

AO21x1_ASAP7_75t_L g423 ( 
.A1(n_380),
.A2(n_336),
.B(n_236),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_342),
.A2(n_337),
.B(n_315),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_384),
.A2(n_371),
.B(n_391),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_311),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_237),
.C(n_264),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_341),
.A2(n_338),
.B1(n_361),
.B2(n_366),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_361),
.A2(n_315),
.B1(n_322),
.B2(n_306),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_393),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_355),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_306),
.B1(n_317),
.B2(n_311),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_337),
.A2(n_332),
.B(n_307),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_400),
.B(n_344),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_343),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_224),
.C(n_7),
.Y(n_429)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_402),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_395),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_403),
.B(n_405),
.Y(n_439)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_394),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_400),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_409),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_370),
.A2(n_357),
.B1(n_363),
.B2(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_414),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_348),
.Y(n_411)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_412),
.B(n_396),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_413),
.A2(n_415),
.B(n_419),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_370),
.A2(n_369),
.B1(n_367),
.B2(n_362),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_353),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_354),
.Y(n_416)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_416),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_387),
.A2(n_358),
.B1(n_307),
.B2(n_318),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_427),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_377),
.Y(n_435)
);

OAI31xp33_ASAP7_75t_L g421 ( 
.A1(n_380),
.A2(n_336),
.A3(n_237),
.B(n_240),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_421),
.A2(n_423),
.B(n_381),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_400),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_422),
.B(n_426),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_382),
.B(n_236),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_429),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_398),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_336),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_372),
.C(n_378),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_432),
.C(n_444),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_415),
.B(n_428),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_420),
.C(n_376),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_450),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_386),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_436),
.B(n_448),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_397),
.C(n_388),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_425),
.C(n_413),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_432),
.C(n_435),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_384),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_375),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_423),
.Y(n_470)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_439),
.Y(n_453)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_426),
.Y(n_454)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_424),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_456),
.Y(n_481)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_438),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_462),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_470),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_407),
.B1(n_415),
.B2(n_422),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_459),
.A2(n_461),
.B1(n_463),
.B2(n_468),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_434),
.A2(n_403),
.B1(n_402),
.B2(n_409),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_411),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_440),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_421),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_464),
.A2(n_467),
.B1(n_431),
.B2(n_452),
.Y(n_473)
);

FAx1_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_428),
.CI(n_380),
.CON(n_465),
.SN(n_465)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_423),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_418),
.B1(n_406),
.B2(n_428),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_471),
.A2(n_414),
.B(n_416),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_430),
.C(n_448),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_475),
.C(n_476),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_480),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_437),
.C(n_444),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_437),
.C(n_436),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_442),
.B1(n_404),
.B2(n_433),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_478),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_483),
.B(n_484),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_450),
.C(n_373),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_385),
.C(n_427),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_487),
.C(n_488),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_385),
.C(n_379),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_467),
.C(n_465),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_486),
.Y(n_490)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_481),
.A2(n_458),
.B(n_465),
.Y(n_491)
);

AO21x1_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_492),
.B(n_6),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_472),
.A2(n_488),
.B(n_479),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_482),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_494),
.Y(n_504)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_464),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_496),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_390),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_389),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_501),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_399),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_399),
.B1(n_380),
.B2(n_224),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_502),
.A2(n_487),
.B1(n_8),
.B2(n_10),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_503),
.A2(n_489),
.B1(n_11),
.B2(n_12),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_506),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_497),
.B(n_6),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_509),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_6),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_489),
.C(n_496),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_511),
.A2(n_11),
.B(n_12),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_495),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_512),
.A2(n_504),
.B(n_511),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_8),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g517 ( 
.A1(n_513),
.A2(n_499),
.B(n_500),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_507),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_519),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_520),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_11),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_521),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_517),
.B(n_516),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_527),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_523),
.B(n_510),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_524),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_522),
.B1(n_515),
.B2(n_514),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_528),
.B(n_13),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_12),
.C(n_13),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_13),
.C(n_15),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_15),
.B(n_16),
.Y(n_534)
);


endmodule