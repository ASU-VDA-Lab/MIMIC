module fake_jpeg_24964_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_28),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_21),
.B1(n_20),
.B2(n_34),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_69),
.B1(n_42),
.B2(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_21),
.B1(n_20),
.B2(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_34),
.B1(n_22),
.B2(n_28),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_22),
.B(n_23),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_47),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_47),
.C(n_40),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_92),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_47),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_94),
.B(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_83),
.Y(n_108)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_93),
.B1(n_92),
.B2(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_91),
.Y(n_119)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_87),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_39),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_97),
.B1(n_55),
.B2(n_76),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_40),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_29),
.B1(n_23),
.B2(n_41),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_41),
.B1(n_37),
.B2(n_45),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_96),
.B(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_39),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_47),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_40),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_126),
.B(n_131),
.Y(n_142)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_116),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_117),
.B1(n_103),
.B2(n_48),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_132),
.B1(n_84),
.B2(n_76),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_75),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_29),
.B(n_89),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_129),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_134),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_40),
.B(n_52),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_77),
.A2(n_48),
.B1(n_45),
.B2(n_37),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_40),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_68),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_141),
.B1(n_157),
.B2(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_152),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_80),
.B1(n_100),
.B2(n_82),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_102),
.B1(n_88),
.B2(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

AO22x1_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_106),
.B1(n_94),
.B2(n_103),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_124),
.B1(n_120),
.B2(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_88),
.B1(n_90),
.B2(n_106),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_161),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_73),
.B1(n_99),
.B2(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_17),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_83),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_89),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_25),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_39),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_167),
.Y(n_195)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_26),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_25),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_25),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_22),
.B(n_19),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_166),
.A2(n_136),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_17),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_122),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_175),
.C(n_194),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_169),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_150),
.B(n_166),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_173),
.B(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_172),
.B(n_178),
.Y(n_227)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_150),
.B(n_167),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_115),
.B1(n_112),
.B2(n_107),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_181),
.B1(n_139),
.B2(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_196),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_183),
.A2(n_189),
.B1(n_7),
.B2(n_14),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_111),
.B1(n_124),
.B2(n_120),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_111),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_200),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_146),
.A2(n_114),
.B(n_110),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_129),
.B1(n_30),
.B2(n_36),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_156),
.A2(n_31),
.B(n_33),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_201),
.B1(n_138),
.B2(n_24),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_25),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_31),
.B1(n_24),
.B2(n_17),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_24),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_219),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_159),
.B(n_137),
.C(n_157),
.D(n_24),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_207),
.B(n_15),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_181),
.B(n_187),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_232),
.B(n_173),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_230),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_138),
.B1(n_149),
.B2(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_149),
.B1(n_25),
.B2(n_2),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_231),
.B1(n_180),
.B2(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_193),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_228),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_16),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_182),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_233),
.A2(n_237),
.B1(n_243),
.B2(n_258),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_171),
.B1(n_197),
.B2(n_184),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_168),
.C(n_195),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_252),
.C(n_253),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_175),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_247),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_183),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_194),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_250),
.B(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_188),
.C(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_189),
.C(n_1),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

HAxp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_229),
.CON(n_259),
.SN(n_259)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_259),
.A2(n_265),
.B(n_274),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_205),
.B1(n_219),
.B2(n_215),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_267),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_271),
.Y(n_285)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_224),
.B(n_208),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_208),
.B1(n_204),
.B2(n_221),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_222),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_210),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_244),
.B(n_231),
.CI(n_207),
.CON(n_273),
.SN(n_273)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_SL g274 ( 
.A(n_243),
.B(n_218),
.C(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_247),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_220),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_287),
.C(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_217),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_286),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_259),
.A2(n_233),
.B1(n_239),
.B2(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_263),
.B1(n_206),
.B2(n_276),
.Y(n_303)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_295),
.C(n_206),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_273),
.B(n_255),
.Y(n_294)
);

AO22x1_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_298),
.B1(n_263),
.B2(n_252),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_261),
.C(n_270),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx11_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_SL g298 ( 
.A1(n_261),
.A2(n_217),
.B(n_235),
.C(n_253),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_299),
.B(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_236),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_301),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_235),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_298),
.B1(n_3),
.B2(n_4),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_304),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_295),
.C(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_6),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_311),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_287),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_309),
.A2(n_298),
.B1(n_12),
.B2(n_13),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_0),
.C(n_1),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_281),
.A2(n_14),
.B(n_10),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_292),
.A2(n_5),
.B(n_11),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_294),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_11),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_324),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_294),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_305),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_293),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_320),
.C(n_304),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_322),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_285),
.B1(n_288),
.B2(n_291),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_284),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_SL g330 ( 
.A(n_321),
.B(n_307),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_332),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_314),
.A2(n_311),
.B(n_310),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_330),
.B(n_331),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_308),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_302),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_323),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_325),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_339),
.B(n_327),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

AOI21x1_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_327),
.B(n_315),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_342),
.A2(n_343),
.B(n_335),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_336),
.B(n_341),
.C(n_318),
.Y(n_345)
);

AOI321xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_12),
.A3(n_13),
.B1(n_4),
.B2(n_0),
.C(n_3),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_4),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_4),
.Y(n_348)
);


endmodule