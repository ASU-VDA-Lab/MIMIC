module fake_jpeg_25596_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_31),
.B1(n_23),
.B2(n_24),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_54),
.B1(n_63),
.B2(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_23),
.B1(n_31),
.B2(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_25),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_23),
.B1(n_33),
.B2(n_24),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_64),
.B1(n_25),
.B2(n_22),
.Y(n_80)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_21),
.B1(n_27),
.B2(n_17),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_25),
.B1(n_22),
.B2(n_17),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_55),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_83),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_11),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_86),
.Y(n_92)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_87),
.B(n_89),
.C(n_58),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_64),
.B1(n_61),
.B2(n_53),
.Y(n_110)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_88),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_9),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_44),
.B(n_28),
.CI(n_32),
.CON(n_87),
.SN(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_32),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_102),
.Y(n_137)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_51),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_79),
.C(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_109),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_89),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_48),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_81),
.B1(n_67),
.B2(n_65),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_77),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_59),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_53),
.B1(n_43),
.B2(n_62),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_81),
.B1(n_67),
.B2(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_49),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_70),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_78),
.B1(n_84),
.B2(n_79),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_108),
.B1(n_98),
.B2(n_109),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_139),
.B(n_98),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_105),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_120),
.B1(n_128),
.B2(n_134),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_87),
.C(n_66),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_99),
.C(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_68),
.B1(n_74),
.B2(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_131),
.Y(n_146)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_16),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_16),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_0),
.B(n_15),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_95),
.B(n_0),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_104),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_143),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_107),
.B1(n_108),
.B2(n_99),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_156),
.B(n_141),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_111),
.B(n_108),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_122),
.B(n_125),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_167),
.Y(n_171)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_0),
.B(n_101),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_91),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_118),
.C(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_104),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_91),
.B1(n_104),
.B2(n_4),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_119),
.B1(n_132),
.B2(n_131),
.Y(n_177)
);

NAND2xp33_ASAP7_75t_R g166 ( 
.A(n_134),
.B(n_139),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_124),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_175),
.A2(n_176),
.B(n_187),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_164),
.B1(n_163),
.B2(n_161),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_189),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_135),
.B1(n_124),
.B2(n_121),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_184),
.B1(n_154),
.B2(n_165),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_147),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_127),
.B1(n_125),
.B2(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_159),
.C(n_144),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_198),
.C(n_210),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_192),
.B1(n_185),
.B2(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_182),
.C(n_183),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_184),
.B1(n_176),
.B2(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_150),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_174),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_149),
.C(n_146),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_146),
.C(n_145),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_168),
.C(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_171),
.B1(n_169),
.B2(n_177),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_225),
.B1(n_211),
.B2(n_210),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_224),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_223),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_174),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_198),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_172),
.C(n_151),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_151),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_200),
.B1(n_167),
.B2(n_194),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_212),
.B(n_204),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_231),
.A2(n_240),
.B(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_203),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_234),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_217),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_200),
.B(n_199),
.C(n_170),
.D(n_179),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_239),
.C(n_8),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_199),
.B(n_156),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_155),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_220),
.C(n_221),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_242),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_249),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_217),
.C(n_224),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_15),
.C(n_9),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_216),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_250),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_226),
.B(n_3),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_251),
.B(n_6),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_237),
.C(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_257),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_251),
.B1(n_255),
.B2(n_257),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_8),
.B(n_9),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.C(n_261),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_252),
.A2(n_8),
.B(n_10),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_10),
.C(n_13),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_266),
.B(n_13),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_269),
.B(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_10),
.Y(n_272)
);


endmodule