module fake_jpeg_24696_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_16),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_42),
.B1(n_23),
.B2(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_40),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_27),
.B(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_56),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_23),
.Y(n_48)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_52),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_33),
.B(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_17),
.B1(n_21),
.B2(n_27),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_20),
.B1(n_26),
.B2(n_30),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_17),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_37),
.C(n_34),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_62),
.A2(n_24),
.B(n_31),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_65),
.Y(n_91)
);

AOI22x1_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_34),
.B1(n_35),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_78),
.B1(n_47),
.B2(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_75),
.C(n_85),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_37),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_41),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_82),
.B(n_65),
.C(n_80),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_53),
.B1(n_39),
.B2(n_45),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_29),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_35),
.B1(n_41),
.B2(n_38),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_83),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_38),
.CI(n_41),
.CON(n_82),
.SN(n_82)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_55),
.CI(n_53),
.CON(n_94),
.SN(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_2),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_92),
.B1(n_101),
.B2(n_81),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_24),
.C(n_31),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_98),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_39),
.B(n_40),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_94),
.B(n_102),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_55),
.B1(n_44),
.B2(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_71),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_53),
.B1(n_60),
.B2(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_53),
.B1(n_79),
.B2(n_60),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_72),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_102),
.B(n_91),
.Y(n_135)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_38),
.Y(n_134)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_67),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_87),
.C(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_101),
.B1(n_102),
.B2(n_94),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_82),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_68),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_79),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_111),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_134),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_116),
.B1(n_129),
.B2(n_132),
.C(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_147),
.C(n_151),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_112),
.B1(n_133),
.B2(n_115),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_88),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_154),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_93),
.C(n_110),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_25),
.C(n_18),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_94),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_29),
.B(n_25),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_116),
.C(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_63),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_85),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_114),
.B(n_73),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_120),
.C(n_124),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_151),
.C(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_109),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_117),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_165),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_175),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_114),
.B(n_69),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_113),
.B1(n_117),
.B2(n_103),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_147),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_113),
.B1(n_103),
.B2(n_109),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_38),
.Y(n_171)
);

OAI22x1_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_70),
.B1(n_21),
.B2(n_27),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_109),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_99),
.B1(n_52),
.B2(n_44),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_146),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_191),
.B(n_192),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_136),
.C(n_144),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_188),
.C(n_168),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_149),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_166),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_144),
.C(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_145),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_143),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_199),
.C(n_201),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_175),
.C(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_197),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_174),
.CI(n_166),
.CON(n_196),
.SN(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_180),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_172),
.B1(n_163),
.B2(n_156),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_189),
.B1(n_184),
.B2(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_171),
.C(n_170),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_184),
.A2(n_18),
.B(n_3),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_2),
.B(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_182),
.B1(n_187),
.B2(n_22),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_206),
.B1(n_201),
.B2(n_8),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_182),
.B1(n_3),
.B2(n_4),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_19),
.C(n_5),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_210),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_7),
.B(n_8),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_5),
.C(n_6),
.Y(n_210)
);

OAI221xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_198),
.B1(n_202),
.B2(n_203),
.C(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_200),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_218),
.B(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_217),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_210),
.B(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_219),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_208),
.B(n_207),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_208),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_228),
.A3(n_224),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_230),
.B1(n_226),
.B2(n_11),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_225),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_14),
.Y(n_232)
);


endmodule