module real_jpeg_218_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_25),
.C(n_38),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_7),
.B(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_23),
.C(n_30),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_7),
.B(n_54),
.C(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_58),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_7),
.B(n_69),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_8),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_94),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_93),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_80),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_61),
.C(n_76),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_46),
.B2(n_60),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_17),
.A2(n_18),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_35),
.B2(n_45),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_45),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_19),
.A2(n_20),
.B1(n_67),
.B2(n_68),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_19),
.A2(n_20),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_19),
.A2(n_68),
.B(n_79),
.C(n_152),
.Y(n_155)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_67),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_20),
.B(n_51),
.C(n_104),
.Y(n_103)
);

AO21x2_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_22)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

OA22x2_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_25),
.B(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_29),
.Y(n_137)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_30),
.A2(n_32),
.B1(n_70),
.B2(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_30),
.B(n_131),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_35),
.A2(n_45),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AO21x2_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_44),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

AOI211xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_68),
.B(n_78),
.C(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_50),
.A2(n_51),
.B1(n_104),
.B2(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_50),
.A2(n_51),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_50),
.A2(n_51),
.B1(n_118),
.B2(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_51),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_51),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_67),
.C(n_136),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_58),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_54),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_54),
.B(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_76),
.B1(n_77),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_75),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_68),
.B1(n_89),
.B2(n_92),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_113),
.C(n_117),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_68),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_68),
.B1(n_129),
.B2(n_130),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_67),
.A2(n_68),
.B1(n_117),
.B2(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_129),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B(n_74),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_73),
.Y(n_72)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_109),
.B(n_161),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_97),
.B(n_106),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_103),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_99),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_101),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_124),
.B(n_160),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_121),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_154),
.B(n_159),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_148),
.B(n_153),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_138),
.B(n_147),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_132),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);


endmodule