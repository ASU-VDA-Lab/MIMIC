module fake_jpeg_12348_n_615 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_615);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_615;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_0),
.B(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_7),
.B(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx8_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_61),
.Y(n_205)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_64),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_65),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_68),
.B(n_110),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_88),
.Y(n_133)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_89),
.B(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_93),
.Y(n_198)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_94),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_25),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_114),
.Y(n_182)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_97),
.Y(n_208)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_34),
.B(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_126),
.Y(n_150)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

CKINVDCx6p67_ASAP7_75t_R g179 ( 
.A(n_109),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_113),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_115),
.B(n_122),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_24),
.Y(n_119)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_34),
.B(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_128),
.Y(n_197)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_29),
.Y(n_169)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_27),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_28),
.B1(n_44),
.B2(n_50),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_131),
.A2(n_191),
.B1(n_9),
.B2(n_10),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_67),
.A2(n_44),
.B1(n_39),
.B2(n_27),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_138),
.A2(n_146),
.B1(n_154),
.B2(n_155),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_69),
.A2(n_39),
.B1(n_37),
.B2(n_49),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_139),
.A2(n_185),
.B1(n_196),
.B2(n_203),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_74),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_95),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_153),
.B(n_159),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_29),
.B1(n_51),
.B2(n_38),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_84),
.A2(n_29),
.B1(n_51),
.B2(n_40),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_90),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_58),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_204),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_169),
.B(n_201),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_98),
.A2(n_40),
.B1(n_43),
.B2(n_58),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_172),
.A2(n_186),
.B1(n_194),
.B2(n_9),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_68),
.B(n_49),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_210),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_66),
.A2(n_26),
.B1(n_50),
.B2(n_23),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_111),
.A2(n_43),
.B1(n_23),
.B2(n_26),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_72),
.A2(n_78),
.B1(n_126),
.B2(n_121),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_118),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_73),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_64),
.B(n_2),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_200),
.B(n_202),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_127),
.B(n_3),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_79),
.B(n_3),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_80),
.A2(n_52),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_83),
.B(n_52),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_92),
.B(n_5),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_5),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_97),
.B(n_5),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_99),
.A2(n_52),
.B1(n_7),
.B2(n_8),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_215),
.B(n_272),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_217),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_120),
.C(n_117),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_218),
.B(n_287),
.C(n_198),
.Y(n_297)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_221),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_116),
.B1(n_113),
.B2(n_100),
.Y(n_222)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_222),
.A2(n_154),
.B1(n_164),
.B2(n_161),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_223),
.B(n_234),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_150),
.B(n_8),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_224),
.B(n_271),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_226),
.Y(n_336)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_229),
.Y(n_323)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_231),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_136),
.Y(n_232)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_233),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_131),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_236),
.A2(n_243),
.B1(n_254),
.B2(n_199),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_134),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_240),
.A2(n_214),
.B1(n_222),
.B2(n_287),
.Y(n_337)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_242),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_9),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_244),
.B(n_269),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_245),
.A2(n_257),
.B1(n_278),
.B2(n_241),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_136),
.Y(n_246)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_133),
.B(n_12),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_248),
.B(n_252),
.Y(n_309)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_160),
.B(n_15),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_182),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_253),
.B(n_261),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_191),
.A2(n_16),
.B1(n_185),
.B2(n_211),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_143),
.Y(n_255)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_255),
.Y(n_313)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_186),
.A2(n_16),
.B1(n_138),
.B2(n_172),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_201),
.A2(n_209),
.B(n_176),
.C(n_155),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_258),
.B(n_266),
.Y(n_342)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_137),
.Y(n_259)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_173),
.Y(n_260)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_165),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_136),
.Y(n_263)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_143),
.Y(n_264)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_268),
.Y(n_341)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_142),
.Y(n_266)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_144),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_157),
.B(n_149),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_213),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_147),
.B(n_181),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_130),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_273),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_274),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_132),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_275),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_157),
.B(n_145),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_277),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_205),
.A2(n_162),
.B1(n_140),
.B2(n_189),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_175),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_279),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_137),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_284),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_179),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_141),
.B(n_148),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_286),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_179),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_192),
.B(n_140),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_161),
.B(n_208),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_222),
.Y(n_343)
);

AOI32xp33_ASAP7_75t_L g290 ( 
.A1(n_238),
.A2(n_198),
.A3(n_146),
.B1(n_205),
.B2(n_194),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_290),
.A2(n_301),
.B(n_300),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_296),
.A2(n_308),
.B1(n_326),
.B2(n_287),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_297),
.B(n_276),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_237),
.A2(n_177),
.B(n_175),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_301),
.A2(n_281),
.B(n_226),
.Y(n_367)
);

AO21x2_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_208),
.B(n_184),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_305),
.A2(n_310),
.B1(n_337),
.B2(n_260),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_216),
.A2(n_164),
.B1(n_177),
.B2(n_174),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g310 ( 
.A1(n_216),
.A2(n_184),
.B1(n_174),
.B2(n_168),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_258),
.B(n_271),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_321),
.A2(n_276),
.B(n_240),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_220),
.A2(n_214),
.B1(n_168),
.B2(n_199),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_255),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_224),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_346),
.B(n_350),
.Y(n_416)
);

AO21x1_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_368),
.B(n_381),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_348),
.B(n_358),
.C(n_361),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_349),
.A2(n_356),
.B1(n_372),
.B2(n_373),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_276),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_352),
.A2(n_296),
.B1(n_344),
.B2(n_334),
.Y(n_390)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

NAND2x1_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_222),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_355),
.A2(n_316),
.B(n_292),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_218),
.B1(n_282),
.B2(n_225),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_268),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_357),
.B(n_363),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_267),
.Y(n_358)
);

INVx5_ASAP7_75t_SL g359 ( 
.A(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_359),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_334),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_360),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_266),
.C(n_272),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_306),
.B(n_247),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_291),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_365),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_318),
.B(n_259),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_366),
.A2(n_331),
.B1(n_311),
.B2(n_304),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_367),
.A2(n_379),
.B(n_383),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_321),
.B(n_219),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_368),
.B(n_374),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_342),
.B(n_273),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_369),
.B(n_382),
.Y(n_411)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_371),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_315),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_305),
.A2(n_230),
.B1(n_264),
.B2(n_274),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_300),
.A2(n_221),
.B1(n_235),
.B2(n_280),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_295),
.B(n_279),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_249),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_375),
.B(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_239),
.B1(n_232),
.B2(n_246),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_377),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_308),
.A2(n_217),
.B1(n_283),
.B2(n_263),
.Y(n_378)
);

INVx3_ASAP7_75t_SL g403 ( 
.A(n_378),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_322),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_297),
.B(n_273),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_381),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_342),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_305),
.B(n_315),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_309),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_299),
.B(n_330),
.C(n_340),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_389),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_329),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_386),
.Y(n_398)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_387),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_305),
.A2(n_296),
.B1(n_310),
.B2(n_298),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_331),
.B1(n_344),
.B2(n_320),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_305),
.B(n_303),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_390),
.A2(n_425),
.B1(n_426),
.B2(n_373),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_397),
.A2(n_400),
.B1(n_414),
.B2(n_366),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_388),
.A2(n_294),
.B1(n_311),
.B2(n_325),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_361),
.A2(n_367),
.B(n_371),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_406),
.A2(n_413),
.B(n_417),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_407),
.A2(n_412),
.B(n_369),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_359),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_419),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_354),
.A2(n_289),
.B(n_292),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_349),
.A2(n_294),
.B1(n_323),
.B2(n_302),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_289),
.B(n_317),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_307),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_374),
.C(n_375),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_359),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_362),
.A2(n_335),
.B1(n_307),
.B2(n_332),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_347),
.A2(n_335),
.B1(n_319),
.B2(n_316),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_402),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_433),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_389),
.B(n_380),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_430),
.A2(n_457),
.B(n_399),
.Y(n_486)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_358),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_444),
.C(n_448),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_357),
.Y(n_435)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g480 ( 
.A1(n_436),
.A2(n_441),
.B1(n_403),
.B2(n_423),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_420),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_411),
.Y(n_474)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_439),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_415),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_440),
.B(n_449),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_394),
.B(n_383),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_442),
.B(n_456),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_346),
.Y(n_443)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_420),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_392),
.A2(n_379),
.B1(n_355),
.B2(n_350),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_445),
.A2(n_446),
.B1(n_452),
.B2(n_453),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_392),
.A2(n_355),
.B1(n_356),
.B2(n_372),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_447),
.A2(n_422),
.B1(n_412),
.B2(n_417),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_363),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_415),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_391),
.Y(n_462)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_458),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_400),
.A2(n_365),
.B1(n_384),
.B2(n_353),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_404),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_385),
.B1(n_376),
.B2(n_370),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_454),
.A2(n_460),
.B1(n_390),
.B2(n_423),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_394),
.B(n_319),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_401),
.A2(n_317),
.B(n_304),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_414),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_416),
.B(n_364),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_459),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_404),
.A2(n_351),
.B1(n_329),
.B2(n_324),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_462),
.B(n_443),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_391),
.C(n_411),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_478),
.C(n_479),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_471),
.A2(n_480),
.B1(n_447),
.B2(n_455),
.Y(n_505)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_474),
.B(n_437),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_427),
.A2(n_416),
.B1(n_407),
.B2(n_403),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_398),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_432),
.B(n_406),
.C(n_405),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_405),
.C(n_426),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_423),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_429),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_446),
.A2(n_403),
.B1(n_425),
.B2(n_422),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_482),
.A2(n_486),
.B1(n_487),
.B2(n_457),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_434),
.A2(n_419),
.B(n_409),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_483),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_454),
.Y(n_484)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_458),
.A2(n_445),
.B1(n_453),
.B2(n_441),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_456),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_491),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_399),
.Y(n_490)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_490),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_442),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_492),
.B(n_496),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_476),
.Y(n_495)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_495),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_450),
.C(n_434),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_502),
.C(n_504),
.Y(n_541)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_490),
.Y(n_501)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_463),
.B(n_438),
.C(n_431),
.Y(n_502)
);

MAJx2_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_511),
.C(n_513),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_430),
.C(n_428),
.Y(n_504)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_452),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_506),
.B(n_518),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_475),
.A2(n_433),
.B1(n_449),
.B2(n_440),
.Y(n_507)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_507),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_462),
.B(n_479),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_510),
.Y(n_522)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_435),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_460),
.C(n_451),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_512),
.A2(n_486),
.B(n_489),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_474),
.B(n_459),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_439),
.Y(n_514)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_514),
.Y(n_536)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_465),
.A2(n_398),
.B1(n_436),
.B2(n_393),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_471),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_489),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_469),
.B(n_393),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_477),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_497),
.A2(n_465),
.B1(n_487),
.B2(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_521),
.Y(n_551)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_494),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_533),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_483),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_531),
.B(n_535),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_514),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_534),
.A2(n_542),
.B1(n_467),
.B2(n_500),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_469),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_516),
.A2(n_473),
.B(n_482),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_537),
.B(n_533),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_SL g539 ( 
.A(n_504),
.B(n_498),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_540),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_473),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_510),
.C(n_493),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_545),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_493),
.C(n_511),
.Y(n_545)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_546),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_541),
.B(n_516),
.C(n_496),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_547),
.B(n_554),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_499),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_548),
.B(n_552),
.Y(n_571)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_524),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_549),
.B(n_467),
.Y(n_568)
);

CKINVDCx14_ASAP7_75t_R g552 ( 
.A(n_523),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_497),
.C(n_513),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_540),
.C(n_528),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_555),
.B(n_557),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_492),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_560),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_526),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_532),
.B(n_509),
.C(n_512),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_558),
.B(n_527),
.C(n_535),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_525),
.B(n_464),
.C(n_500),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_559),
.B(n_521),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_563),
.B(n_573),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_560),
.A2(n_537),
.B(n_527),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_564),
.A2(n_395),
.B(n_424),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_543),
.B(n_529),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_556),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_567),
.Y(n_578)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_551),
.A2(n_525),
.B1(n_536),
.B2(n_542),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_570),
.B(n_576),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_520),
.C(n_530),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_545),
.B(n_519),
.C(n_538),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_544),
.C(n_550),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_558),
.B(n_395),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_575),
.B(n_468),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_548),
.A2(n_461),
.B(n_468),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_561),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_572),
.A2(n_461),
.B1(n_549),
.B2(n_550),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_579),
.B(n_583),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_574),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_582),
.B(n_561),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_564),
.A2(n_553),
.B1(n_436),
.B2(n_424),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_553),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_588),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_586),
.B(n_576),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_571),
.B(n_328),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_587),
.A2(n_562),
.B(n_569),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_590),
.A2(n_578),
.B(n_586),
.Y(n_603)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_591),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_577),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_573),
.C(n_563),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_595),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_596),
.B(n_597),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_571),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_570),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_581),
.Y(n_602)
);

AOI31xp33_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_589),
.A3(n_579),
.B(n_591),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_603),
.B(n_604),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_594),
.A2(n_581),
.B(n_588),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_605),
.B(n_593),
.C(n_592),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_606),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_607),
.A2(n_608),
.B(n_600),
.Y(n_610)
);

OAI311xp33_ASAP7_75t_L g608 ( 
.A1(n_599),
.A2(n_583),
.A3(n_566),
.B1(n_320),
.C1(n_314),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_610),
.B(n_601),
.C(n_606),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_612),
.A2(n_611),
.B1(n_609),
.B2(n_336),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_613),
.B(n_336),
.Y(n_614)
);

HAxp5_ASAP7_75t_SL g615 ( 
.A(n_614),
.B(n_328),
.CON(n_615),
.SN(n_615)
);


endmodule