module fake_jpeg_10128_n_227 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_46),
.Y(n_74)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_54),
.B1(n_58),
.B2(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_51),
.B1(n_17),
.B2(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_15),
.B1(n_27),
.B2(n_26),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_35),
.B1(n_39),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_17),
.B1(n_28),
.B2(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_55),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_31),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_23),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_67),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_64),
.B1(n_73),
.B2(n_75),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_38),
.B(n_34),
.C(n_39),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_74),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_38),
.B1(n_34),
.B2(n_35),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_40),
.B1(n_36),
.B2(n_23),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_23),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_47),
.C(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_82),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_40),
.B1(n_36),
.B2(n_23),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_102),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_36),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_55),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_40),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_71),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_78),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_107),
.B(n_123),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_116),
.B1(n_119),
.B2(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_82),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_66),
.B1(n_65),
.B2(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_81),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_83),
.B(n_90),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_56),
.B1(n_42),
.B2(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_64),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_88),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_45),
.B1(n_60),
.B2(n_43),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_45),
.B1(n_81),
.B2(n_77),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_93),
.B1(n_84),
.B2(n_100),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_138),
.B1(n_147),
.B2(n_117),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_134),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_90),
.Y(n_135)
);

NOR2x1_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_143),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_145),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_97),
.B1(n_85),
.B2(n_91),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_123),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_85),
.B1(n_45),
.B2(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_157),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_113),
.C(n_115),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_133),
.C(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_158),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_109),
.B1(n_121),
.B2(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_107),
.B1(n_122),
.B2(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_162),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_111),
.B1(n_52),
.B2(n_77),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_145),
.B(n_130),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_133),
.C(n_143),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g170 ( 
.A(n_164),
.B(n_134),
.C(n_135),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_174),
.B1(n_165),
.B2(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_146),
.C(n_135),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_152),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_154),
.B1(n_150),
.B2(n_157),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_53),
.B1(n_18),
.B2(n_5),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_184),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_154),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_187),
.B1(n_184),
.B2(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_81),
.B1(n_86),
.B2(n_92),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_176),
.B1(n_86),
.B2(n_53),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_201),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_168),
.C(n_167),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_196),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_200),
.B1(n_3),
.B2(n_5),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_180),
.B(n_2),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_188),
.B1(n_185),
.B2(n_186),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_209),
.B1(n_194),
.B2(n_9),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_197),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_207),
.B(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_6),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_189),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_213),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_8),
.C(n_10),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_206),
.B(n_10),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_211),
.A3(n_215),
.B1(n_206),
.B2(n_13),
.C1(n_11),
.C2(n_12),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_11),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_218),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_224),
.C(n_12),
.Y(n_227)
);


endmodule