module fake_ariane_1771_n_770 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_770);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_770;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_515;
wire n_445;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_3),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_8),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_56),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_13),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_16),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_10),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_103),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_43),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_16),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_17),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_57),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_93),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_2),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_104),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_55),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_47),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_25),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_22),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_8),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_24),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_86),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_50),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_6),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_28),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_36),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_21),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_0),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_0),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_152),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_3),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_161),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_4),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_5),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_5),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_7),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_145),
.B(n_7),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_9),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_153),
.B(n_9),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_148),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_148),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_146),
.B(n_165),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_10),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_147),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_149),
.B(n_11),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_196),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_159),
.B1(n_191),
.B2(n_186),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_159),
.B1(n_191),
.B2(n_202),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_196),
.B1(n_193),
.B2(n_177),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_176),
.B1(n_180),
.B2(n_178),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_192),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_185),
.B1(n_183),
.B2(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_162),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_163),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_179),
.B1(n_173),
.B2(n_170),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_205),
.A2(n_222),
.B1(n_212),
.B2(n_225),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_164),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_169),
.B1(n_168),
.B2(n_167),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_202),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_217),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_19),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_202),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_23),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_23),
.Y(n_264)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_265)
);

AOI22x1_ASAP7_75t_SL g266 ( 
.A1(n_229),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_31),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_209),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_217),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_207),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_219),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

OR2x6_ASAP7_75t_L g274 ( 
.A(n_199),
.B(n_48),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_216),
.B(n_49),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_216),
.B(n_142),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_218),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_224),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_199),
.B(n_61),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_236),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

BUFx8_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_218),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_247),
.A2(n_237),
.B(n_226),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_226),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_239),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_235),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx4_ASAP7_75t_SL g309 ( 
.A(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_280),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_235),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

OR2x6_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_225),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_237),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_255),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_246),
.B(n_198),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_218),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_258),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_243),
.B(n_218),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_232),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_203),
.B(n_221),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_244),
.B(n_233),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_268),
.A2(n_211),
.B(n_220),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

NAND2x1p5_ASAP7_75t_L g343 ( 
.A(n_266),
.B(n_208),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_238),
.B(n_232),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_248),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_248),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_248),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_248),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_232),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_213),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_346),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_299),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_289),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_346),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_286),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_291),
.A2(n_232),
.B1(n_214),
.B2(n_206),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_232),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_305),
.B(n_200),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_296),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_298),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_200),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_296),
.B(n_206),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_296),
.B(n_206),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_206),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_329),
.B(n_230),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_214),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_324),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_294),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_290),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_287),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_301),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_301),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_214),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_214),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_67),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_318),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_323),
.B(n_214),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_319),
.B(n_200),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_331),
.B(n_68),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_69),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_318),
.B(n_70),
.Y(n_393)
);

OR2x2_ASAP7_75t_SL g394 ( 
.A(n_320),
.B(n_71),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_330),
.B(n_72),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_200),
.Y(n_396)
);

BUFx8_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_323),
.B(n_200),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_306),
.B(n_200),
.Y(n_400)
);

BUFx12f_ASAP7_75t_L g401 ( 
.A(n_289),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_317),
.B(n_73),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_307),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_308),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_317),
.B(n_74),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_334),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_75),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_141),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_310),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_311),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_292),
.B(n_76),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_330),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_292),
.B(n_138),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_337),
.B(n_77),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_322),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_401),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_380),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_378),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_321),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_315),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_313),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_303),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_328),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_327),
.Y(n_429)
);

OR2x6_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_343),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_338),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_339),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_375),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_289),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_78),
.Y(n_441)
);

INVx8_ASAP7_75t_L g442 ( 
.A(n_383),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_369),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_364),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_365),
.B(n_343),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_406),
.B(n_79),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_80),
.Y(n_452)
);

NAND2x1p5_ASAP7_75t_L g453 ( 
.A(n_351),
.B(n_81),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_365),
.B(n_82),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_403),
.B(n_377),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_403),
.B(n_83),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_354),
.Y(n_458)
);

NAND2x1p5_ASAP7_75t_L g459 ( 
.A(n_354),
.B(n_407),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_364),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_365),
.B(n_84),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_85),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_383),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_377),
.B(n_87),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_350),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_88),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_372),
.B(n_90),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_393),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_377),
.B(n_91),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_399),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_423),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_420),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_447),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_419),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_447),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_417),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_424),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_434),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_442),
.Y(n_487)
);

CKINVDCx6p67_ASAP7_75t_R g488 ( 
.A(n_430),
.Y(n_488)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

NAND2x1p5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_393),
.Y(n_491)
);

NOR2x1_ASAP7_75t_SL g492 ( 
.A(n_448),
.B(n_414),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_418),
.Y(n_493)
);

BUFx2_ASAP7_75t_R g494 ( 
.A(n_438),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_442),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_456),
.A2(n_390),
.B1(n_405),
.B2(n_402),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_442),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_430),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_448),
.B(n_393),
.Y(n_502)
);

BUFx8_ASAP7_75t_L g503 ( 
.A(n_440),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_451),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_418),
.Y(n_506)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_430),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_417),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_466),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_393),
.Y(n_515)
);

BUFx12f_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_425),
.B(n_402),
.Y(n_518)
);

BUFx4_ASAP7_75t_SL g519 ( 
.A(n_449),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_478),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_484),
.Y(n_521)
);

OAI22x1_ASAP7_75t_L g522 ( 
.A1(n_483),
.A2(n_464),
.B1(n_392),
.B2(n_471),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_499),
.A2(n_409),
.B(n_357),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_456),
.B1(n_440),
.B2(n_464),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_485),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_518),
.A2(n_440),
.B1(n_429),
.B2(n_392),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_486),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_494),
.Y(n_528)
);

CKINVDCx11_ASAP7_75t_R g529 ( 
.A(n_480),
.Y(n_529)
);

CKINVDCx11_ASAP7_75t_R g530 ( 
.A(n_480),
.Y(n_530)
);

BUFx4f_ASAP7_75t_SL g531 ( 
.A(n_481),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_514),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_504),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_493),
.Y(n_534)
);

BUFx8_ASAP7_75t_L g535 ( 
.A(n_516),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_493),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_503),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_510),
.Y(n_538)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_503),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_496),
.A2(n_440),
.B1(n_429),
.B2(n_379),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_516),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_477),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_475),
.A2(n_429),
.B1(n_405),
.B2(n_422),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_500),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_509),
.A2(n_429),
.B1(n_470),
.B2(n_443),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_475),
.A2(n_429),
.B1(n_422),
.B2(n_435),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_517),
.A2(n_470),
.B1(n_425),
.B2(n_356),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_509),
.A2(n_470),
.B1(n_356),
.B2(n_363),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_506),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_488),
.A2(n_363),
.B1(n_446),
.B2(n_461),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_504),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_515),
.A2(n_459),
.B1(n_472),
.B2(n_467),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_506),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_488),
.A2(n_363),
.B1(n_446),
.B2(n_461),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_510),
.A2(n_386),
.B1(n_384),
.B2(n_459),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_489),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_511),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_513),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_513),
.B(n_426),
.Y(n_560)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_503),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_520),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_537),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_543),
.A2(n_394),
.B1(n_515),
.B2(n_472),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_526),
.A2(n_515),
.B(n_394),
.Y(n_565)
);

AOI222xp33_ASAP7_75t_L g566 ( 
.A1(n_522),
.A2(n_397),
.B1(n_399),
.B2(n_391),
.C1(n_427),
.C2(n_353),
.Y(n_566)
);

OAI222xp33_ASAP7_75t_L g567 ( 
.A1(n_547),
.A2(n_454),
.B1(n_449),
.B2(n_501),
.C1(n_467),
.C2(n_491),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_521),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_522),
.A2(n_397),
.B1(n_489),
.B2(n_502),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_528),
.B(n_481),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_548),
.A2(n_489),
.B1(n_479),
.B2(n_482),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_545),
.A2(n_502),
.B(n_491),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_527),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_529),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_540),
.A2(n_431),
.B(n_452),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_524),
.A2(n_431),
.B(n_452),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_546),
.A2(n_384),
.B1(n_386),
.B2(n_376),
.Y(n_578)
);

INVx5_ASAP7_75t_SL g579 ( 
.A(n_535),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_542),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_531),
.A2(n_501),
.B1(n_449),
.B2(n_489),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_536),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_523),
.A2(n_395),
.B(n_412),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_532),
.B(n_370),
.C(n_367),
.Y(n_584)
);

OAI21xp33_ASAP7_75t_L g585 ( 
.A1(n_560),
.A2(n_349),
.B(n_373),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_561),
.A2(n_397),
.B1(n_431),
.B2(n_350),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_536),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_555),
.A2(n_490),
.B1(n_505),
.B2(n_455),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_541),
.B(n_495),
.Y(n_589)
);

BUFx4f_ASAP7_75t_SL g590 ( 
.A(n_535),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_537),
.A2(n_376),
.B1(n_350),
.B2(n_368),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_529),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_550),
.A2(n_490),
.B1(n_505),
.B2(n_454),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_537),
.A2(n_376),
.B1(n_350),
.B2(n_368),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_537),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_539),
.A2(n_350),
.B1(n_454),
.B2(n_373),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_539),
.A2(n_350),
.B1(n_359),
.B2(n_361),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_553),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_556),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_534),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_554),
.A2(n_505),
.B1(n_487),
.B2(n_498),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_541),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_539),
.A2(n_350),
.B1(n_359),
.B2(n_361),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_557),
.A2(n_497),
.B1(n_519),
.B2(n_385),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_561),
.A2(n_437),
.B1(n_444),
.B2(n_382),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_565),
.A2(n_557),
.B(n_453),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_580),
.B(n_549),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_566),
.A2(n_530),
.B1(n_561),
.B2(n_444),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_570),
.A2(n_530),
.B1(n_561),
.B2(n_437),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_564),
.A2(n_510),
.B1(n_382),
.B2(n_465),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_576),
.A2(n_500),
.B1(n_510),
.B2(n_538),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_586),
.A2(n_465),
.B1(n_558),
.B2(n_559),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_581),
.A2(n_463),
.B1(n_453),
.B2(n_469),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_596),
.B1(n_578),
.B2(n_584),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_572),
.A2(n_552),
.B1(n_497),
.B2(n_487),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_596),
.A2(n_450),
.B1(n_463),
.B2(n_469),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_579),
.A2(n_505),
.B1(n_498),
.B2(n_395),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_578),
.A2(n_469),
.B1(n_458),
.B2(n_462),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_608),
.A2(n_469),
.B1(n_458),
.B2(n_462),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_571),
.B(n_495),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_608),
.A2(n_410),
.B1(n_411),
.B2(n_416),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_603),
.A2(n_410),
.B1(n_411),
.B2(n_360),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_568),
.B(n_535),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_577),
.A2(n_370),
.B1(n_441),
.B2(n_500),
.Y(n_628)
);

AOI222xp33_ASAP7_75t_L g629 ( 
.A1(n_567),
.A2(n_388),
.B1(n_396),
.B2(n_371),
.C1(n_381),
.C2(n_374),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_569),
.A2(n_388),
.B1(n_415),
.B2(n_396),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_SL g631 ( 
.A1(n_593),
.A2(n_607),
.B1(n_583),
.B2(n_595),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_574),
.B(n_551),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_573),
.A2(n_441),
.B1(n_500),
.B2(n_457),
.Y(n_633)
);

AOI222xp33_ASAP7_75t_L g634 ( 
.A1(n_597),
.A2(n_374),
.B1(n_441),
.B2(n_387),
.C1(n_411),
.C2(n_410),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_589),
.B(n_551),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_597),
.A2(n_500),
.B1(n_544),
.B2(n_538),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_591),
.A2(n_468),
.B1(n_473),
.B2(n_538),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_579),
.A2(n_505),
.B1(n_533),
.B2(n_551),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_591),
.A2(n_538),
.B1(n_400),
.B2(n_404),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_594),
.A2(n_606),
.B1(n_587),
.B2(n_602),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_594),
.A2(n_538),
.B1(n_404),
.B2(n_398),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_606),
.A2(n_404),
.B1(n_476),
.B2(n_432),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_588),
.A2(n_544),
.B1(n_507),
.B2(n_476),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_582),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_590),
.A2(n_563),
.B1(n_595),
.B2(n_579),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_628),
.A2(n_575),
.B1(n_592),
.B2(n_590),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_615),
.B(n_605),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_632),
.B(n_599),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_610),
.B(n_589),
.C(n_563),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_600),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_L g652 ( 
.A1(n_611),
.A2(n_604),
.B1(n_600),
.B2(n_563),
.C(n_601),
.Y(n_652)
);

OA211x2_ASAP7_75t_L g653 ( 
.A1(n_646),
.A2(n_595),
.B(n_563),
.C(n_544),
.Y(n_653)
);

AND2x2_ASAP7_75t_SL g654 ( 
.A(n_633),
.B(n_595),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_599),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_618),
.B(n_631),
.C(n_609),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_624),
.B(n_645),
.Y(n_657)
);

NAND4xp25_ASAP7_75t_L g658 ( 
.A(n_627),
.B(n_533),
.C(n_404),
.D(n_476),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_SL g659 ( 
.A1(n_646),
.A2(n_533),
.B(n_504),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_644),
.B(n_598),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_614),
.B(n_598),
.Y(n_661)
);

OAI221xp5_ASAP7_75t_SL g662 ( 
.A1(n_611),
.A2(n_582),
.B1(n_436),
.B2(n_95),
.C(n_96),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_612),
.A2(n_507),
.B1(n_508),
.B2(n_474),
.C(n_436),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_630),
.B(n_508),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_639),
.B(n_507),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_613),
.B(n_508),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_630),
.B(n_508),
.C(n_474),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_619),
.B(n_641),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_508),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_637),
.B(n_474),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_638),
.B(n_474),
.Y(n_671)
);

OAI221xp5_ASAP7_75t_L g672 ( 
.A1(n_617),
.A2(n_507),
.B1(n_474),
.B2(n_436),
.C(n_445),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_623),
.B(n_92),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_655),
.Y(n_674)
);

OAI211xp5_ASAP7_75t_L g675 ( 
.A1(n_656),
.A2(n_620),
.B(n_643),
.C(n_634),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_649),
.B(n_616),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_668),
.A2(n_629),
.B1(n_622),
.B2(n_626),
.Y(n_677)
);

AO21x2_ASAP7_75t_L g678 ( 
.A1(n_669),
.A2(n_621),
.B(n_492),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_657),
.B(n_642),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_650),
.B(n_640),
.C(n_625),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_657),
.B(n_94),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_649),
.B(n_98),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_658),
.B(n_99),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_L g684 ( 
.A(n_667),
.B(n_445),
.C(n_432),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_648),
.B(n_100),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_654),
.B(n_659),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_654),
.Y(n_687)
);

AO21x2_ASAP7_75t_L g688 ( 
.A1(n_661),
.A2(n_101),
.B(n_107),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_655),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_662),
.B(n_445),
.C(n_432),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_674),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_674),
.B(n_648),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_679),
.B(n_651),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_689),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_689),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_685),
.B(n_647),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_676),
.Y(n_697)
);

XNOR2x2_ASAP7_75t_L g698 ( 
.A(n_686),
.B(n_663),
.Y(n_698)
);

XNOR2xp5_ASAP7_75t_L g699 ( 
.A(n_681),
.B(n_653),
.Y(n_699)
);

NAND4xp75_ASAP7_75t_L g700 ( 
.A(n_681),
.B(n_653),
.C(n_652),
.D(n_670),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_675),
.A2(n_670),
.B1(n_671),
.B2(n_665),
.Y(n_701)
);

XOR2x2_ASAP7_75t_L g702 ( 
.A(n_699),
.B(n_700),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_691),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_695),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_698),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_696),
.B(n_683),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_703),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_702),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_705),
.A2(n_696),
.B1(n_701),
.B2(n_680),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_707),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_708),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_711),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_709),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_715),
.A2(n_705),
.B1(n_710),
.B2(n_697),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_714),
.Y(n_717)
);

OAI22x1_ASAP7_75t_L g718 ( 
.A1(n_714),
.A2(n_710),
.B1(n_691),
.B2(n_682),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_717),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_716),
.Y(n_720)
);

OAI221xp5_ASAP7_75t_L g721 ( 
.A1(n_718),
.A2(n_713),
.B1(n_712),
.B2(n_677),
.C(n_690),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_717),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_722),
.B(n_687),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_720),
.A2(n_688),
.B1(n_678),
.B2(n_682),
.Y(n_724)
);

NOR2x1_ASAP7_75t_L g725 ( 
.A(n_721),
.B(n_688),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_719),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_722),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_719),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_727),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_726),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_728),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_729),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_725),
.B(n_693),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_723),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_724),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_725),
.A2(n_688),
.B1(n_678),
.B2(n_679),
.Y(n_737)
);

NOR4xp75_ASAP7_75t_L g738 ( 
.A(n_734),
.B(n_692),
.C(n_673),
.D(n_672),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_735),
.A2(n_687),
.B1(n_694),
.B2(n_695),
.Y(n_739)
);

OA22x2_ASAP7_75t_L g740 ( 
.A1(n_733),
.A2(n_673),
.B1(n_664),
.B2(n_671),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_678),
.B1(n_687),
.B2(n_676),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_730),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_730),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_731),
.B(n_687),
.Y(n_744)
);

NOR3xp33_ASAP7_75t_L g745 ( 
.A(n_732),
.B(n_737),
.C(n_684),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_660),
.B1(n_666),
.B2(n_687),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_743),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_740),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_745),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_741),
.B(n_666),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_738),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_739),
.Y(n_753)
);

OAI22x1_ASAP7_75t_L g754 ( 
.A1(n_747),
.A2(n_445),
.B1(n_432),
.B2(n_110),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_748),
.Y(n_755)
);

OA22x2_ASAP7_75t_L g756 ( 
.A1(n_749),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_750),
.Y(n_757)
);

AO22x2_ASAP7_75t_L g758 ( 
.A1(n_753),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_752),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_755),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_757),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_754),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_761),
.A2(n_759),
.B1(n_756),
.B2(n_751),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_762),
.A2(n_758),
.B1(n_746),
.B2(n_120),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_760),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_764),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_763),
.B1(n_765),
.B2(n_125),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_767),
.Y(n_768)
);

AOI221xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.C(n_128),
.Y(n_769)
);

AOI211xp5_ASAP7_75t_L g770 ( 
.A1(n_769),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_770)
);


endmodule