module fake_jpeg_18409_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_16),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_51),
.A2(n_18),
.B1(n_22),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_22),
.B2(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_26),
.B1(n_32),
.B2(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_32),
.B1(n_18),
.B2(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_30),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_24),
.B(n_16),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_21),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_82),
.B1(n_20),
.B2(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_17),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_27),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_43),
.B(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_29),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_23),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_101),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_107),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_98),
.B1(n_103),
.B2(n_106),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_56),
.B1(n_41),
.B2(n_46),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_23),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_23),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_108),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_41),
.B1(n_52),
.B2(n_29),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_52),
.B1(n_23),
.B2(n_3),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_1),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_23),
.B1(n_9),
.B2(n_10),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_67),
.B1(n_71),
.B2(n_81),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_64),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_60),
.B(n_80),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_123),
.B(n_127),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_86),
.B(n_84),
.C(n_82),
.D(n_60),
.Y(n_123)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_86),
.C(n_88),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_107),
.C(n_96),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_87),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_72),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_74),
.B1(n_73),
.B2(n_69),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_98),
.B1(n_93),
.B2(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_137),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_71),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_93),
.B(n_89),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_73),
.B1(n_69),
.B2(n_71),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_101),
.B1(n_112),
.B2(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_78),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_9),
.B(n_13),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_7),
.B(n_13),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_96),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_119),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_152),
.B(n_161),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_97),
.B1(n_107),
.B2(n_92),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_107),
.B1(n_97),
.B2(n_109),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_165),
.B1(n_128),
.B2(n_134),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_107),
.B(n_115),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_169),
.C(n_171),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_163),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_110),
.B(n_96),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_72),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_74),
.B1(n_113),
.B2(n_9),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_114),
.B(n_3),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_135),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_8),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_123),
.A2(n_127),
.B(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_119),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_117),
.B(n_8),
.Y(n_171)
);

AOI22x1_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_172)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_122),
.B1(n_132),
.B2(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_186),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2x1_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_138),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_145),
.B1(n_150),
.B2(n_188),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_157),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_182),
.B(n_183),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_141),
.C(n_117),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_191),
.C(n_169),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_160),
.B1(n_165),
.B2(n_147),
.Y(n_205)
);

BUFx12f_ASAP7_75t_SL g189 ( 
.A(n_168),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_131),
.C(n_125),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

NAND5xp2_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_120),
.C(n_139),
.D(n_116),
.E(n_140),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_174),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_194),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_160),
.B1(n_153),
.B2(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_152),
.B1(n_159),
.B2(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_179),
.A2(n_159),
.B1(n_148),
.B2(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_148),
.B1(n_171),
.B2(n_161),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_214),
.C(n_178),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_136),
.C(n_120),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_196),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_191),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_224),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_178),
.C(n_184),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_230),
.C(n_218),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_210),
.A2(n_185),
.B1(n_189),
.B2(n_176),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_201),
.B1(n_200),
.B2(n_215),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_210),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_202),
.C(n_209),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_240),
.Y(n_247)
);

XOR2x1_ASAP7_75t_SL g237 ( 
.A(n_230),
.B(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_239),
.A2(n_244),
.B1(n_222),
.B2(n_204),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_199),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_198),
.B(n_173),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_180),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_190),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_175),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_250),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_225),
.B(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_195),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_253),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_242),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_256),
.B(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_242),
.C(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_263),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_243),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_243),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_6),
.B(n_12),
.Y(n_269)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_250),
.B(n_246),
.Y(n_265)
);

OAI321xp33_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_266),
.A3(n_267),
.B1(n_14),
.B2(n_4),
.C(n_2),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_247),
.C(n_3),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_269),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_2),
.B(n_3),
.Y(n_274)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_262),
.B1(n_5),
.B2(n_11),
.C(n_14),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_265),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_276),
.A2(n_272),
.B(n_2),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_275),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_4),
.Y(n_279)
);


endmodule