module real_aes_9594_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_102;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_397;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_0), .A2(n_3), .B1(n_623), .B2(n_625), .C(n_629), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_0), .A2(n_3), .B1(n_649), .B2(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_1), .B(n_194), .Y(n_219) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_2), .Y(n_594) );
INVx1_ASAP7_75t_L g621 ( .A(n_2), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_4), .A2(n_72), .B1(n_487), .B2(n_497), .Y(n_486) );
INVx1_ASAP7_75t_L g607 ( .A(n_4), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_5), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_6), .B(n_162), .Y(n_218) );
INVx2_ASAP7_75t_L g491 ( .A(n_7), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_8), .A2(n_70), .B1(n_579), .B2(n_584), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_8), .A2(n_70), .B1(n_649), .B2(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g539 ( .A(n_9), .Y(n_539) );
BUFx2_ASAP7_75t_L g591 ( .A(n_9), .Y(n_591) );
INVx1_ASAP7_75t_L g619 ( .A(n_9), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_10), .B(n_179), .Y(n_243) );
INVx1_ASAP7_75t_L g686 ( .A(n_10), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_11), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_12), .B(n_157), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_13), .B(n_140), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_14), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_15), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_15), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_16), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_17), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_18), .B(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_19), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_20), .B(n_157), .Y(n_163) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_21), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_22), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_23), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_24), .B(n_124), .Y(n_144) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_25), .A2(n_517), .B(n_521), .C(n_526), .Y(n_516) );
INVx1_ASAP7_75t_L g610 ( .A(n_25), .Y(n_610) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_26), .Y(n_674) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_27), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_28), .B(n_140), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_29), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g537 ( .A(n_30), .Y(n_537) );
INVx1_ASAP7_75t_L g708 ( .A(n_30), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_31), .Y(n_632) );
NAND2xp33_ASAP7_75t_SL g122 ( .A(n_32), .B(n_91), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_33), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_34), .B(n_118), .Y(n_242) );
OAI21x1_ASAP7_75t_L g112 ( .A1(n_35), .A2(n_53), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_36), .B(n_166), .Y(n_182) );
AND2x6_ASAP7_75t_L g84 ( .A(n_37), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_37), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_37), .B(n_662), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_38), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_39), .B(n_109), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_40), .B(n_109), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_41), .B(n_176), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_42), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_43), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_44), .A2(n_48), .B1(n_502), .B2(n_510), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_44), .A2(n_72), .B1(n_597), .B2(n_603), .C(n_606), .Y(n_596) );
INVx1_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_45), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_46), .B(n_191), .Y(n_190) );
NAND2xp33_ASAP7_75t_L g119 ( .A(n_47), .B(n_91), .Y(n_119) );
INVx1_ASAP7_75t_L g570 ( .A(n_48), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_49), .B(n_124), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_50), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_51), .B(n_192), .Y(n_203) );
INVx2_ASAP7_75t_L g551 ( .A(n_52), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_54), .B(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_54), .Y(n_710) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_55), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_56), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_57), .B(n_166), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_58), .Y(n_531) );
BUFx10_ASAP7_75t_L g702 ( .A(n_59), .Y(n_702) );
INVx1_ASAP7_75t_L g554 ( .A(n_60), .Y(n_554) );
INVx2_ASAP7_75t_L g563 ( .A(n_60), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_61), .B(n_140), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_62), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_63), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_64), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_65), .B(n_157), .Y(n_174) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_65), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_66), .Y(n_534) );
INVx2_ASAP7_75t_L g113 ( .A(n_67), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_68), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_69), .B(n_138), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_71), .B(n_179), .Y(n_207) );
INVx2_ASAP7_75t_L g549 ( .A(n_73), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_74), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_75), .Y(n_543) );
INVx1_ASAP7_75t_L g494 ( .A(n_76), .Y(n_494) );
BUFx3_ASAP7_75t_L g500 ( .A(n_76), .Y(n_500) );
INVx1_ASAP7_75t_L g496 ( .A(n_77), .Y(n_496) );
BUFx3_ASAP7_75t_L g509 ( .A(n_77), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_96), .B(n_480), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx2_ASAP7_75t_SL g127 ( .A(n_83), .Y(n_127) );
INVx8_ASAP7_75t_L g145 ( .A(n_83), .Y(n_145) );
INVx8_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_84), .A2(n_173), .B(n_177), .Y(n_172) );
OAI21x1_ASAP7_75t_SL g200 ( .A1(n_84), .A2(n_201), .B(n_204), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_84), .A2(n_126), .B(n_213), .C(n_216), .Y(n_212) );
INVxp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AO21x1_ASAP7_75t_L g720 ( .A1(n_87), .A2(n_721), .B(n_722), .Y(n_720) );
NAND2xp33_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g206 ( .A(n_91), .Y(n_206) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g118 ( .A(n_92), .Y(n_118) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_92), .Y(n_125) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
INVx1_ASAP7_75t_L g180 ( .A(n_92), .Y(n_180) );
BUFx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_94), .A2(n_205), .B(n_207), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_94), .A2(n_217), .B(n_218), .Y(n_216) );
BUFx12f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx5_ASAP7_75t_L g120 ( .A(n_95), .Y(n_120) );
INVx5_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_359), .Y(n_99) );
NOR3xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_289), .C(n_330), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_102), .B(n_272), .Y(n_101) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_169), .B1(n_220), .B2(n_223), .C(n_256), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_129), .Y(n_104) );
INVx1_ASAP7_75t_L g271 ( .A(n_105), .Y(n_271) );
INVx1_ASAP7_75t_L g285 ( .A(n_105), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_105), .B(n_259), .Y(n_358) );
INVx1_ASAP7_75t_L g410 ( .A(n_105), .Y(n_410) );
AND2x2_ASAP7_75t_L g459 ( .A(n_105), .B(n_349), .Y(n_459) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g261 ( .A(n_106), .B(n_222), .Y(n_261) );
AND2x2_ASAP7_75t_L g452 ( .A(n_106), .B(n_400), .Y(n_452) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_107), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_107), .B(n_222), .Y(n_336) );
INVx2_ASAP7_75t_L g365 ( .A(n_107), .Y(n_365) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g250 ( .A(n_108), .B(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_108), .Y(n_429) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_114), .B(n_128), .Y(n_108) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_109), .A2(n_172), .B(n_182), .Y(n_171) );
INVx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g209 ( .A(n_110), .Y(n_209) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx5_ASAP7_75t_L g134 ( .A(n_111), .Y(n_134) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g168 ( .A(n_112), .Y(n_168) );
OAI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_121), .B(n_127), .Y(n_114) );
O2A1O1Ixp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B(n_119), .C(n_120), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g213 ( .A1(n_118), .A2(n_140), .B1(n_214), .B2(n_215), .Y(n_213) );
INVx2_ASAP7_75t_SL g126 ( .A(n_120), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_120), .A2(n_137), .B(n_139), .Y(n_136) );
INVx2_ASAP7_75t_SL g158 ( .A(n_120), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_120), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B(n_126), .Y(n_121) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
INVx2_ASAP7_75t_L g155 ( .A(n_125), .Y(n_155) );
INVx2_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_126), .A2(n_142), .B(n_144), .Y(n_141) );
AOI21x1_ASAP7_75t_L g188 ( .A1(n_126), .A2(n_189), .B(n_190), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_127), .A2(n_153), .B(n_159), .Y(n_152) );
OAI21x1_ASAP7_75t_L g184 ( .A1(n_127), .A2(n_185), .B(n_188), .Y(n_184) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_130), .B(n_250), .Y(n_296) );
INVx1_ASAP7_75t_L g320 ( .A(n_130), .Y(n_320) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_130), .Y(n_369) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_130), .B(n_348), .Y(n_411) );
AND2x2_ASAP7_75t_L g456 ( .A(n_130), .B(n_398), .Y(n_456) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_148), .Y(n_130) );
INVx3_ASAP7_75t_L g357 ( .A(n_131), .Y(n_357) );
BUFx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g282 ( .A(n_132), .Y(n_282) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g222 ( .A(n_133), .Y(n_222) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_146), .Y(n_133) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_134), .A2(n_152), .B(n_165), .Y(n_151) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_134), .A2(n_212), .B(n_219), .Y(n_211) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_134), .A2(n_237), .B(n_244), .Y(n_236) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .B(n_145), .Y(n_135) );
OAI21x1_ASAP7_75t_L g237 ( .A1(n_145), .A2(n_238), .B(n_241), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_148), .B(n_300), .Y(n_378) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_149), .B(n_282), .Y(n_366) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g269 ( .A(n_150), .Y(n_269) );
AND2x2_ASAP7_75t_L g326 ( .A(n_150), .B(n_235), .Y(n_326) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g260 ( .A(n_151), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_158), .Y(n_153) );
INVx5_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_158), .A2(n_178), .B(n_181), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_158), .A2(n_239), .B(n_240), .Y(n_238) );
O2A1O1Ixp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_163), .C(n_164), .Y(n_159) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_174), .B(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_164), .A2(n_179), .B(n_202), .C(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_164), .A2(n_242), .B(n_243), .Y(n_241) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_168), .Y(n_194) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_196), .Y(n_169) );
INVx2_ASAP7_75t_L g262 ( .A(n_170), .Y(n_262) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_170), .Y(n_313) );
AND2x2_ASAP7_75t_L g338 ( .A(n_170), .B(n_278), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_170), .B(n_353), .Y(n_432) );
AND2x2_ASAP7_75t_L g435 ( .A(n_170), .B(n_387), .Y(n_435) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_183), .Y(n_170) );
INVx2_ASAP7_75t_L g228 ( .A(n_171), .Y(n_228) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g192 ( .A(n_180), .Y(n_192) );
BUFx2_ASAP7_75t_L g275 ( .A(n_183), .Y(n_275) );
AND2x2_ASAP7_75t_L g294 ( .A(n_183), .B(n_228), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_193), .B(n_195), .Y(n_183) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_184), .A2(n_193), .B(n_195), .Y(n_231) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_200), .B(n_208), .Y(n_199) );
BUFx2_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_197), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_210), .Y(n_197) );
INVx1_ASAP7_75t_L g227 ( .A(n_198), .Y(n_227) );
INVx2_ASAP7_75t_SL g255 ( .A(n_198), .Y(n_255) );
AND2x2_ASAP7_75t_L g316 ( .A(n_198), .B(n_228), .Y(n_316) );
AND2x2_ASAP7_75t_L g387 ( .A(n_198), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g416 ( .A(n_198), .Y(n_416) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_198), .Y(n_439) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g303 ( .A(n_199), .B(n_211), .Y(n_303) );
AND2x2_ASAP7_75t_L g229 ( .A(n_210), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g278 ( .A(n_210), .B(n_255), .Y(n_278) );
AND2x2_ASAP7_75t_L g310 ( .A(n_210), .B(n_282), .Y(n_310) );
INVx1_ASAP7_75t_L g388 ( .A(n_210), .Y(n_388) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g266 ( .A(n_211), .B(n_230), .Y(n_266) );
INVx2_ASAP7_75t_L g329 ( .A(n_211), .Y(n_329) );
BUFx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_221), .B(n_260), .Y(n_350) );
INVx2_ASAP7_75t_L g474 ( .A(n_221), .Y(n_474) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OAI221xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_232), .B1(n_245), .B2(n_249), .C(n_252), .Y(n_223) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_224), .A2(n_469), .B1(n_472), .B2(n_475), .C(n_477), .Y(n_471) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_229), .Y(n_225) );
NOR2xp67_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_227), .Y(n_404) );
AND2x2_ASAP7_75t_L g254 ( .A(n_228), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
INVx1_ASAP7_75t_L g395 ( .A(n_228), .Y(n_395) );
INVx1_ASAP7_75t_L g414 ( .A(n_228), .Y(n_414) );
AND2x2_ASAP7_75t_L g253 ( .A(n_229), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g318 ( .A(n_229), .Y(n_318) );
INVx2_ASAP7_75t_SL g248 ( .A(n_230), .Y(n_248) );
AND2x4_ASAP7_75t_L g394 ( .A(n_230), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVxp67_ASAP7_75t_R g346 ( .A(n_231), .Y(n_346) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_233), .A2(n_320), .B(n_437), .C(n_478), .Y(n_477) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g428 ( .A(n_234), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g251 ( .A(n_235), .Y(n_251) );
AND2x2_ASAP7_75t_L g284 ( .A(n_235), .B(n_269), .Y(n_284) );
INVx1_ASAP7_75t_L g300 ( .A(n_235), .Y(n_300) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_245), .Y(n_354) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g381 ( .A(n_248), .B(n_316), .Y(n_381) );
NAND4xp25_ASAP7_75t_SL g407 ( .A(n_249), .B(n_385), .C(n_408), .D(n_411), .Y(n_407) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_250), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_250), .B(n_268), .Y(n_464) );
INVx1_ASAP7_75t_L g400 ( .A(n_251), .Y(n_400) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g265 ( .A(n_254), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g328 ( .A(n_254), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g342 ( .A(n_254), .B(n_343), .Y(n_342) );
OAI32xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_262), .A3(n_263), .B1(n_264), .B2(n_267), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_258), .A2(n_298), .B(n_301), .Y(n_297) );
AND2x4_ASAP7_75t_SL g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g409 ( .A(n_259), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g373 ( .A(n_261), .B(n_299), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_263), .A2(n_273), .B1(n_279), .B2(n_286), .Y(n_272) );
INVx1_ASAP7_75t_L g457 ( .A(n_263), .Y(n_457) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
O2A1O1Ixp5_ASAP7_75t_SL g443 ( .A1(n_265), .A2(n_444), .B(n_446), .C(n_450), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g299 ( .A(n_269), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_269), .Y(n_334) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g377 ( .A(n_271), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g343 ( .A(n_275), .Y(n_343) );
AND2x2_ASAP7_75t_L g415 ( .A(n_275), .B(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x6_ASAP7_75t_L g292 ( .A(n_277), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g370 ( .A(n_278), .B(n_346), .Y(n_370) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g286 ( .A(n_281), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g298 ( .A(n_281), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g325 ( .A(n_281), .B(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_283), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g418 ( .A(n_283), .Y(n_418) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g287 ( .A(n_284), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
AND2x2_ASAP7_75t_L g323 ( .A(n_288), .B(n_299), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_307), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B(n_297), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g431 ( .A(n_299), .Y(n_431) );
BUFx2_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_303), .B(n_305), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_303), .A2(n_455), .B1(n_457), .B2(n_458), .Y(n_454) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI221xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_313), .B1(n_314), .B2(n_319), .C(n_321), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_311), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g385 ( .A(n_312), .B(n_357), .Y(n_385) );
INVx1_ASAP7_75t_L g470 ( .A(n_312), .Y(n_470) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp33_ASAP7_75t_SL g463 ( .A1(n_315), .A2(n_445), .B1(n_464), .B2(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g345 ( .A(n_316), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g352 ( .A(n_316), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g476 ( .A(n_316), .Y(n_476) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B(n_327), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g382 ( .A(n_323), .Y(n_382) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g441 ( .A(n_326), .B(n_410), .Y(n_441) );
INVx1_ASAP7_75t_L g449 ( .A(n_326), .Y(n_449) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx4_ASAP7_75t_L g353 ( .A(n_329), .Y(n_353) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_329), .B(n_394), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_337), .B(n_339), .C(n_351), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_331), .A2(n_397), .B(n_401), .C(n_403), .Y(n_396) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g391 ( .A(n_336), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_337), .A2(n_420), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
AND2x2_ASAP7_75t_L g386 ( .A(n_343), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g465 ( .A(n_345), .Y(n_465) );
AND2x2_ASAP7_75t_L g438 ( .A(n_346), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g420 ( .A(n_350), .B(n_364), .Y(n_420) );
INVx1_ASAP7_75t_L g426 ( .A(n_350), .Y(n_426) );
OAI21xp33_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_354), .B(n_355), .Y(n_351) );
INVx1_ASAP7_75t_L g376 ( .A(n_353), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_353), .B(n_394), .Y(n_421) );
OR2x2_ASAP7_75t_L g475 ( .A(n_353), .B(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g445 ( .A(n_357), .B(n_399), .Y(n_445) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_357), .B(n_449), .Y(n_448) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_442), .Y(n_359) );
NAND4xp25_ASAP7_75t_L g360 ( .A(n_361), .B(n_383), .C(n_406), .D(n_422), .Y(n_360) );
O2A1O1Ixp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_367), .B(n_370), .C(n_371), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
OR2x2_ASAP7_75t_L g430 ( .A(n_364), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g478 ( .A(n_364), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g399 ( .A(n_365), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
INVx1_ASAP7_75t_L g479 ( .A(n_366), .Y(n_479) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
OAI322xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .A3(n_376), .B1(n_377), .B2(n_379), .C1(n_380), .C2(n_382), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g467 ( .A(n_376), .B(n_381), .Y(n_467) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B1(n_389), .B2(n_392), .C(n_396), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g419 ( .A(n_386), .Y(n_419) );
AND2x2_ASAP7_75t_L g413 ( .A(n_388), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g405 ( .A(n_394), .Y(n_405) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_412), .B(n_417), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_413), .B(n_415), .Y(n_424) );
AND2x4_ASAP7_75t_L g437 ( .A(n_413), .B(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_433), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_430), .B2(n_432), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_453), .C(n_466), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp67_ASAP7_75t_SL g473 ( .A(n_452), .B(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_460), .B(n_463), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_471), .Y(n_466) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B1(n_660), .B2(n_665), .C(n_715), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_483), .A2(n_710), .B1(n_716), .B2(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND3x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_540), .C(n_595), .Y(n_484) );
OAI31xp33_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_501), .A3(n_516), .B(n_535), .Y(n_485) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_492), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x6_ASAP7_75t_L g498 ( .A(n_489), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g523 ( .A(n_489), .Y(n_523) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x6_ASAP7_75t_L g532 ( .A(n_490), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_491), .Y(n_505) );
INVx1_ASAP7_75t_L g513 ( .A(n_491), .Y(n_513) );
AND2x2_ASAP7_75t_L g642 ( .A(n_491), .B(n_537), .Y(n_642) );
INVx2_ASAP7_75t_L g654 ( .A(n_491), .Y(n_654) );
INVx2_ASAP7_75t_L g645 ( .A(n_492), .Y(n_645) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g520 ( .A(n_493), .B(n_495), .Y(n_520) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g515 ( .A(n_494), .B(n_509), .Y(n_515) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g499 ( .A(n_496), .B(n_500), .Y(n_499) );
CKINVDCx6p67_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_499), .Y(n_649) );
INVx2_ASAP7_75t_L g507 ( .A(n_500), .Y(n_507) );
AND2x2_ASAP7_75t_L g525 ( .A(n_500), .B(n_509), .Y(n_525) );
INVx4_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
AND2x4_ASAP7_75t_L g527 ( .A(n_504), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g533 ( .A(n_507), .Y(n_533) );
INVx1_ASAP7_75t_L g530 ( .A(n_508), .Y(n_530) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_514), .Y(n_650) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_515), .Y(n_659) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g647 ( .A(n_520), .Y(n_647) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_520), .Y(n_657) );
CKINVDCx8_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_531), .B1(n_532), .B2(n_534), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g700 ( .A(n_530), .Y(n_700) );
AOI222xp33_ASAP7_75t_SL g542 ( .A1(n_531), .A2(n_534), .B1(n_543), .B2(n_544), .C1(n_552), .C2(n_556), .Y(n_542) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g653 ( .A(n_537), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g637 ( .A(n_539), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_578), .B(n_589), .Y(n_540) );
NAND3xp33_ASAP7_75t_SL g541 ( .A(n_542), .B(n_564), .C(n_575), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_543), .A2(n_565), .B1(n_644), .B2(n_656), .C(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g576 ( .A(n_547), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g559 ( .A(n_549), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_549), .B(n_551), .Y(n_569) );
INVx2_ASAP7_75t_L g583 ( .A(n_549), .Y(n_583) );
AND2x4_ASAP7_75t_L g588 ( .A(n_549), .B(n_550), .Y(n_588) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g555 ( .A(n_551), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_551), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g602 ( .A(n_551), .Y(n_602) );
INVx1_ASAP7_75t_L g615 ( .A(n_551), .Y(n_615) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
OR2x6_ASAP7_75t_L g567 ( .A(n_553), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g638 ( .A(n_554), .B(n_593), .Y(n_638) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_559), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g634 ( .A(n_559), .B(n_615), .Y(n_634) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g577 ( .A(n_561), .Y(n_577) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_562), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g574 ( .A(n_563), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_570), .B2(n_571), .Y(n_564) );
INVx8_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x6_ASAP7_75t_L g572 ( .A(n_568), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_SL g609 ( .A(n_568), .Y(n_609) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_568), .Y(n_631) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx4_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g580 ( .A(n_573), .Y(n_580) );
AND2x4_ASAP7_75t_L g585 ( .A(n_573), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx11_ASAP7_75t_R g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
BUFx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g600 ( .A(n_583), .B(n_601), .Y(n_600) );
INVx5_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_588), .Y(n_605) );
INVx3_ASAP7_75t_L g628 ( .A(n_588), .Y(n_628) );
CKINVDCx16_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
OR2x6_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x4_ASAP7_75t_L g652 ( .A(n_591), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_616), .B1(n_622), .B2(n_635), .C(n_639), .Y(n_595) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g624 ( .A(n_600), .Y(n_624) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_610), .B2(n_611), .Y(n_606) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx6_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x6_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_630), .A2(n_632), .B1(n_644), .B2(n_646), .C(n_648), .Y(n_643) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OR2x2_ASAP7_75t_L g640 ( .A(n_637), .B(n_641), .Y(n_640) );
OAI22xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_643), .B1(n_651), .B2(n_655), .Y(n_639) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_SL g696 ( .A(n_642), .Y(n_696) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx4_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g706 ( .A(n_654), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_662), .B(n_664), .Y(n_692) );
INVx1_ASAP7_75t_SL g721 ( .A(n_662), .Y(n_721) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_689), .B1(n_710), .B2(n_711), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_666), .A2(n_710), .B1(n_717), .B2(n_718), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_678), .B1(n_679), .B2(n_688), .Y(n_666) );
INVx1_ASAP7_75t_L g688 ( .A(n_667), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_676), .B2(n_677), .Y(n_667) );
CKINVDCx16_ASAP7_75t_R g676 ( .A(n_668), .Y(n_676) );
XOR2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g677 ( .A(n_671), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_672), .Y(n_675) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_679) );
INVx1_ASAP7_75t_L g687 ( .A(n_680), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_683), .B2(n_684), .Y(n_680) );
INVx4_ASAP7_75t_L g684 ( .A(n_681), .Y(n_684) );
INVx1_ASAP7_75t_L g683 ( .A(n_682), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_691), .Y(n_717) );
OR2x6_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
OR2x4_ASAP7_75t_L g714 ( .A(n_692), .B(n_694), .Y(n_714) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI31xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .A3(n_701), .B(n_703), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g709 ( .A(n_700), .Y(n_709) );
INVx6_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx5_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx8_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g718 ( .A(n_713), .Y(n_718) );
INVx8_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx3_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
endmodule