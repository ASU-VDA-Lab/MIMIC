module fake_jpeg_20160_n_31 (n_3, n_2, n_1, n_0, n_4, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_SL g6 ( 
.A(n_1),
.B(n_5),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx4f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_14),
.B1(n_15),
.B2(n_11),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_7),
.B1(n_14),
.B2(n_8),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_21),
.B1(n_16),
.B2(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_9),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.C(n_24),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_11),
.B(n_10),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_9),
.C(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_10),
.B(n_3),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_28),
.B(n_4),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_9),
.Y(n_31)
);


endmodule