module fake_jpeg_11385_n_183 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_10),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_21),
.Y(n_56)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_44),
.B1(n_23),
.B2(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_20),
.Y(n_53)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_56),
.B(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_15),
.Y(n_61)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_21),
.CON(n_66),
.SN(n_66)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_19),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_47),
.B1(n_37),
.B2(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_88),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_91),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_27),
.B1(n_17),
.B2(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_16),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_40),
.B1(n_34),
.B2(n_17),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_67),
.A3(n_66),
.B1(n_70),
.B2(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_27),
.B1(n_45),
.B2(n_30),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_55),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_16),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_16),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_70),
.C(n_40),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_109),
.C(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_11),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_122),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_109),
.B1(n_99),
.B2(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_131),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_8),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_14),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_77),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_109),
.B(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_130),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_127),
.B1(n_122),
.B2(n_125),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_145),
.B1(n_75),
.B2(n_73),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_103),
.B(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_118),
.B(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_75),
.B1(n_97),
.B2(n_64),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_119),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_97),
.C(n_91),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_150),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_151),
.B1(n_139),
.B2(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_103),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_143),
.B1(n_132),
.B2(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_4),
.C(n_5),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_146),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_142),
.A3(n_141),
.B1(n_145),
.B2(n_7),
.C1(n_2),
.C2(n_1),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_152),
.B1(n_154),
.B2(n_148),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_142),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_164),
.B1(n_160),
.B2(n_3),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_150),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_159),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_1),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_171),
.B(n_174),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_177),
.C(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_2),
.Y(n_183)
);


endmodule