module real_aes_7673_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_1), .A2(n_150), .B(n_155), .C(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_2), .A2(n_145), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g462 ( .A(n_3), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_4), .A2(n_104), .B1(n_118), .B2(n_736), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_5), .B(n_169), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_6), .A2(n_16), .B1(n_724), .B2(n_725), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_6), .Y(n_725) );
AOI21xp33_ASAP7_75t_L g479 ( .A1(n_7), .A2(n_145), .B(n_480), .Y(n_479) );
AND2x6_ASAP7_75t_L g150 ( .A(n_8), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g179 ( .A(n_9), .Y(n_179) );
INVx1_ASAP7_75t_L g110 ( .A(n_10), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_10), .B(n_44), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_11), .A2(n_257), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_12), .B(n_160), .Y(n_196) );
INVx1_ASAP7_75t_L g484 ( .A(n_13), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_14), .B(n_159), .Y(n_532) );
INVx1_ASAP7_75t_L g143 ( .A(n_15), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_16), .Y(n_724) );
INVx1_ASAP7_75t_L g544 ( .A(n_17), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_18), .A2(n_180), .B(n_205), .C(n_207), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_19), .B(n_169), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_20), .B(n_473), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_21), .B(n_145), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_22), .B(n_265), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_23), .A2(n_159), .B(n_161), .C(n_165), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_24), .B(n_169), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_25), .B(n_160), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_26), .A2(n_163), .B(n_207), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_27), .B(n_160), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_28), .Y(n_225) );
INVx1_ASAP7_75t_L g239 ( .A(n_29), .Y(n_239) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_30), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_31), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_32), .B(n_160), .Y(n_463) );
INVx1_ASAP7_75t_L g262 ( .A(n_33), .Y(n_262) );
INVx1_ASAP7_75t_L g497 ( .A(n_34), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_35), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g148 ( .A(n_36), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_37), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_38), .A2(n_159), .B(n_218), .C(n_220), .Y(n_217) );
INVxp67_ASAP7_75t_L g263 ( .A(n_39), .Y(n_263) );
CKINVDCx14_ASAP7_75t_R g216 ( .A(n_40), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_41), .A2(n_155), .B(n_238), .C(n_244), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_42), .A2(n_150), .B(n_155), .C(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_43), .A2(n_92), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_43), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_44), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g496 ( .A(n_45), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_46), .A2(n_177), .B(n_178), .C(n_181), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_47), .B(n_160), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_48), .A2(n_126), .B1(n_438), .B2(n_439), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_48), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_49), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_50), .Y(n_259) );
INVx1_ASAP7_75t_L g153 ( .A(n_51), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_52), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_53), .B(n_145), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_54), .A2(n_155), .B1(n_165), .B2(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_55), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_56), .Y(n_459) );
CKINVDCx14_ASAP7_75t_R g175 ( .A(n_57), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_58), .A2(n_177), .B(n_220), .C(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_59), .Y(n_525) );
INVx1_ASAP7_75t_L g481 ( .A(n_60), .Y(n_481) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
INVx1_ASAP7_75t_L g142 ( .A(n_62), .Y(n_142) );
INVx1_ASAP7_75t_SL g219 ( .A(n_63), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_64), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_65), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g228 ( .A(n_66), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_SL g472 ( .A1(n_67), .A2(n_220), .B(n_473), .C(n_474), .Y(n_472) );
INVxp67_ASAP7_75t_L g475 ( .A(n_68), .Y(n_475) );
INVx1_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_70), .A2(n_145), .B(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_71), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_72), .A2(n_145), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_73), .Y(n_500) );
INVx1_ASAP7_75t_L g519 ( .A(n_74), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_75), .A2(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g203 ( .A(n_76), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_77), .Y(n_236) );
AOI222xp33_ASAP7_75t_L g449 ( .A1(n_78), .A2(n_450), .B1(n_721), .B2(n_727), .C1(n_731), .C2(n_732), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_79), .A2(n_150), .B(n_155), .C(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_80), .A2(n_145), .B(n_152), .Y(n_144) );
INVx1_ASAP7_75t_L g206 ( .A(n_81), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_82), .B(n_240), .Y(n_513) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
INVx1_ASAP7_75t_L g193 ( .A(n_84), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_85), .B(n_473), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_86), .A2(n_150), .B(n_155), .C(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g114 ( .A(n_87), .Y(n_114) );
OR2x2_ASAP7_75t_L g442 ( .A(n_87), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g720 ( .A(n_87), .B(n_444), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_88), .A2(n_155), .B(n_227), .C(n_230), .Y(n_226) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_89), .A2(n_722), .B1(n_723), .B2(n_726), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_89), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_90), .B(n_172), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_91), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_92), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_93), .A2(n_150), .B(n_155), .C(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_94), .Y(n_536) );
INVx1_ASAP7_75t_L g471 ( .A(n_95), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_96), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_97), .B(n_240), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_98), .B(n_138), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_99), .B(n_138), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_100), .B(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g162 ( .A(n_101), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_102), .A2(n_145), .B(n_470), .Y(n_469) );
BUFx4f_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g736 ( .A(n_107), .Y(n_736) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g444 ( .A(n_113), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g719 ( .A(n_114), .B(n_444), .Y(n_719) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_114), .B(n_443), .Y(n_734) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
AO21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_448), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g735 ( .A(n_121), .Y(n_735) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_440), .B(n_446), .Y(n_124) );
INVx1_ASAP7_75t_L g439 ( .A(n_126), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_436), .B2(n_437), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_127), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_130), .A2(n_719), .B1(n_728), .B2(n_729), .Y(n_727) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g437 ( .A(n_131), .Y(n_437) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_362), .Y(n_131) );
NOR4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_304), .C(n_334), .D(n_344), .Y(n_132) );
OAI211xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_209), .B(n_267), .C(n_294), .Y(n_133) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_134), .A2(n_309), .B1(n_390), .B2(n_391), .C1(n_392), .C2(n_393), .Y(n_389) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_184), .Y(n_134) );
AOI33xp33_ASAP7_75t_L g315 ( .A1(n_135), .A2(n_302), .A3(n_303), .B1(n_316), .B2(n_321), .B3(n_323), .Y(n_315) );
OAI211xp5_ASAP7_75t_SL g372 ( .A1(n_135), .A2(n_373), .B(n_375), .C(n_377), .Y(n_372) );
OR2x2_ASAP7_75t_L g388 ( .A(n_135), .B(n_374), .Y(n_388) );
INVx1_ASAP7_75t_L g421 ( .A(n_135), .Y(n_421) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_171), .Y(n_135) );
INVx2_ASAP7_75t_L g298 ( .A(n_136), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_136), .B(n_200), .Y(n_314) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_136), .Y(n_349) );
AND2x2_ASAP7_75t_L g378 ( .A(n_136), .B(n_171), .Y(n_378) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_168), .Y(n_136) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_137), .A2(n_201), .B(n_208), .Y(n_200) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_137), .A2(n_214), .B(n_222), .Y(n_213) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_138), .A2(n_469), .B(n_476), .Y(n_468) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g255 ( .A(n_139), .Y(n_255) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_140), .B(n_141), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g257 ( .A(n_145), .Y(n_257) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_146), .B(n_150), .Y(n_190) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g243 ( .A(n_147), .Y(n_243) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
INVx1_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
INVx1_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
INVx3_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
INVx1_ASAP7_75t_L g473 ( .A(n_149), .Y(n_473) );
INVx4_ASAP7_75t_SL g167 ( .A(n_150), .Y(n_167) );
BUFx3_ASAP7_75t_L g244 ( .A(n_150), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g152 ( .A1(n_153), .A2(n_154), .B(n_158), .C(n_167), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_154), .A2(n_167), .B(n_175), .C(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_154), .A2(n_167), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_154), .A2(n_167), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_154), .A2(n_167), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_154), .A2(n_167), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_154), .A2(n_167), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_154), .A2(n_167), .B(n_541), .C(n_542), .Y(n_540) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx3_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_156), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_159), .B(n_219), .Y(n_218) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_163), .B(n_206), .Y(n_205) );
OAI22xp33_ASAP7_75t_L g261 ( .A1(n_163), .A2(n_240), .B1(n_262), .B2(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_163), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_164), .A2(n_195), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g464 ( .A(n_165), .Y(n_464) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g230 ( .A(n_167), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_167), .A2(n_190), .B1(n_494), .B2(n_498), .Y(n_493) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_169), .A2(n_479), .B(n_485), .Y(n_478) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_170), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_170), .A2(n_224), .B(n_231), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_170), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_SL g515 ( .A(n_170), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g278 ( .A(n_171), .Y(n_278) );
BUFx3_ASAP7_75t_L g286 ( .A(n_171), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_171), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g297 ( .A(n_171), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_171), .B(n_185), .Y(n_326) );
AND2x2_ASAP7_75t_L g395 ( .A(n_171), .B(n_329), .Y(n_395) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_183), .Y(n_171) );
INVx1_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
INVx2_ASAP7_75t_L g233 ( .A(n_172), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_172), .A2(n_190), .B(n_236), .C(n_237), .Y(n_235) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_172), .A2(n_539), .B(n_545), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx5_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_180), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_180), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g197 ( .A(n_181), .Y(n_197) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g207 ( .A(n_182), .Y(n_207) );
INVx2_ASAP7_75t_SL g289 ( .A(n_184), .Y(n_289) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_185), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g331 ( .A(n_185), .Y(n_331) );
AND2x2_ASAP7_75t_L g342 ( .A(n_185), .B(n_298), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_185), .B(n_327), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_185), .B(n_329), .Y(n_374) );
AND2x2_ASAP7_75t_L g433 ( .A(n_185), .B(n_378), .Y(n_433) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g303 ( .A(n_186), .B(n_200), .Y(n_303) );
AND2x2_ASAP7_75t_L g313 ( .A(n_186), .B(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g335 ( .A(n_186), .Y(n_335) );
AND3x2_ASAP7_75t_L g394 ( .A(n_186), .B(n_395), .C(n_396), .Y(n_394) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_198), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_187), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_187), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_187), .B(n_536), .Y(n_535) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_190), .A2(n_225), .B(n_226), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_190), .A2(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_190), .A2(n_519), .B(n_520), .Y(n_518) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_197), .B(n_228), .C(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_197), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_197), .A2(n_522), .B(n_523), .Y(n_521) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_200), .Y(n_285) );
INVx1_ASAP7_75t_SL g329 ( .A(n_200), .Y(n_329) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_200), .B(n_278), .C(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_247), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g364 ( .A1(n_210), .A2(n_313), .B(n_365), .C(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_212), .B(n_234), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_212), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g381 ( .A(n_212), .Y(n_381) );
AND2x2_ASAP7_75t_L g402 ( .A(n_212), .B(n_249), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_212), .B(n_311), .Y(n_430) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AND2x2_ASAP7_75t_L g275 ( .A(n_213), .B(n_266), .Y(n_275) );
INVx2_ASAP7_75t_L g282 ( .A(n_213), .Y(n_282) );
AND2x2_ASAP7_75t_L g302 ( .A(n_213), .B(n_249), .Y(n_302) );
AND2x2_ASAP7_75t_L g352 ( .A(n_213), .B(n_234), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_213), .Y(n_356) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_221), .Y(n_533) );
INVx2_ASAP7_75t_SL g266 ( .A(n_223), .Y(n_266) );
BUFx2_ASAP7_75t_L g292 ( .A(n_223), .Y(n_292) );
AND2x2_ASAP7_75t_L g419 ( .A(n_223), .B(n_234), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
INVx1_ASAP7_75t_L g265 ( .A(n_233), .Y(n_265) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_233), .A2(n_528), .B(n_535), .Y(n_527) );
INVx3_ASAP7_75t_SL g249 ( .A(n_234), .Y(n_249) );
AND2x2_ASAP7_75t_L g274 ( .A(n_234), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g281 ( .A(n_234), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g311 ( .A(n_234), .B(n_271), .Y(n_311) );
OR2x2_ASAP7_75t_L g320 ( .A(n_234), .B(n_266), .Y(n_320) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_234), .Y(n_338) );
AND2x2_ASAP7_75t_L g343 ( .A(n_234), .B(n_296), .Y(n_343) );
AND2x2_ASAP7_75t_L g371 ( .A(n_234), .B(n_251), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_234), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g409 ( .A(n_234), .B(n_250), .Y(n_409) );
OR2x6_ASAP7_75t_L g234 ( .A(n_235), .B(n_245), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_241), .C(n_242), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_240), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_243), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x2_ASAP7_75t_L g333 ( .A(n_249), .B(n_282), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_249), .B(n_275), .Y(n_361) );
AND2x2_ASAP7_75t_L g379 ( .A(n_249), .B(n_296), .Y(n_379) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_266), .Y(n_250) );
AND2x2_ASAP7_75t_L g280 ( .A(n_251), .B(n_266), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_251), .B(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g318 ( .A(n_251), .Y(n_318) );
OR2x2_ASAP7_75t_L g366 ( .A(n_251), .B(n_286), .Y(n_366) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_256), .B(n_264), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_253), .A2(n_272), .B(n_273), .Y(n_271) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_253), .A2(n_518), .B(n_524), .Y(n_517) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_254), .A2(n_510), .B(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_255), .A2(n_458), .B(n_465), .Y(n_457) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_255), .A2(n_493), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_255), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g272 ( .A(n_256), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_264), .Y(n_273) );
AND2x2_ASAP7_75t_L g301 ( .A(n_266), .B(n_271), .Y(n_301) );
INVx1_ASAP7_75t_L g309 ( .A(n_266), .Y(n_309) );
AND2x2_ASAP7_75t_L g404 ( .A(n_266), .B(n_282), .Y(n_404) );
AOI222xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_276), .B1(n_279), .B2(n_283), .C1(n_287), .C2(n_290), .Y(n_267) );
INVx1_ASAP7_75t_L g399 ( .A(n_268), .Y(n_399) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_274), .Y(n_268) );
AND2x2_ASAP7_75t_L g295 ( .A(n_269), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g306 ( .A(n_269), .B(n_275), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_269), .B(n_297), .Y(n_322) );
OAI222xp33_ASAP7_75t_L g344 ( .A1(n_269), .A2(n_345), .B1(n_350), .B2(n_351), .C1(n_359), .C2(n_361), .Y(n_344) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g332 ( .A(n_271), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_271), .B(n_352), .Y(n_392) );
AND2x2_ASAP7_75t_L g403 ( .A(n_271), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g411 ( .A(n_274), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_276), .B(n_327), .Y(n_390) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_278), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g348 ( .A(n_278), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx3_ASAP7_75t_L g293 ( .A(n_281), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g383 ( .A1(n_281), .A2(n_384), .B(n_387), .C(n_389), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_281), .B(n_318), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_281), .B(n_301), .Y(n_423) );
AND2x2_ASAP7_75t_L g296 ( .A(n_282), .B(n_292), .Y(n_296) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g323 ( .A(n_285), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_286), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g375 ( .A(n_286), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g414 ( .A(n_286), .B(n_314), .Y(n_414) );
INVx1_ASAP7_75t_L g426 ( .A(n_286), .Y(n_426) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_289), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g407 ( .A(n_292), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_299), .C(n_303), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_295), .A2(n_325), .B1(n_340), .B2(n_343), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_296), .B(n_310), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_296), .B(n_318), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_297), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g360 ( .A(n_297), .Y(n_360) );
AND2x2_ASAP7_75t_L g367 ( .A(n_297), .B(n_347), .Y(n_367) );
INVx2_ASAP7_75t_L g328 ( .A(n_298), .Y(n_328) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NOR4xp25_ASAP7_75t_L g305 ( .A(n_302), .B(n_306), .C(n_307), .D(n_310), .Y(n_305) );
INVx1_ASAP7_75t_SL g376 ( .A(n_303), .Y(n_376) );
AND2x2_ASAP7_75t_L g420 ( .A(n_303), .B(n_421), .Y(n_420) );
OAI211xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_312), .B(n_315), .C(n_324), .Y(n_304) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_311), .B(n_381), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_313), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_431) );
INVx1_ASAP7_75t_SL g386 ( .A(n_314), .Y(n_386) );
AND2x2_ASAP7_75t_L g425 ( .A(n_314), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_318), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_322), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_323), .B(n_348), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_330), .B(n_332), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g400 ( .A(n_327), .Y(n_400) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g428 ( .A(n_328), .Y(n_428) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
OAI21xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B(n_339), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g347 ( .A(n_335), .Y(n_347) );
OR2x2_ASAP7_75t_L g385 ( .A(n_335), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI21xp33_ASAP7_75t_SL g380 ( .A1(n_338), .A2(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_369), .B1(n_372), .B2(n_379), .C(n_380), .Y(n_368) );
INVx1_ASAP7_75t_SL g412 ( .A(n_343), .Y(n_412) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
OR2x2_ASAP7_75t_L g359 ( .A(n_347), .B(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_356), .B2(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g391 ( .A(n_352), .Y(n_391) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_355), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_397), .C(n_410), .D(n_422), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g363 ( .A(n_364), .B(n_368), .C(n_383), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_366), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_373), .B(n_378), .Y(n_382) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_385), .A2(n_411), .B1(n_412), .B2(n_413), .C(n_415), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_387), .A2(n_402), .B(n_403), .C(n_405), .Y(n_401) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_388), .A2(n_406), .B1(n_408), .B2(n_409), .Y(n_405) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_400), .C(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g416 ( .A(n_409), .Y(n_416) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI221xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .B1(n_427), .B2(n_429), .C(n_431), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_437), .A2(n_451), .B1(n_719), .B2(n_720), .Y(n_450) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g447 ( .A(n_442), .Y(n_447) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI21xp33_ASAP7_75t_SL g448 ( .A1(n_446), .A2(n_449), .B(n_735), .Y(n_448) );
INVx1_ASAP7_75t_L g728 ( .A(n_451), .Y(n_728) );
NAND2x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_635), .Y(n_451) );
NOR5xp2_ASAP7_75t_L g452 ( .A(n_453), .B(n_558), .C(n_590), .D(n_605), .E(n_622), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_486), .B(n_505), .C(n_546), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_467), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_455), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_455), .B(n_610), .Y(n_673) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_456), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_456), .B(n_502), .Y(n_559) );
AND2x2_ASAP7_75t_L g600 ( .A(n_456), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_456), .B(n_569), .Y(n_604) );
OR2x2_ASAP7_75t_L g641 ( .A(n_456), .B(n_492), .Y(n_641) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g491 ( .A(n_457), .B(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
OR2x2_ASAP7_75t_L g712 ( .A(n_457), .B(n_552), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_467), .A2(n_615), .B1(n_616), .B2(n_619), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_467), .B(n_549), .Y(n_698) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
AND2x2_ASAP7_75t_L g504 ( .A(n_468), .B(n_492), .Y(n_504) );
AND2x2_ASAP7_75t_L g551 ( .A(n_468), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g556 ( .A(n_468), .Y(n_556) );
INVx3_ASAP7_75t_L g569 ( .A(n_468), .Y(n_569) );
OR2x2_ASAP7_75t_L g589 ( .A(n_468), .B(n_552), .Y(n_589) );
AND2x2_ASAP7_75t_L g608 ( .A(n_468), .B(n_478), .Y(n_608) );
BUFx2_ASAP7_75t_L g640 ( .A(n_468), .Y(n_640) );
AND2x4_ASAP7_75t_L g555 ( .A(n_477), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g490 ( .A(n_478), .Y(n_490) );
INVx2_ASAP7_75t_L g503 ( .A(n_478), .Y(n_503) );
OR2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_552), .Y(n_571) );
AND2x2_ASAP7_75t_L g601 ( .A(n_478), .B(n_492), .Y(n_601) );
AND2x2_ASAP7_75t_L g618 ( .A(n_478), .B(n_549), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_478), .B(n_569), .Y(n_658) );
AND2x2_ASAP7_75t_SL g694 ( .A(n_478), .B(n_504), .Y(n_694) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp33_ASAP7_75t_SL g487 ( .A(n_488), .B(n_501), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_489), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_490), .A2(n_504), .B(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_490), .B(n_492), .Y(n_688) );
AND2x2_ASAP7_75t_L g624 ( .A(n_491), .B(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_492), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_501), .B(n_549), .Y(n_717) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_502), .A2(n_660), .B1(n_661), .B2(n_666), .Y(n_659) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_L g550 ( .A(n_503), .B(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g588 ( .A(n_503), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g625 ( .A(n_503), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_504), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g679 ( .A(n_504), .Y(n_679) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_526), .Y(n_506) );
INVx4_ASAP7_75t_L g565 ( .A(n_507), .Y(n_565) );
AND2x2_ASAP7_75t_L g643 ( .A(n_507), .B(n_610), .Y(n_643) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
INVx3_ASAP7_75t_L g562 ( .A(n_508), .Y(n_562) );
AND2x2_ASAP7_75t_L g576 ( .A(n_508), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
INVx2_ASAP7_75t_L g594 ( .A(n_508), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_508), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g651 ( .A(n_508), .B(n_646), .Y(n_651) );
AND2x2_ASAP7_75t_L g716 ( .A(n_508), .B(n_686), .Y(n_716) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
AND2x2_ASAP7_75t_L g557 ( .A(n_517), .B(n_538), .Y(n_557) );
INVx2_ASAP7_75t_L g577 ( .A(n_517), .Y(n_577) );
INVx1_ASAP7_75t_L g582 ( .A(n_526), .Y(n_582) );
AND2x2_ASAP7_75t_L g628 ( .A(n_526), .B(n_576), .Y(n_628) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
INVx2_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
INVx1_ASAP7_75t_L g575 ( .A(n_527), .Y(n_575) );
AND2x2_ASAP7_75t_L g593 ( .A(n_527), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_527), .B(n_577), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_534), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g610 ( .A(n_537), .B(n_567), .Y(n_610) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g563 ( .A(n_538), .Y(n_563) );
AND2x2_ASAP7_75t_L g646 ( .A(n_538), .B(n_577), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_553), .B(n_557), .Y(n_546) );
INVx1_ASAP7_75t_SL g591 ( .A(n_547), .Y(n_591) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_548), .B(n_555), .Y(n_648) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g597 ( .A(n_549), .B(n_552), .Y(n_597) );
AND2x2_ASAP7_75t_L g626 ( .A(n_549), .B(n_570), .Y(n_626) );
OR2x2_ASAP7_75t_L g629 ( .A(n_549), .B(n_589), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g693 ( .A1(n_550), .A2(n_642), .B1(n_694), .B2(n_695), .C1(n_697), .C2(n_699), .Y(n_693) );
BUFx2_ASAP7_75t_L g607 ( .A(n_552), .Y(n_607) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g596 ( .A(n_555), .B(n_597), .Y(n_596) );
INVx3_ASAP7_75t_SL g613 ( .A(n_555), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_555), .B(n_607), .Y(n_667) );
AND2x2_ASAP7_75t_L g602 ( .A(n_557), .B(n_562), .Y(n_602) );
INVx1_ASAP7_75t_L g621 ( .A(n_557), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_560), .B1(n_564), .B2(n_568), .C(n_572), .Y(n_558) );
OR2x2_ASAP7_75t_L g630 ( .A(n_560), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g615 ( .A(n_562), .B(n_585), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_562), .B(n_575), .Y(n_655) );
AND2x2_ASAP7_75t_L g660 ( .A(n_562), .B(n_610), .Y(n_660) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_562), .Y(n_670) );
NAND2x1_ASAP7_75t_SL g681 ( .A(n_562), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g566 ( .A(n_563), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g586 ( .A(n_563), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_563), .B(n_581), .Y(n_612) );
INVx1_ASAP7_75t_L g678 ( .A(n_563), .Y(n_678) );
INVx1_ASAP7_75t_L g653 ( .A(n_564), .Y(n_653) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g665 ( .A(n_565), .Y(n_665) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_565), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g682 ( .A(n_566), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_566), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g585 ( .A(n_567), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_567), .B(n_577), .Y(n_598) );
INVx1_ASAP7_75t_L g664 ( .A(n_567), .Y(n_664) );
INVx1_ASAP7_75t_L g685 ( .A(n_568), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_578), .B(n_587), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
AND2x2_ASAP7_75t_L g718 ( .A(n_574), .B(n_651), .Y(n_718) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g686 ( .A(n_575), .B(n_646), .Y(n_686) );
AOI32xp33_ASAP7_75t_L g599 ( .A1(n_576), .A2(n_582), .A3(n_600), .B1(n_602), .B2(n_603), .Y(n_599) );
AOI322xp5_ASAP7_75t_L g701 ( .A1(n_576), .A2(n_608), .A3(n_691), .B1(n_702), .B2(n_703), .C1(n_704), .C2(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g581 ( .A(n_577), .Y(n_581) );
INVx1_ASAP7_75t_L g691 ( .A(n_577), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B1(n_583), .B2(n_584), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_579), .B(n_585), .Y(n_634) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_580), .B(n_646), .Y(n_696) );
INVx1_ASAP7_75t_L g583 ( .A(n_581), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_581), .B(n_610), .Y(n_700) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_589), .B(n_684), .Y(n_683) );
OAI221xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_592), .B1(n_595), .B2(n_598), .C(n_599), .Y(n_590) );
OR2x2_ASAP7_75t_L g611 ( .A(n_592), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g620 ( .A(n_592), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g645 ( .A(n_593), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g649 ( .A(n_603), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B1(n_611), .B2(n_613), .C(n_614), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_607), .A2(n_638), .B1(n_642), .B2(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_608), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_608), .Y(n_713) );
INVx1_ASAP7_75t_L g707 ( .A(n_610), .Y(n_707) );
INVx1_ASAP7_75t_SL g642 ( .A(n_611), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_613), .B(n_641), .Y(n_703) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_618), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g684 ( .A(n_618), .Y(n_684) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_627), .B1(n_629), .B2(n_630), .C(n_632), .Y(n_622) );
NOR2xp33_ASAP7_75t_SL g623 ( .A(n_624), .B(n_626), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_624), .A2(n_642), .B1(n_688), .B2(n_689), .Y(n_687) );
CKINVDCx14_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_629), .A2(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR3xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_668), .C(n_692), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_637), .B(n_644), .C(n_652), .D(n_659), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g715 ( .A(n_640), .Y(n_715) );
INVx3_ASAP7_75t_SL g709 ( .A(n_641), .Y(n_709) );
OR2x2_ASAP7_75t_L g714 ( .A(n_641), .B(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_651), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_646), .B(n_664), .Y(n_705) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_656), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_671), .B(n_674), .C(n_687), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g702 ( .A(n_673), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B1(n_680), .B2(n_683), .C1(n_685), .C2(n_686), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND4xp25_ASAP7_75t_SL g711 ( .A(n_684), .B(n_712), .C(n_713), .D(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_701), .C(n_710), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_710) );
INVx1_ASAP7_75t_L g730 ( .A(n_720), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_721), .Y(n_731) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
endmodule