module fake_jpeg_17417_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_20),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_27),
.B1(n_30),
.B2(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_18),
.B1(n_22),
.B2(n_33),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_27),
.B1(n_16),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_80),
.Y(n_100)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_27),
.B1(n_30),
.B2(n_18),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_67),
.B1(n_82),
.B2(n_83),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_75),
.B1(n_79),
.B2(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_43),
.B1(n_44),
.B2(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_86),
.B1(n_88),
.B2(n_0),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_78),
.A2(n_13),
.B(n_15),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_91),
.B1(n_53),
.B2(n_29),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_43),
.B1(n_25),
.B2(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_32),
.A3(n_20),
.B1(n_19),
.B2(n_39),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_93),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_107),
.B1(n_113),
.B2(n_115),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_37),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_112),
.B(n_114),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_104),
.Y(n_139)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_54),
.B1(n_51),
.B2(n_62),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_51),
.B1(n_53),
.B2(n_19),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_19),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_116),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_29),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_35),
.C(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_138),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_107),
.B1(n_114),
.B2(n_97),
.Y(n_151)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_67),
.B1(n_73),
.B2(n_71),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_130),
.B1(n_113),
.B2(n_102),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_73),
.B1(n_84),
.B2(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_84),
.B1(n_68),
.B2(n_70),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_141),
.B1(n_110),
.B2(n_102),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_35),
.C(n_37),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_100),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_87),
.B1(n_85),
.B2(n_35),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_85),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_147),
.B(n_168),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_105),
.B(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_148),
.A2(n_157),
.B(n_170),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_171),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_154),
.B1(n_165),
.B2(n_137),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_95),
.B1(n_101),
.B2(n_97),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_156),
.B1(n_163),
.B2(n_127),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_101),
.B1(n_120),
.B2(n_121),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_121),
.B(n_20),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_109),
.C(n_19),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_138),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_120),
.B1(n_108),
.B2(n_12),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_124),
.A2(n_108),
.B1(n_89),
.B2(n_57),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_125),
.B(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_19),
.B1(n_108),
.B2(n_29),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_122),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_145),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_187),
.C(n_190),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_202),
.B1(n_171),
.B2(n_173),
.Y(n_204)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_189),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_164),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_142),
.C(n_137),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_150),
.B1(n_156),
.B2(n_154),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_142),
.B(n_135),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_193),
.A2(n_159),
.B(n_170),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_141),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_195),
.C(n_196),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_129),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_136),
.C(n_134),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_122),
.B1(n_1),
.B2(n_2),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_119),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_163),
.A2(n_31),
.B1(n_29),
.B2(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_29),
.B1(n_31),
.B2(n_8),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_164),
.B1(n_159),
.B2(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_196),
.B1(n_183),
.B2(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_209),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_160),
.C(n_31),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_226),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_193),
.B(n_177),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_223),
.A2(n_225),
.B(n_201),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_8),
.B(n_15),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_190),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_239),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_194),
.B1(n_187),
.B2(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_198),
.C(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_10),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_246),
.B1(n_225),
.B2(n_206),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_10),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_219),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_251),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_214),
.C(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_258),
.C(n_243),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_214),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_259),
.C(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_215),
.B1(n_204),
.B2(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_223),
.C(n_220),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_216),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_213),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_211),
.B1(n_213),
.B2(n_212),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_262),
.A2(n_233),
.B1(n_238),
.B2(n_247),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_224),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_236),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_241),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_240),
.B1(n_264),
.B2(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_228),
.B1(n_11),
.B2(n_7),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_227),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_248),
.B1(n_235),
.B2(n_230),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_248),
.B1(n_228),
.B2(n_12),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_251),
.C(n_252),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_270),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_286),
.B1(n_14),
.B2(n_5),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_290),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_266),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_256),
.B1(n_259),
.B2(n_250),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_277),
.B(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_273),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_4),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_299),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_268),
.C(n_274),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_300),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_7),
.CI(n_11),
.CON(n_299),
.SN(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_31),
.C(n_5),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_11),
.B1(n_14),
.B2(n_6),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_303),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_14),
.CI(n_5),
.CON(n_302),
.SN(n_302)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_287),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_303),
.B(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_302),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_297),
.B(n_302),
.C(n_296),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_286),
.B1(n_281),
.B2(n_6),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_312),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_305),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_316),
.C(n_311),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_315),
.B(n_308),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_298),
.B(n_300),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_307),
.C(n_314),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_299),
.B(n_4),
.C(n_31),
.Y(n_324)
);


endmodule