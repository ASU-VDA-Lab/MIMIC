module fake_jpeg_6401_n_126 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_28),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_26),
.B1(n_15),
.B2(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_11),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_46),
.B1(n_49),
.B2(n_59),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_50),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_27),
.B1(n_29),
.B2(n_35),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_26),
.B(n_15),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_3),
.B(n_4),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_61),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_39),
.B1(n_21),
.B2(n_17),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_21),
.B1(n_18),
.B2(n_16),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_44),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_19),
.C(n_39),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_77),
.C(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_45),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_78),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_45),
.B1(n_41),
.B2(n_52),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_42),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_9),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_66),
.B1(n_78),
.B2(n_75),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_88),
.Y(n_99)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_92),
.C(n_76),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_44),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_77),
.C(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_61),
.B1(n_54),
.B2(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_67),
.B1(n_70),
.B2(n_74),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_43),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_62),
.B1(n_68),
.B2(n_64),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_94),
.B1(n_48),
.B2(n_43),
.Y(n_109)
);

OAI21x1_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_72),
.B(n_65),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_82),
.B(n_89),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_81),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_88),
.B(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_78),
.B1(n_48),
.B2(n_10),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_80),
.C(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_94),
.B(n_80),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_107),
.C(n_109),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_90),
.B(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_113),
.B(n_110),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_48),
.B(n_6),
.Y(n_123)
);

OAI33xp33_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_123),
.A3(n_121),
.B1(n_7),
.B2(n_6),
.B3(n_5),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_7),
.Y(n_126)
);


endmodule