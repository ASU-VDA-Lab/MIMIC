module fake_jpeg_17196_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_34),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_24),
.B1(n_22),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_60),
.B1(n_64),
.B2(n_47),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_59),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_45),
.B1(n_22),
.B2(n_41),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_59),
.B1(n_53),
.B2(n_51),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_34),
.B1(n_18),
.B2(n_26),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_1),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_68),
.B1(n_31),
.B2(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_27),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_13),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_62),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_69),
.B(n_96),
.C(n_50),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_71),
.B1(n_80),
.B2(n_81),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_38),
.B1(n_35),
.B2(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_49),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_98),
.C(n_100),
.Y(n_117)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_76),
.A2(n_84),
.B1(n_94),
.B2(n_15),
.Y(n_125)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_30),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_97),
.B1(n_10),
.B2(n_11),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_35),
.B1(n_32),
.B2(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_25),
.B1(n_21),
.B2(n_31),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_25),
.B1(n_30),
.B2(n_5),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_86),
.B1(n_101),
.B2(n_11),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_87),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_29),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_17),
.B1(n_28),
.B2(n_40),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_48),
.B1(n_67),
.B2(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_17),
.B1(n_29),
.B2(n_6),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_29),
.B1(n_3),
.B2(n_6),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_43),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_2),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_29),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_121),
.Y(n_129)
);

NOR2x1_ASAP7_75t_SL g104 ( 
.A(n_69),
.B(n_79),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_110),
.B(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_43),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_43),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_125),
.B1(n_76),
.B2(n_97),
.Y(n_151)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_115),
.Y(n_132)
);

XNOR2x2_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_40),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_91),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_74),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_80),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_126),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_40),
.B1(n_43),
.B2(n_50),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_40),
.B1(n_15),
.B2(n_16),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_71),
.Y(n_150)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_16),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_82),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_146),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_75),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_140),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_150),
.B(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_130),
.B1(n_151),
.B2(n_152),
.C(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_102),
.B1(n_103),
.B2(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_174),
.B1(n_129),
.B2(n_150),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_119),
.C(n_96),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_164),
.C(n_165),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_111),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_109),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_96),
.C(n_121),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_175),
.C(n_97),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_121),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_129),
.B(n_130),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_77),
.B1(n_89),
.B2(n_72),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_107),
.C(n_87),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_186),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_192),
.C(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_185),
.B1(n_189),
.B2(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_156),
.B(n_134),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_129),
.B(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_145),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_190),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_138),
.B(n_128),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_168),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_92),
.B1(n_171),
.B2(n_158),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_171),
.B1(n_169),
.B2(n_166),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_196),
.A2(n_204),
.B1(n_189),
.B2(n_185),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_179),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_157),
.B1(n_175),
.B2(n_160),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_157),
.C(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_192),
.Y(n_216)
);

AOI321xp33_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_155),
.A3(n_162),
.B1(n_174),
.B2(n_167),
.C(n_172),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_216),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_181),
.B1(n_195),
.B2(n_182),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_221),
.B(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_227),
.Y(n_235)
);

OAI221xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_220),
.B1(n_208),
.B2(n_213),
.C(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_197),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_231),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_213),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_200),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_217),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_239),
.B(n_240),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_178),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_243),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_223),
.CI(n_205),
.CON(n_243),
.SN(n_243)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_238),
.B(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_222),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_245),
.B(n_237),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_92),
.Y(n_248)
);


endmodule