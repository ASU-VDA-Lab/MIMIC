module fake_netlist_1_206_n_1350 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1350);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1350;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g309 ( .A(n_117), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_27), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_24), .Y(n_311) );
CKINVDCx14_ASAP7_75t_R g312 ( .A(n_223), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_274), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_123), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_232), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_265), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_98), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_199), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_58), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g320 ( .A(n_36), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_78), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_273), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_99), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_139), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_150), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_137), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_266), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_221), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_67), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_28), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_165), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_8), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_56), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_172), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_24), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_185), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_282), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_209), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_261), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_181), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_156), .Y(n_341) );
INVxp67_ASAP7_75t_SL g342 ( .A(n_7), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_241), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_196), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_254), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_45), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_82), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_127), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_125), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
BUFx2_ASAP7_75t_SL g352 ( .A(n_49), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_205), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_89), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_16), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_291), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_234), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_250), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_300), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_54), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_30), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_40), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_296), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_9), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_27), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_37), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_192), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_279), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_286), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_50), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_162), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_141), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_42), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_288), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_245), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_171), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_216), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_145), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_242), .Y(n_379) );
BUFx8_ASAP7_75t_SL g380 ( .A(n_174), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_36), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_270), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_236), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_230), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_260), .B(n_175), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_132), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_244), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_7), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_202), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_0), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_61), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_9), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_75), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_62), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_103), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_298), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_68), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_59), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_146), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_1), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_289), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_276), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_91), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_64), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_106), .Y(n_405) );
INVxp33_ASAP7_75t_L g406 ( .A(n_136), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_271), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_210), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_214), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_39), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_114), .Y(n_411) );
INVxp33_ASAP7_75t_L g412 ( .A(n_157), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_81), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g414 ( .A(n_5), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_255), .Y(n_415) );
BUFx10_ASAP7_75t_L g416 ( .A(n_297), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_112), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_240), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_88), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_59), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_243), .Y(n_421) );
CKINVDCx16_ASAP7_75t_R g422 ( .A(n_249), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_187), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_97), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_224), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_107), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_10), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_195), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_219), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_239), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_268), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_49), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_15), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_170), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_182), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_306), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_84), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_90), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_67), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_108), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_278), .Y(n_441) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_218), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_168), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_262), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_280), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_54), .Y(n_446) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_68), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_301), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_188), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_211), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_251), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_63), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_30), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_152), .B(n_124), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_159), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_48), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_61), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_20), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_126), .Y(n_459) );
INVxp33_ASAP7_75t_SL g460 ( .A(n_304), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_269), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_259), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_277), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_197), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_143), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_120), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_155), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_184), .B(n_6), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_267), .Y(n_469) );
BUFx10_ASAP7_75t_L g470 ( .A(n_290), .Y(n_470) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_130), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_311), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_431), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_311), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_380), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_431), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_419), .B(n_0), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_410), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_341), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_410), .Y(n_480) );
INVx5_ASAP7_75t_L g481 ( .A(n_448), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_375), .B(n_1), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_448), .Y(n_483) );
AND2x2_ASAP7_75t_SL g484 ( .A(n_408), .B(n_385), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_448), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_432), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_448), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_419), .B(n_2), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_341), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_432), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_446), .B(n_2), .Y(n_491) );
NOR2xp33_ASAP7_75t_SL g492 ( .A(n_389), .B(n_96), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_344), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_344), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_320), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_406), .B(n_3), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_349), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_452), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_453), .B(n_4), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_382), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_349), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_380), .Y(n_502) );
OAI22x1_ASAP7_75t_SL g503 ( .A1(n_393), .A2(n_10), .B1(n_6), .B2(n_8), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_425), .B(n_11), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_374), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_382), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_406), .B(n_11), .Y(n_507) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_374), .A2(n_101), .B(n_100), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_386), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_377), .B(n_12), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_436), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_436), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_479), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_496), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_496), .B(n_329), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_487), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_487), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_484), .B(n_412), .Y(n_519) );
NOR2x1p5_ASAP7_75t_L g520 ( .A(n_475), .B(n_319), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_484), .B(n_407), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_487), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_507), .B(n_412), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_493), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_487), .Y(n_525) );
BUFx10_ASAP7_75t_L g526 ( .A(n_484), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_507), .B(n_422), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_493), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_479), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_492), .B(n_477), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_487), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_487), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_489), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_479), .B(n_411), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
NAND2xp33_ASAP7_75t_L g539 ( .A(n_489), .B(n_313), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_511), .B(n_414), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_489), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_508), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_489), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_509), .B(n_319), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_494), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_509), .B(n_473), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_473), .B(n_353), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_489), .Y(n_548) );
XOR2xp5_ASAP7_75t_L g549 ( .A(n_503), .B(n_393), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_502), .B(n_456), .Y(n_550) );
CKINVDCx11_ASAP7_75t_R g551 ( .A(n_495), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_509), .B(n_321), .Y(n_552) );
OR2x6_ASAP7_75t_L g553 ( .A(n_495), .B(n_352), .Y(n_553) );
INVx4_ASAP7_75t_L g554 ( .A(n_477), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_503), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_477), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_508), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_488), .B(n_312), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_494), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_553), .A2(n_343), .B1(n_426), .B2(n_334), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_523), .B(n_488), .Y(n_562) );
NAND2x1_ASAP7_75t_L g563 ( .A(n_554), .B(n_488), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_523), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_551), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_515), .B(n_488), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_530), .B(n_476), .Y(n_567) );
BUFx3_ASAP7_75t_L g568 ( .A(n_524), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_542), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_520), .B(n_499), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_540), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g572 ( .A(n_540), .B(n_516), .Y(n_572) );
BUFx5_ASAP7_75t_L g573 ( .A(n_514), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_516), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_527), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_550), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_536), .B(n_482), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_550), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g580 ( .A1(n_519), .A2(n_499), .B(n_491), .C(n_420), .Y(n_580) );
INVx4_ASAP7_75t_L g581 ( .A(n_554), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_554), .A2(n_504), .B1(n_460), .B2(n_476), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_559), .B(n_322), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_514), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_530), .B(n_476), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_530), .B(n_460), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_554), .A2(n_312), .B1(n_471), .B2(n_335), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_524), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_528), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_526), .B(n_321), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_521), .A2(n_343), .B1(n_426), .B2(n_334), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_544), .B(n_322), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_556), .B(n_337), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_552), .B(n_337), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_547), .B(n_339), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_531), .A2(n_501), .B(n_497), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_553), .A2(n_437), .B1(n_466), .B2(n_361), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_528), .B(n_339), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_529), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_520), .B(n_466), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_526), .B(n_461), .Y(n_602) );
AND2x6_ASAP7_75t_SL g603 ( .A(n_553), .B(n_333), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_526), .A2(n_361), .B1(n_310), .B2(n_332), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_553), .B(n_354), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_534), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
INVx5_ASAP7_75t_L g608 ( .A(n_542), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_538), .B(n_443), .Y(n_609) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_545), .B(n_497), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_560), .B(n_443), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_560), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g613 ( .A(n_555), .B(n_501), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_546), .B(n_444), .Y(n_614) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_542), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_542), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_542), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_553), .B(n_403), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_542), .A2(n_362), .B1(n_370), .B2(n_330), .Y(n_619) );
AND2x6_ASAP7_75t_SL g620 ( .A(n_549), .B(n_347), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_549), .B(n_381), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_557), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_557), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_557), .B(n_449), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_557), .B(n_400), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_557), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_539), .B(n_449), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_535), .A2(n_437), .B1(n_458), .B2(n_427), .Y(n_628) );
O2A1O1Ixp5_ASAP7_75t_L g629 ( .A1(n_541), .A2(n_434), .B(n_442), .C(n_338), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_537), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_541), .A2(n_471), .B1(n_348), .B2(n_364), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_543), .B(n_463), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_537), .B(n_342), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_548), .A2(n_360), .B1(n_366), .B2(n_365), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_543), .B(n_463), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_548), .A2(n_512), .B(n_505), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_558), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_558), .B(n_512), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_558), .B(n_512), .Y(n_639) );
NAND2x1_ASAP7_75t_L g640 ( .A(n_517), .B(n_513), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_522), .B(n_416), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_517), .B(n_513), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_517), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_518), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_571), .B(n_373), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_575), .B(n_447), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_564), .A2(n_390), .B(n_391), .C(n_388), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_616), .A2(n_445), .B(n_314), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_572), .B(n_394), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_574), .A2(n_398), .B(n_404), .C(n_397), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_626), .A2(n_317), .B(n_309), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_622), .A2(n_323), .B(n_318), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_562), .A2(n_438), .B(n_457), .C(n_433), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_566), .B(n_472), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_591), .A2(n_392), .B1(n_413), .B2(n_355), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_576), .B(n_472), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_561), .B(n_478), .C(n_474), .Y(n_657) );
INVx4_ASAP7_75t_L g658 ( .A(n_581), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_581), .B(n_315), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_580), .A2(n_513), .B(n_478), .C(n_480), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_563), .A2(n_326), .B(n_325), .Y(n_661) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_568), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_567), .A2(n_328), .B(n_327), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_567), .A2(n_340), .B(n_336), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_579), .B(n_486), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_590), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_597), .A2(n_468), .B(n_490), .C(n_486), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_605), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_570), .B(n_490), .Y(n_669) );
OR2x6_ASAP7_75t_L g670 ( .A(n_601), .B(n_498), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_585), .A2(n_346), .B(n_345), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_585), .A2(n_351), .B(n_350), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_586), .A2(n_358), .B(n_357), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_570), .B(n_498), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_633), .Y(n_675) );
INVx4_ASAP7_75t_L g676 ( .A(n_603), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_604), .B(n_416), .Y(n_677) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_598), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_586), .A2(n_363), .B(n_359), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_624), .A2(n_368), .B(n_367), .Y(n_680) );
BUFx8_ASAP7_75t_L g681 ( .A(n_618), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_595), .A2(n_372), .B(n_369), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_613), .B(n_510), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_606), .Y(n_684) );
BUFx8_ASAP7_75t_L g685 ( .A(n_621), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_599), .A2(n_510), .B1(n_454), .B2(n_392), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_599), .B(n_316), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_625), .A2(n_392), .B1(n_413), .B2(n_355), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_595), .A2(n_378), .B(n_376), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_609), .B(n_470), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_SL g691 ( .A1(n_642), .A2(n_395), .B(n_399), .C(n_387), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_609), .B(n_611), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_611), .A2(n_402), .B(n_401), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_592), .A2(n_392), .B1(n_413), .B2(n_355), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_614), .B(n_324), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_569), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_608), .A2(n_409), .B(n_405), .Y(n_697) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_578), .A2(n_356), .B(n_331), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_614), .B(n_371), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_594), .B(n_470), .Y(n_700) );
BUFx12f_ASAP7_75t_L g701 ( .A(n_620), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_588), .Y(n_702) );
BUFx3_ASAP7_75t_L g703 ( .A(n_610), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_594), .B(n_470), .Y(n_704) );
OAI21xp33_ASAP7_75t_SL g705 ( .A1(n_589), .A2(n_423), .B(n_421), .Y(n_705) );
AO21x1_ASAP7_75t_L g706 ( .A1(n_636), .A2(n_428), .B(n_424), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_583), .B(n_379), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_582), .A2(n_413), .B1(n_439), .B2(n_355), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_596), .B(n_383), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_587), .A2(n_439), .B1(n_430), .B2(n_435), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_602), .A2(n_439), .B1(n_506), .B2(n_500), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_607), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_628), .B(n_384), .Y(n_713) );
NAND2x2_ASAP7_75t_L g714 ( .A(n_565), .B(n_386), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g715 ( .A(n_623), .B(n_396), .Y(n_715) );
NOR2xp33_ASAP7_75t_SL g716 ( .A(n_573), .B(n_415), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_596), .B(n_417), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_593), .B(n_418), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_577), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_612), .A2(n_439), .B1(n_441), .B2(n_440), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_617), .A2(n_455), .B(n_450), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_619), .B(n_429), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_569), .A2(n_464), .B(n_459), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_634), .Y(n_724) );
O2A1O1Ixp5_ASAP7_75t_L g725 ( .A1(n_635), .A2(n_462), .B(n_465), .C(n_467), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_569), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_634), .B(n_469), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_631), .B(n_13), .Y(n_728) );
AND2x4_ASAP7_75t_L g729 ( .A(n_584), .B(n_451), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_573), .B(n_627), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_615), .A2(n_465), .B(n_462), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_573), .B(n_13), .Y(n_732) );
BUFx8_ASAP7_75t_L g733 ( .A(n_600), .Y(n_733) );
AOI21x1_ASAP7_75t_L g734 ( .A1(n_640), .A2(n_525), .B(n_518), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_632), .A2(n_506), .B1(n_500), .B2(n_483), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g736 ( .A1(n_642), .A2(n_506), .B(n_485), .Y(n_736) );
INVx4_ASAP7_75t_L g737 ( .A(n_615), .Y(n_737) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_615), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_637), .B(n_14), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_638), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_630), .A2(n_532), .B(n_525), .Y(n_741) );
NOR2xp33_ASAP7_75t_SL g742 ( .A(n_639), .B(n_506), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_639), .B(n_14), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_643), .B(n_15), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_644), .B(n_506), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_571), .B(n_16), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_568), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_568), .Y(n_748) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_571), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_571), .A2(n_481), .B1(n_533), .B2(n_19), .Y(n_750) );
OAI22x1_ASAP7_75t_L g751 ( .A1(n_592), .A2(n_19), .B1(n_17), .B2(n_18), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_616), .A2(n_533), .B(n_481), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_571), .B(n_17), .Y(n_753) );
AO32x1_ASAP7_75t_L g754 ( .A1(n_626), .A2(n_522), .A3(n_481), .B1(n_21), .B2(n_22), .Y(n_754) );
O2A1O1Ixp5_ASAP7_75t_SL g755 ( .A1(n_641), .A2(n_522), .B(n_481), .C(n_104), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_568), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_561), .B(n_20), .C(n_21), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_572), .A2(n_481), .B1(n_522), .B2(n_26), .Y(n_758) );
OAI21xp33_ASAP7_75t_L g759 ( .A1(n_571), .A2(n_23), .B(n_25), .Y(n_759) );
OA22x2_ASAP7_75t_L g760 ( .A1(n_561), .A2(n_28), .B1(n_23), .B2(n_25), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_571), .B(n_29), .Y(n_761) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_568), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_571), .B(n_31), .Y(n_763) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_568), .Y(n_764) );
OAI21xp5_ASAP7_75t_L g765 ( .A1(n_629), .A2(n_105), .B(n_102), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_571), .B(n_32), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_568), .Y(n_767) );
INVxp67_ASAP7_75t_SL g768 ( .A(n_561), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g769 ( .A1(n_562), .A2(n_35), .B(n_33), .C(n_34), .Y(n_769) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_572), .B(n_34), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_568), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_724), .A2(n_38), .B1(n_35), .B2(n_37), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_669), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_692), .A2(n_110), .B(n_109), .Y(n_774) );
OR2x6_ASAP7_75t_L g775 ( .A(n_701), .B(n_38), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_749), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_668), .B(n_41), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_733), .Y(n_778) );
AO31x2_ASAP7_75t_L g779 ( .A1(n_706), .A2(n_42), .A3(n_43), .B(n_44), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_730), .A2(n_113), .B(n_111), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_650), .B(n_43), .C(n_44), .Y(n_781) );
AO31x2_ASAP7_75t_L g782 ( .A1(n_667), .A2(n_45), .A3(n_46), .B(n_47), .Y(n_782) );
AO31x2_ASAP7_75t_L g783 ( .A1(n_732), .A2(n_46), .A3(n_47), .B(n_48), .Y(n_783) );
BUFx2_ASAP7_75t_L g784 ( .A(n_733), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_666), .B(n_51), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_768), .B(n_51), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_696), .A2(n_116), .B(n_115), .Y(n_787) );
AO31x2_ASAP7_75t_L g788 ( .A1(n_686), .A2(n_52), .A3(n_53), .B(n_55), .Y(n_788) );
AO21x2_ASAP7_75t_L g789 ( .A1(n_765), .A2(n_119), .B(n_118), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_662), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_740), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_674), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_656), .B(n_52), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_675), .B(n_53), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_753), .B(n_55), .Y(n_795) );
AO21x1_ASAP7_75t_L g796 ( .A1(n_731), .A2(n_122), .B(n_121), .Y(n_796) );
AO31x2_ASAP7_75t_L g797 ( .A1(n_708), .A2(n_769), .A3(n_750), .B(n_710), .Y(n_797) );
NAND2x1p5_ASAP7_75t_L g798 ( .A(n_662), .B(n_56), .Y(n_798) );
O2A1O1Ixp5_ASAP7_75t_SL g799 ( .A1(n_720), .A2(n_194), .B(n_303), .C(n_302), .Y(n_799) );
AOI31xp67_ASAP7_75t_L g800 ( .A1(n_735), .A2(n_191), .A3(n_299), .B(n_295), .Y(n_800) );
BUFx3_ASAP7_75t_L g801 ( .A(n_762), .Y(n_801) );
BUFx2_ASAP7_75t_L g802 ( .A(n_762), .Y(n_802) );
BUFx4f_ASAP7_75t_SL g803 ( .A(n_685), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_678), .B(n_57), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_726), .A2(n_129), .B(n_128), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_752), .A2(n_133), .B(n_131), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_702), .Y(n_807) );
BUFx3_ASAP7_75t_L g808 ( .A(n_762), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_657), .B(n_57), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_665), .B(n_58), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_670), .B(n_677), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_670), .B(n_60), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g813 ( .A1(n_682), .A2(n_135), .B(n_134), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_689), .A2(n_62), .B(n_63), .C(n_64), .Y(n_814) );
INVx5_ASAP7_75t_L g815 ( .A(n_764), .Y(n_815) );
OAI22xp33_ASAP7_75t_L g816 ( .A1(n_760), .A2(n_65), .B1(n_66), .B2(n_69), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_761), .B(n_66), .Y(n_817) );
BUFx4f_ASAP7_75t_L g818 ( .A(n_744), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_712), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_744), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_684), .Y(n_821) );
OAI21x1_ASAP7_75t_L g822 ( .A1(n_741), .A2(n_203), .B(n_294), .Y(n_822) );
INVx2_ASAP7_75t_SL g823 ( .A(n_685), .Y(n_823) );
BUFx12f_ASAP7_75t_L g824 ( .A(n_681), .Y(n_824) );
BUFx2_ASAP7_75t_L g825 ( .A(n_764), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_763), .Y(n_826) );
AO31x2_ASAP7_75t_L g827 ( .A1(n_751), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_654), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_743), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_738), .A2(n_204), .B(n_293), .Y(n_830) );
OR2x6_ASAP7_75t_L g831 ( .A(n_676), .B(n_71), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_693), .A2(n_206), .B(n_292), .Y(n_832) );
AO31x2_ASAP7_75t_L g833 ( .A1(n_737), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_833) );
BUFx3_ASAP7_75t_L g834 ( .A(n_681), .Y(n_834) );
O2A1O1Ixp33_ASAP7_75t_L g835 ( .A1(n_653), .A2(n_72), .B(n_73), .C(n_74), .Y(n_835) );
BUFx2_ASAP7_75t_L g836 ( .A(n_658), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_658), .Y(n_837) );
AO31x2_ASAP7_75t_L g838 ( .A1(n_737), .A2(n_75), .A3(n_76), .B(n_77), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_719), .Y(n_839) );
NAND2xp5_ASAP7_75t_SL g840 ( .A(n_715), .B(n_76), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_746), .B(n_77), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_646), .B(n_78), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_766), .B(n_79), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g844 ( .A1(n_673), .A2(n_212), .B(n_287), .Y(n_844) );
O2A1O1Ixp33_ASAP7_75t_L g845 ( .A1(n_647), .A2(n_80), .B(n_81), .C(n_82), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_649), .B(n_80), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_651), .A2(n_208), .B(n_285), .Y(n_847) );
AOI21xp5_ASAP7_75t_L g848 ( .A1(n_690), .A2(n_207), .B(n_284), .Y(n_848) );
AO31x2_ASAP7_75t_L g849 ( .A1(n_680), .A2(n_83), .A3(n_84), .B(n_85), .Y(n_849) );
AO31x2_ASAP7_75t_L g850 ( .A1(n_679), .A2(n_83), .A3(n_85), .B(n_86), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_688), .B(n_87), .C(n_88), .Y(n_851) );
O2A1O1Ixp33_ASAP7_75t_L g852 ( .A1(n_705), .A2(n_87), .B(n_89), .C(n_90), .Y(n_852) );
A2O1A1Ixp33_ASAP7_75t_L g853 ( .A1(n_660), .A2(n_91), .B(n_92), .C(n_93), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_687), .A2(n_220), .B(n_283), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g855 ( .A(n_716), .B(n_92), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_645), .B(n_93), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_757), .A2(n_94), .B1(n_95), .B2(n_138), .Y(n_857) );
BUFx4f_ASAP7_75t_L g858 ( .A(n_683), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_648), .A2(n_222), .B(n_140), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_683), .B(n_94), .Y(n_860) );
AO31x2_ASAP7_75t_L g861 ( .A1(n_663), .A2(n_142), .A3(n_144), .B(n_147), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_695), .A2(n_148), .B(n_149), .Y(n_862) );
AO31x2_ASAP7_75t_L g863 ( .A1(n_664), .A2(n_151), .A3(n_153), .B(n_154), .Y(n_863) );
AO31x2_ASAP7_75t_L g864 ( .A1(n_671), .A2(n_158), .A3(n_160), .B(n_161), .Y(n_864) );
NAND2xp5_ASAP7_75t_SL g865 ( .A(n_747), .B(n_163), .Y(n_865) );
AO21x1_ASAP7_75t_L g866 ( .A1(n_652), .A2(n_164), .B(n_166), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_700), .B(n_167), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_699), .A2(n_169), .B(n_173), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_704), .A2(n_176), .B(n_177), .Y(n_869) );
AO31x2_ASAP7_75t_L g870 ( .A1(n_672), .A2(n_178), .A3(n_179), .B(n_180), .Y(n_870) );
A2O1A1Ixp33_ASAP7_75t_L g871 ( .A1(n_759), .A2(n_183), .B(n_186), .C(n_189), .Y(n_871) );
INVx5_ASAP7_75t_L g872 ( .A(n_748), .Y(n_872) );
O2A1O1Ixp33_ASAP7_75t_L g873 ( .A1(n_694), .A2(n_190), .B(n_193), .C(n_198), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_661), .A2(n_200), .B(n_201), .C(n_213), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_721), .A2(n_215), .B(n_217), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_723), .A2(n_225), .B(n_226), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_709), .A2(n_227), .B(n_228), .Y(n_877) );
INVxp67_ASAP7_75t_SL g878 ( .A(n_767), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_770), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_756), .B(n_308), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_717), .A2(n_229), .B(n_231), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_728), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_727), .A2(n_233), .B(n_235), .C(n_237), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_718), .A2(n_238), .B(n_246), .Y(n_884) );
O2A1O1Ixp33_ASAP7_75t_SL g885 ( .A1(n_722), .A2(n_247), .B(n_248), .C(n_252), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_707), .A2(n_253), .B(n_256), .Y(n_886) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_725), .A2(n_257), .B(n_258), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_771), .B(n_739), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g889 ( .A1(n_697), .A2(n_263), .B(n_264), .Y(n_889) );
OR2x6_ASAP7_75t_L g890 ( .A(n_659), .B(n_272), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_698), .B(n_275), .Y(n_891) );
CKINVDCx6p67_ASAP7_75t_R g892 ( .A(n_703), .Y(n_892) );
INVx2_ASAP7_75t_SL g893 ( .A(n_714), .Y(n_893) );
OAI21xp5_ASAP7_75t_SL g894 ( .A1(n_713), .A2(n_281), .B(n_758), .Y(n_894) );
BUFx2_ASAP7_75t_L g895 ( .A(n_729), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_691), .Y(n_896) );
BUFx2_ASAP7_75t_L g897 ( .A(n_745), .Y(n_897) );
AO32x2_ASAP7_75t_L g898 ( .A1(n_754), .A2(n_742), .A3(n_736), .B1(n_711), .B2(n_655), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_754), .A2(n_622), .B(n_626), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_754), .A2(n_622), .B(n_626), .Y(n_900) );
NOR2xp33_ASAP7_75t_SL g901 ( .A(n_701), .B(n_561), .Y(n_901) );
OAI21x1_ASAP7_75t_L g902 ( .A1(n_755), .A2(n_616), .B(n_734), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_692), .A2(n_622), .B(n_626), .Y(n_903) );
AOI21xp5_ASAP7_75t_L g904 ( .A1(n_692), .A2(n_622), .B(n_626), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_749), .B(n_571), .Y(n_905) );
INVx4_ASAP7_75t_L g906 ( .A(n_662), .Y(n_906) );
NOR2xp33_ASAP7_75t_SL g907 ( .A(n_701), .B(n_561), .Y(n_907) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_662), .Y(n_908) );
INVx1_ASAP7_75t_SL g909 ( .A(n_749), .Y(n_909) );
AO22x2_ASAP7_75t_L g910 ( .A1(n_768), .A2(n_561), .B1(n_744), .B2(n_678), .Y(n_910) );
AOI21xp5_ASAP7_75t_L g911 ( .A1(n_692), .A2(n_622), .B(n_626), .Y(n_911) );
AND2x4_ASAP7_75t_L g912 ( .A(n_658), .B(n_572), .Y(n_912) );
INVx3_ASAP7_75t_L g913 ( .A(n_733), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_749), .B(n_571), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_899), .A2(n_900), .B(n_902), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_807), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_824), .Y(n_917) );
OR2x2_ASAP7_75t_L g918 ( .A(n_914), .B(n_909), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_903), .A2(n_911), .B(n_829), .Y(n_919) );
INVxp67_ASAP7_75t_L g920 ( .A(n_905), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_828), .B(n_791), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_819), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_821), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_794), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_793), .Y(n_925) );
AO21x2_ASAP7_75t_L g926 ( .A1(n_887), .A2(n_896), .B(n_789), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_784), .Y(n_927) );
OAI21x1_ASAP7_75t_SL g928 ( .A1(n_844), .A2(n_813), .B(n_832), .Y(n_928) );
CKINVDCx14_ASAP7_75t_R g929 ( .A(n_775), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g930 ( .A(n_811), .B(n_826), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_901), .B(n_907), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_882), .B(n_773), .Y(n_932) );
BUFx3_ASAP7_75t_L g933 ( .A(n_913), .Y(n_933) );
NAND2x1p5_ASAP7_75t_L g934 ( .A(n_815), .B(n_906), .Y(n_934) );
OA21x2_ASAP7_75t_L g935 ( .A1(n_822), .A2(n_871), .B(n_806), .Y(n_935) );
INVx3_ASAP7_75t_L g936 ( .A(n_815), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_778), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_804), .A2(n_853), .B(n_809), .Y(n_938) );
BUFx3_ASAP7_75t_L g939 ( .A(n_803), .Y(n_939) );
OAI21x1_ASAP7_75t_L g940 ( .A1(n_799), .A2(n_787), .B(n_805), .Y(n_940) );
AO21x2_ASAP7_75t_L g941 ( .A1(n_866), .A2(n_875), .B(n_889), .Y(n_941) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_846), .A2(n_843), .B(n_841), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_839), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_810), .Y(n_944) );
INVx3_ASAP7_75t_L g945 ( .A(n_801), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_858), .B(n_812), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_792), .B(n_910), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_842), .Y(n_948) );
A2O1A1Ixp33_ASAP7_75t_L g949 ( .A1(n_835), .A2(n_856), .B(n_852), .C(n_845), .Y(n_949) );
OR2x2_ASAP7_75t_L g950 ( .A(n_795), .B(n_834), .Y(n_950) );
BUFx12f_ASAP7_75t_L g951 ( .A(n_775), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_786), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_785), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_860), .Y(n_954) );
OA21x2_ASAP7_75t_L g955 ( .A1(n_796), .A2(n_876), .B(n_774), .Y(n_955) );
OAI21x1_ASAP7_75t_L g956 ( .A1(n_830), .A2(n_881), .B(n_877), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_777), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_788), .Y(n_958) );
OA21x2_ASAP7_75t_L g959 ( .A1(n_886), .A2(n_884), .B(n_874), .Y(n_959) );
OAI21xp5_ASAP7_75t_L g960 ( .A1(n_848), .A2(n_869), .B(n_814), .Y(n_960) );
OAI21x1_ASAP7_75t_L g961 ( .A1(n_780), .A2(n_865), .B(n_862), .Y(n_961) );
AO31x2_ASAP7_75t_L g962 ( .A1(n_883), .A2(n_891), .A3(n_772), .B(n_859), .Y(n_962) );
AND2x4_ASAP7_75t_L g963 ( .A(n_912), .B(n_837), .Y(n_963) );
INVxp67_ASAP7_75t_SL g964 ( .A(n_897), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_912), .B(n_888), .Y(n_965) );
AND2x4_ASAP7_75t_L g966 ( .A(n_836), .B(n_880), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_910), .B(n_820), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_831), .Y(n_968) );
INVx3_ASAP7_75t_L g969 ( .A(n_808), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_868), .A2(n_854), .B(n_847), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_788), .Y(n_971) );
AO21x2_ASAP7_75t_L g972 ( .A1(n_898), .A2(n_816), .B(n_894), .Y(n_972) );
OR2x2_ASAP7_75t_L g973 ( .A(n_823), .B(n_892), .Y(n_973) );
OAI21x1_ASAP7_75t_L g974 ( .A1(n_873), .A2(n_798), .B(n_879), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_831), .B(n_895), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_850), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_797), .B(n_817), .Y(n_977) );
OA21x2_ASAP7_75t_L g978 ( .A1(n_898), .A2(n_857), .B(n_851), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_850), .Y(n_979) );
OAI21x1_ASAP7_75t_L g980 ( .A1(n_855), .A2(n_867), .B(n_908), .Y(n_980) );
OAI21xp5_ASAP7_75t_L g981 ( .A1(n_781), .A2(n_800), .B(n_776), .Y(n_981) );
AO31x2_ASAP7_75t_L g982 ( .A1(n_898), .A2(n_870), .A3(n_864), .B(n_863), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_797), .B(n_878), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_783), .Y(n_984) );
AO21x2_ASAP7_75t_L g985 ( .A1(n_885), .A2(n_840), .B(n_880), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_783), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_890), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_890), .A2(n_872), .B1(n_802), .B2(n_825), .Y(n_988) );
NOR3xp33_ASAP7_75t_L g989 ( .A(n_893), .B(n_827), .C(n_782), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_872), .B(n_783), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_849), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_779), .B(n_782), .Y(n_992) );
OA21x2_ASAP7_75t_L g993 ( .A1(n_861), .A2(n_863), .B(n_782), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_849), .A2(n_827), .B1(n_779), .B2(n_833), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_849), .B(n_833), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_838), .B(n_571), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_838), .Y(n_997) );
BUFx2_ASAP7_75t_R g998 ( .A(n_834), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_807), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_909), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_909), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_905), .B(n_571), .Y(n_1002) );
BUFx8_ASAP7_75t_SL g1003 ( .A(n_824), .Y(n_1003) );
INVx4_ASAP7_75t_SL g1004 ( .A(n_803), .Y(n_1004) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_828), .B(n_791), .Y(n_1005) );
O2A1O1Ixp33_ASAP7_75t_L g1006 ( .A1(n_781), .A2(n_574), .B(n_521), .C(n_845), .Y(n_1006) );
NAND2x1p5_ASAP7_75t_L g1007 ( .A(n_818), .B(n_815), .Y(n_1007) );
AO21x1_ASAP7_75t_L g1008 ( .A1(n_816), .A2(n_896), .B(n_852), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1009 ( .A(n_828), .B(n_791), .Y(n_1009) );
AOI21xp5_ASAP7_75t_L g1010 ( .A1(n_899), .A2(n_900), .B(n_622), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g1011 ( .A(n_790), .Y(n_1011) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_828), .B(n_791), .Y(n_1012) );
NAND2x1p5_ASAP7_75t_L g1013 ( .A(n_818), .B(n_815), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_905), .B(n_571), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_828), .B(n_791), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_914), .B(n_749), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_818), .A2(n_910), .B1(n_744), .B2(n_768), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_818), .A2(n_561), .B1(n_768), .B2(n_901), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_828), .B(n_791), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_807), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_807), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1022 ( .A(n_909), .Y(n_1022) );
AND2x4_ASAP7_75t_L g1023 ( .A(n_828), .B(n_791), .Y(n_1023) );
INVx4_ASAP7_75t_L g1024 ( .A(n_803), .Y(n_1024) );
OAI21xp5_ASAP7_75t_L g1025 ( .A1(n_903), .A2(n_692), .B(n_904), .Y(n_1025) );
BUFx2_ASAP7_75t_R g1026 ( .A(n_834), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_807), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_807), .Y(n_1028) );
AO21x2_ASAP7_75t_L g1029 ( .A1(n_899), .A2(n_900), .B(n_902), .Y(n_1029) );
NOR2xp33_ASAP7_75t_L g1030 ( .A(n_811), .B(n_561), .Y(n_1030) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_1007), .Y(n_1031) );
OR2x6_ASAP7_75t_L g1032 ( .A(n_966), .B(n_987), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_1000), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_916), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_984), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_922), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_999), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_986), .Y(n_1038) );
HB1xp67_ASAP7_75t_L g1039 ( .A(n_1001), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_976), .Y(n_1040) );
CKINVDCx5p33_ASAP7_75t_R g1041 ( .A(n_1003), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_979), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1002), .B(n_1014), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_958), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_1022), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_1005), .B(n_1009), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_947), .B(n_967), .Y(n_1047) );
AO21x1_ASAP7_75t_SL g1048 ( .A1(n_983), .A2(n_988), .B(n_1025), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1016), .B(n_932), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1029), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_1017), .A2(n_1018), .B1(n_1030), .B2(n_1008), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_947), .B(n_967), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1009), .B(n_1012), .Y(n_1053) );
INVx2_ASAP7_75t_L g1054 ( .A(n_915), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_1007), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1020), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1012), .B(n_1023), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_1013), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_918), .Y(n_1059) );
INVxp67_ASAP7_75t_L g1060 ( .A(n_927), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_971), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1021), .Y(n_1062) );
NOR2xp33_ASAP7_75t_SL g1063 ( .A(n_1024), .B(n_998), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_964), .A2(n_1017), .B1(n_1019), .B2(n_1015), .Y(n_1064) );
AO21x2_ASAP7_75t_L g1065 ( .A1(n_1010), .A2(n_928), .B(n_994), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1027), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_921), .B(n_1015), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_921), .B(n_1019), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1028), .Y(n_1069) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_919), .B(n_990), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_943), .B(n_923), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_996), .B(n_932), .Y(n_1072) );
OR2x6_ASAP7_75t_L g1073 ( .A(n_1013), .B(n_934), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_952), .Y(n_1074) );
INVxp67_ASAP7_75t_L g1075 ( .A(n_930), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_948), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1077 ( .A(n_934), .Y(n_1077) );
BUFx3_ASAP7_75t_L g1078 ( .A(n_939), .Y(n_1078) );
BUFx4f_ASAP7_75t_SL g1079 ( .A(n_1024), .Y(n_1079) );
OR2x6_ASAP7_75t_L g1080 ( .A(n_963), .B(n_936), .Y(n_1080) );
BUFx2_ASAP7_75t_L g1081 ( .A(n_983), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_920), .B(n_965), .Y(n_1082) );
BUFx4f_ASAP7_75t_SL g1083 ( .A(n_951), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_995), .B(n_924), .Y(n_1084) );
OAI21xp5_ASAP7_75t_L g1085 ( .A1(n_949), .A2(n_1006), .B(n_938), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_954), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_925), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_944), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_977), .B(n_991), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_997), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_977), .B(n_992), .Y(n_1091) );
OA21x2_ASAP7_75t_L g1092 ( .A1(n_994), .A2(n_981), .B(n_1025), .Y(n_1092) );
AO21x2_ASAP7_75t_L g1093 ( .A1(n_989), .A2(n_981), .B(n_972), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_953), .B(n_950), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_938), .B(n_957), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_937), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_993), .B(n_972), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_993), .B(n_942), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_945), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_1011), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_975), .B(n_946), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_969), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1011), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_973), .Y(n_1104) );
INVx2_ASAP7_75t_SL g1105 ( .A(n_1073), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1076), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1084), .B(n_982), .Y(n_1107) );
INVx4_ASAP7_75t_L g1108 ( .A(n_1073), .Y(n_1108) );
INVxp67_ASAP7_75t_L g1109 ( .A(n_1049), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1074), .Y(n_1110) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1054), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1067), .B(n_931), .Y(n_1112) );
INVxp67_ASAP7_75t_R g1113 ( .A(n_1067), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1044), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1044), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1034), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_1059), .Y(n_1117) );
INVx5_ASAP7_75t_L g1118 ( .A(n_1073), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1084), .B(n_982), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1072), .B(n_978), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_1051), .A2(n_929), .B1(n_968), .B2(n_933), .Y(n_1121) );
OR2x6_ASAP7_75t_SL g1122 ( .A(n_1064), .B(n_917), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1036), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1072), .B(n_978), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1068), .B(n_926), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1068), .B(n_926), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1095), .B(n_1091), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1095), .B(n_985), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1037), .Y(n_1129) );
BUFx4f_ASAP7_75t_L g1130 ( .A(n_1073), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1091), .B(n_941), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1061), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_1047), .B(n_985), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1040), .B(n_941), .Y(n_1134) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_1033), .Y(n_1135) );
AND2x4_ASAP7_75t_L g1136 ( .A(n_1070), .B(n_974), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1040), .B(n_980), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1047), .B(n_962), .Y(n_1138) );
OR2x2_ASAP7_75t_L g1139 ( .A(n_1052), .B(n_962), .Y(n_1139) );
INVxp67_ASAP7_75t_L g1140 ( .A(n_1043), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1042), .B(n_962), .Y(n_1141) );
BUFx2_ASAP7_75t_L g1142 ( .A(n_1081), .Y(n_1142) );
NAND2x1_ASAP7_75t_L g1143 ( .A(n_1081), .B(n_935), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1071), .B(n_1004), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1042), .B(n_955), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_1100), .Y(n_1146) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_1039), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1035), .B(n_1038), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_1075), .A2(n_960), .B1(n_955), .B2(n_959), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1035), .B(n_1004), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1052), .B(n_1089), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1056), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1038), .B(n_960), .Y(n_1153) );
INVx4_ASAP7_75t_L g1154 ( .A(n_1080), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1098), .B(n_935), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1062), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1098), .B(n_959), .Y(n_1157) );
AOI33xp33_ASAP7_75t_L g1158 ( .A1(n_1087), .A2(n_998), .A3(n_1026), .B1(n_940), .B2(n_970), .B3(n_956), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1066), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1160 ( .A(n_1077), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1090), .B(n_961), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1094), .B(n_1026), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1107), .B(n_1092), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1111), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1114), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1151), .B(n_1097), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g1167 ( .A(n_1142), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1114), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1107), .B(n_1092), .Y(n_1169) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_1142), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1115), .Y(n_1171) );
INVx3_ASAP7_75t_SL g1172 ( .A(n_1118), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1119), .B(n_1092), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1115), .Y(n_1174) );
AND2x4_ASAP7_75t_SL g1175 ( .A(n_1108), .B(n_1080), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1119), .B(n_1093), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1127), .B(n_1085), .Y(n_1177) );
BUFx2_ASAP7_75t_SL g1178 ( .A(n_1118), .Y(n_1178) );
NOR2x1_ASAP7_75t_L g1179 ( .A(n_1108), .B(n_1032), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1180 ( .A(n_1151), .B(n_1097), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1124), .B(n_1093), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1124), .B(n_1093), .Y(n_1182) );
NOR2xp67_ASAP7_75t_L g1183 ( .A(n_1118), .B(n_1050), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1127), .B(n_1069), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1120), .B(n_1048), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1120), .B(n_1094), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1138), .B(n_1045), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1125), .B(n_1048), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1189 ( .A(n_1135), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1126), .B(n_1065), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1148), .B(n_1088), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1131), .B(n_1065), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1131), .B(n_1065), .Y(n_1193) );
INVx1_ASAP7_75t_SL g1194 ( .A(n_1146), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1132), .B(n_1086), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1153), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1153), .Y(n_1197) );
INVx3_ASAP7_75t_L g1198 ( .A(n_1143), .Y(n_1198) );
AND2x4_ASAP7_75t_L g1199 ( .A(n_1136), .B(n_1141), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1134), .Y(n_1200) );
INVx3_ASAP7_75t_L g1201 ( .A(n_1198), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1163), .B(n_1157), .Y(n_1202) );
AOI21x1_ASAP7_75t_SL g1203 ( .A1(n_1189), .A2(n_1150), .B(n_1144), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1165), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1163), .B(n_1169), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1169), .B(n_1157), .Y(n_1206) );
INVxp67_ASAP7_75t_L g1207 ( .A(n_1170), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1177), .B(n_1117), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1173), .B(n_1155), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1177), .B(n_1147), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1168), .Y(n_1211) );
NOR2x1_ASAP7_75t_L g1212 ( .A(n_1179), .B(n_1108), .Y(n_1212) );
NAND3xp33_ASAP7_75t_L g1213 ( .A(n_1167), .B(n_1158), .C(n_1162), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1171), .Y(n_1214) );
AND2x4_ASAP7_75t_L g1215 ( .A(n_1199), .B(n_1136), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1196), .B(n_1116), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1173), .B(n_1155), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1176), .B(n_1145), .Y(n_1218) );
NOR2x1_ASAP7_75t_L g1219 ( .A(n_1179), .B(n_1162), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1164), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1176), .B(n_1145), .Y(n_1221) );
AND2x4_ASAP7_75t_L g1222 ( .A(n_1199), .B(n_1136), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1190), .B(n_1161), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1186), .B(n_1138), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1171), .Y(n_1225) );
NAND4xp25_ASAP7_75t_L g1226 ( .A(n_1187), .B(n_1063), .C(n_1121), .D(n_1112), .Y(n_1226) );
AND2x4_ASAP7_75t_L g1227 ( .A(n_1199), .B(n_1161), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1174), .Y(n_1228) );
INVxp67_ASAP7_75t_L g1229 ( .A(n_1170), .Y(n_1229) );
HB1xp67_ASAP7_75t_L g1230 ( .A(n_1167), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1190), .B(n_1139), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1185), .B(n_1139), .Y(n_1232) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1186), .B(n_1133), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1196), .B(n_1123), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_1194), .Y(n_1235) );
NAND2xp5_ASAP7_75t_SL g1236 ( .A(n_1172), .B(n_1130), .Y(n_1236) );
NAND2x1p5_ASAP7_75t_L g1237 ( .A(n_1183), .B(n_1130), .Y(n_1237) );
OR2x2_ASAP7_75t_L g1238 ( .A(n_1166), .B(n_1133), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1185), .B(n_1137), .Y(n_1239) );
INVx3_ASAP7_75t_L g1240 ( .A(n_1198), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1192), .B(n_1137), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1197), .B(n_1129), .Y(n_1242) );
HB1xp67_ASAP7_75t_L g1243 ( .A(n_1194), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1192), .B(n_1128), .Y(n_1244) );
AND2x4_ASAP7_75t_SL g1245 ( .A(n_1199), .B(n_1154), .Y(n_1245) );
NAND2xp5_ASAP7_75t_SL g1246 ( .A(n_1219), .B(n_1130), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1205), .B(n_1181), .Y(n_1247) );
INVx3_ASAP7_75t_L g1248 ( .A(n_1201), .Y(n_1248) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1208), .B(n_1140), .Y(n_1249) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1220), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1204), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1244), .B(n_1197), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1204), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1205), .B(n_1193), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1211), .Y(n_1255) );
NAND2x1_ASAP7_75t_SL g1256 ( .A(n_1212), .B(n_1172), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1211), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1233), .B(n_1181), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1233), .B(n_1182), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1244), .B(n_1184), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1214), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1214), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1231), .B(n_1184), .Y(n_1263) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1226), .B(n_1078), .Y(n_1264) );
INVx1_ASAP7_75t_SL g1265 ( .A(n_1245), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1209), .B(n_1193), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1210), .B(n_1078), .Y(n_1267) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_1213), .A2(n_1109), .B1(n_1096), .B2(n_1191), .C(n_1060), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1225), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g1270 ( .A(n_1235), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1225), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1231), .B(n_1200), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1241), .B(n_1200), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1238), .B(n_1182), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1228), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1216), .B(n_1083), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1258), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1266), .B(n_1223), .Y(n_1278) );
INVx2_ASAP7_75t_L g1279 ( .A(n_1250), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1276), .B(n_1234), .Y(n_1280) );
A2O1A1Ixp33_ASAP7_75t_L g1281 ( .A1(n_1264), .A2(n_1245), .B(n_1175), .C(n_1118), .Y(n_1281) );
INVxp67_ASAP7_75t_L g1282 ( .A(n_1270), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_1268), .A2(n_1113), .B1(n_1227), .B2(n_1188), .Y(n_1283) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_1246), .A2(n_1236), .B(n_1237), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1258), .Y(n_1285) );
AOI32xp33_ASAP7_75t_L g1286 ( .A1(n_1265), .A2(n_1232), .A3(n_1239), .B1(n_1175), .B2(n_1206), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1259), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1266), .B(n_1254), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_1267), .A2(n_1113), .B1(n_1227), .B2(n_1188), .Y(n_1289) );
INVxp67_ASAP7_75t_L g1290 ( .A(n_1249), .Y(n_1290) );
AOI22xp5_ASAP7_75t_L g1291 ( .A1(n_1252), .A2(n_1227), .B1(n_1215), .B2(n_1222), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1259), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1254), .B(n_1223), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1274), .B(n_1218), .Y(n_1294) );
OAI321xp33_ASAP7_75t_L g1295 ( .A1(n_1274), .A2(n_1237), .A3(n_1229), .B1(n_1207), .B2(n_1238), .C(n_1224), .Y(n_1295) );
AOI21xp5_ASAP7_75t_L g1296 ( .A1(n_1248), .A2(n_1237), .B(n_1175), .Y(n_1296) );
OAI221xp5_ASAP7_75t_L g1297 ( .A1(n_1248), .A2(n_1242), .B1(n_1230), .B2(n_1187), .C(n_1224), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_1260), .A2(n_1046), .B1(n_1053), .B2(n_1057), .Y(n_1298) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_1248), .A2(n_1191), .B1(n_1201), .B2(n_1240), .C(n_1243), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1282), .B(n_1218), .Y(n_1300) );
AOI221xp5_ASAP7_75t_L g1301 ( .A1(n_1295), .A2(n_1297), .B1(n_1282), .B2(n_1290), .C(n_1286), .Y(n_1301) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_1283), .A2(n_1247), .B1(n_1263), .B2(n_1256), .C(n_1272), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1277), .B(n_1221), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1285), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_1290), .A2(n_1292), .B1(n_1287), .B2(n_1280), .Y(n_1305) );
AOI22xp5_ASAP7_75t_L g1306 ( .A1(n_1291), .A2(n_1215), .B1(n_1222), .B2(n_1232), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1294), .Y(n_1307) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_1289), .A2(n_1222), .B1(n_1215), .B2(n_1273), .Y(n_1308) );
OAI21xp5_ASAP7_75t_L g1309 ( .A1(n_1284), .A2(n_1256), .B(n_1150), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1279), .Y(n_1310) );
AOI211xp5_ASAP7_75t_L g1311 ( .A1(n_1281), .A2(n_1172), .B(n_1150), .C(n_1041), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1288), .B(n_1202), .Y(n_1312) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_1299), .A2(n_1240), .B1(n_1201), .B2(n_1261), .C(n_1275), .Y(n_1313) );
AOI22xp5_ASAP7_75t_L g1314 ( .A1(n_1298), .A2(n_1239), .B1(n_1241), .B2(n_1206), .Y(n_1314) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_1298), .A2(n_1202), .B1(n_1217), .B2(n_1262), .Y(n_1315) );
NOR4xp25_ASAP7_75t_L g1316 ( .A(n_1293), .B(n_1110), .C(n_1106), .D(n_1156), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1278), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1296), .Y(n_1318) );
NAND2xp5_ASAP7_75t_SL g1319 ( .A(n_1295), .B(n_1240), .Y(n_1319) );
NOR3xp33_ASAP7_75t_L g1320 ( .A(n_1295), .B(n_1104), .C(n_1041), .Y(n_1320) );
NAND4xp75_ASAP7_75t_L g1321 ( .A(n_1283), .B(n_1105), .C(n_1183), .D(n_1101), .Y(n_1321) );
NOR2xp67_ASAP7_75t_SL g1322 ( .A(n_1284), .B(n_1178), .Y(n_1322) );
AOI211xp5_ASAP7_75t_L g1323 ( .A1(n_1295), .A2(n_1166), .B(n_1180), .C(n_1251), .Y(n_1323) );
AOI222xp33_ASAP7_75t_L g1324 ( .A1(n_1295), .A2(n_1257), .B1(n_1251), .B2(n_1253), .C1(n_1269), .C2(n_1255), .Y(n_1324) );
AOI221xp5_ASAP7_75t_SL g1325 ( .A1(n_1290), .A2(n_1217), .B1(n_1253), .B2(n_1269), .C(n_1255), .Y(n_1325) );
O2A1O1Ixp33_ASAP7_75t_SL g1326 ( .A1(n_1281), .A2(n_1105), .B(n_1122), .C(n_1203), .Y(n_1326) );
OAI211xp5_ASAP7_75t_SL g1327 ( .A1(n_1301), .A2(n_1324), .B(n_1320), .C(n_1323), .Y(n_1327) );
A2O1A1Ixp33_ASAP7_75t_L g1328 ( .A1(n_1309), .A2(n_1322), .B(n_1325), .C(n_1311), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1304), .Y(n_1329) );
NAND4xp75_ASAP7_75t_L g1330 ( .A(n_1319), .B(n_1318), .C(n_1308), .D(n_1306), .Y(n_1330) );
NAND4xp25_ASAP7_75t_L g1331 ( .A(n_1305), .B(n_1302), .C(n_1326), .D(n_1315), .Y(n_1331) );
NAND3x1_ASAP7_75t_SL g1332 ( .A(n_1079), .B(n_1316), .C(n_1321), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1317), .B(n_1307), .Y(n_1333) );
NOR3x1_ASAP7_75t_L g1334 ( .A(n_1313), .B(n_1300), .C(n_1303), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1333), .Y(n_1335) );
INVxp67_ASAP7_75t_L g1336 ( .A(n_1330), .Y(n_1336) );
NAND3xp33_ASAP7_75t_L g1337 ( .A(n_1327), .B(n_1314), .C(n_1310), .Y(n_1337) );
NAND4xp75_ASAP7_75t_L g1338 ( .A(n_1334), .B(n_1058), .C(n_1055), .D(n_1082), .Y(n_1338) );
NOR3xp33_ASAP7_75t_L g1339 ( .A(n_1331), .B(n_1058), .C(n_1055), .Y(n_1339) );
AND2x4_ASAP7_75t_L g1340 ( .A(n_1339), .B(n_1335), .Y(n_1340) );
NOR3xp33_ASAP7_75t_L g1341 ( .A(n_1336), .B(n_1332), .C(n_1328), .Y(n_1341) );
NOR2x1_ASAP7_75t_L g1342 ( .A(n_1338), .B(n_1329), .Y(n_1342) );
NOR2x1p5_ASAP7_75t_L g1343 ( .A(n_1337), .B(n_1312), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_1343), .A2(n_1341), .B1(n_1340), .B2(n_1342), .Y(n_1344) );
OAI22xp5_ASAP7_75t_SL g1345 ( .A1(n_1344), .A2(n_1031), .B1(n_1032), .B2(n_1178), .Y(n_1345) );
OR2x2_ASAP7_75t_L g1346 ( .A(n_1345), .B(n_1271), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1347 ( .A1(n_1346), .A2(n_1099), .B1(n_1102), .B2(n_1152), .C(n_1159), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_1347), .A2(n_1122), .B1(n_1160), .B2(n_1149), .Y(n_1348) );
HB1xp67_ASAP7_75t_L g1349 ( .A(n_1348), .Y(n_1349) );
AOI21xp5_ASAP7_75t_L g1350 ( .A1(n_1349), .A2(n_1103), .B(n_1195), .Y(n_1350) );
endmodule