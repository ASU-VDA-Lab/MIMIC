module fake_netlist_1_1290_n_599 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_599);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_599;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_28), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_11), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_14), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_30), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_59), .Y(n_78) );
INVxp67_ASAP7_75t_SL g79 ( .A(n_2), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_25), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_63), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_50), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_2), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_45), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_24), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_46), .Y(n_86) );
INVx2_ASAP7_75t_SL g87 ( .A(n_35), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_52), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_17), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_8), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_60), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
NOR2xp33_ASAP7_75t_L g93 ( .A(n_38), .B(n_10), .Y(n_93) );
BUFx2_ASAP7_75t_SL g94 ( .A(n_20), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_5), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_32), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_36), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_56), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_5), .Y(n_102) );
INVx3_ASAP7_75t_L g103 ( .A(n_16), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_14), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
INVxp33_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_62), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_44), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_48), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_37), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_57), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_19), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_8), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_75), .B(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_103), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_103), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_80), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_110), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_103), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_103), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_113), .B(n_0), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_113), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_92), .B(n_1), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_107), .B(n_1), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_113), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_77), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_110), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_77), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_117), .B(n_3), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_74), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_74), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_78), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_78), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_87), .B(n_4), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_117), .B(n_4), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_84), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_82), .Y(n_151) );
OR2x6_ASAP7_75t_L g152 ( .A(n_94), .B(n_31), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_84), .Y(n_154) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_88), .A2(n_33), .B(n_70), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_91), .B(n_6), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_115), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_85), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_91), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_85), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_128), .B(n_101), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_128), .B(n_95), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
AO22x2_ASAP7_75t_L g167 ( .A1(n_130), .A2(n_108), .B1(n_96), .B2(n_100), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_123), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_137), .B(n_130), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_124), .B(n_109), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_145), .B(n_121), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_125), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_145), .B(n_111), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_126), .B(n_116), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_122), .B(n_101), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_141), .B(n_83), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_148), .A2(n_76), .B(n_89), .C(n_90), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_141), .B(n_116), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_131), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_152), .B(n_76), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g196 ( .A1(n_158), .A2(n_102), .B1(n_127), .B2(n_138), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_143), .B(n_99), .Y(n_197) );
INVx1_ASAP7_75t_SL g198 ( .A(n_140), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_143), .B(n_120), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_122), .B(n_89), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_152), .B(n_105), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_146), .B(n_120), .Y(n_204) );
INVxp67_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_122), .B(n_90), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_152), .A2(n_105), .B1(n_106), .B2(n_79), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_150), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_139), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
NAND3xp33_ASAP7_75t_L g214 ( .A(n_133), .B(n_106), .C(n_118), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_136), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_134), .Y(n_216) );
AO22x2_ASAP7_75t_L g217 ( .A1(n_149), .A2(n_104), .B1(n_118), .B2(n_100), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_152), .A2(n_81), .B1(n_104), .B2(n_112), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_149), .B(n_112), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_136), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_151), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_136), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_136), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_198), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_180), .Y(n_226) );
NAND3xp33_ASAP7_75t_SL g227 ( .A(n_185), .B(n_133), .C(n_134), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_180), .Y(n_228) );
INVx4_ASAP7_75t_L g229 ( .A(n_195), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
OA22x2_ASAP7_75t_L g231 ( .A1(n_210), .A2(n_151), .B1(n_161), .B2(n_160), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_164), .B(n_161), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_163), .B(n_153), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_195), .B(n_153), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_195), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_203), .B(n_163), .Y(n_236) );
NOR2xp33_ASAP7_75t_R g237 ( .A(n_174), .B(n_160), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_203), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_171), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_174), .B(n_156), .Y(n_241) );
NAND2xp33_ASAP7_75t_SL g242 ( .A(n_174), .B(n_108), .Y(n_242) );
NOR3xp33_ASAP7_75t_SL g243 ( .A(n_196), .B(n_147), .C(n_93), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_216), .B(n_162), .Y(n_244) );
NOR2xp33_ASAP7_75t_R g245 ( .A(n_213), .B(n_162), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_171), .Y(n_246) );
AO22x1_ASAP7_75t_L g247 ( .A1(n_213), .A2(n_98), .B1(n_119), .B2(n_135), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_213), .B(n_86), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_199), .B(n_86), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_199), .B(n_86), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_163), .B(n_132), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_218), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_219), .B(n_162), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_180), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_219), .B(n_162), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_171), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_219), .B(n_150), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_207), .B(n_132), .Y(n_259) );
INVx5_ASAP7_75t_L g260 ( .A(n_165), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_205), .B(n_135), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_168), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_167), .A2(n_159), .B1(n_157), .B2(n_94), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_167), .A2(n_159), .B1(n_157), .B2(n_154), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_177), .B(n_159), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
INVx4_ASAP7_75t_L g267 ( .A(n_165), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_167), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_184), .B(n_157), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_175), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_167), .A2(n_154), .B1(n_144), .B2(n_155), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_187), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_168), .Y(n_273) );
OR2x6_ASAP7_75t_L g274 ( .A(n_207), .B(n_155), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_194), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_179), .B(n_114), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_183), .B(n_114), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_187), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_194), .Y(n_279) );
INVxp67_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_209), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_165), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_202), .B(n_154), .Y(n_283) );
BUFx5_ASAP7_75t_L g284 ( .A(n_170), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_209), .Y(n_285) );
INVx5_ASAP7_75t_L g286 ( .A(n_209), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_197), .B(n_114), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_202), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_225), .Y(n_290) );
AO32x2_ASAP7_75t_L g291 ( .A1(n_267), .A2(n_217), .A3(n_155), .B1(n_144), .B2(n_154), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_236), .B(n_186), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_284), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_284), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_235), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_236), .B(n_211), .Y(n_296) );
INVx5_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_234), .B(n_191), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_268), .A2(n_217), .B1(n_214), .B2(n_169), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_239), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_240), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_280), .A2(n_182), .B1(n_173), .B2(n_217), .C(n_221), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_268), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_240), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_248), .A2(n_193), .B(n_200), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_234), .B(n_217), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_239), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_289), .Y(n_310) );
BUFx4f_ASAP7_75t_L g311 ( .A(n_235), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_256), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_235), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_231), .A2(n_189), .B1(n_188), .B2(n_178), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_251), .B(n_204), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_237), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_237), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_256), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_238), .A2(n_189), .B1(n_178), .B2(n_188), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_235), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
OR2x6_ASAP7_75t_SL g323 ( .A(n_252), .B(n_170), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_259), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_238), .A2(n_176), .B1(n_211), .B2(n_222), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_226), .Y(n_328) );
NAND2xp33_ASAP7_75t_L g329 ( .A(n_230), .B(n_176), .Y(n_329) );
NAND3xp33_ASAP7_75t_L g330 ( .A(n_243), .B(n_222), .C(n_208), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_246), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_246), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_280), .B(n_212), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_277), .B(n_208), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_248), .A2(n_155), .B(n_212), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_277), .B(n_7), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_251), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_233), .B(n_9), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_312), .B(n_260), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_324), .B(n_259), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_290), .A2(n_337), .B1(n_310), .B2(n_318), .Y(n_342) );
BUFx10_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_333), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_308), .A2(n_264), .B1(n_263), .B2(n_253), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_304), .A2(n_231), .B1(n_227), .B2(n_267), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_297), .B(n_260), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_333), .B(n_232), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_227), .B1(n_261), .B2(n_260), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_339), .A2(n_264), .B1(n_255), .B2(n_258), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g353 ( .A1(n_303), .A2(n_243), .B(n_276), .C(n_287), .Y(n_353) );
AND2x2_ASAP7_75t_SL g354 ( .A(n_329), .B(n_241), .Y(n_354) );
NAND2xp33_ASAP7_75t_SL g355 ( .A(n_317), .B(n_245), .Y(n_355) );
AND2x6_ASAP7_75t_L g356 ( .A(n_337), .B(n_245), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_297), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_328), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_297), .Y(n_360) );
CKINVDCx14_ASAP7_75t_R g361 ( .A(n_323), .Y(n_361) );
INVxp67_ASAP7_75t_L g362 ( .A(n_323), .Y(n_362) );
INVx5_ASAP7_75t_L g363 ( .A(n_297), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_299), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_318), .B(n_299), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_328), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_311), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_316), .B(n_265), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_329), .A2(n_242), .B1(n_276), .B2(n_247), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_359), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_356), .A2(n_335), .B1(n_320), .B2(n_330), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_357), .A2(n_339), .B1(n_298), .B2(n_326), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_356), .A2(n_335), .B1(n_325), .B2(n_292), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_350), .B(n_335), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_342), .A2(n_315), .B(n_269), .C(n_300), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_361), .A2(n_338), .B1(n_283), .B2(n_332), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_341), .B(n_296), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_341), .A2(n_356), .B1(n_350), .B2(n_362), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_344), .A2(n_336), .B(n_271), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_368), .B(n_296), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_356), .A2(n_299), .B1(n_305), .B2(n_311), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_356), .A2(n_302), .B1(n_305), .B2(n_331), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_354), .A2(n_271), .B1(n_311), .B2(n_293), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_319), .B1(n_301), .B2(n_309), .C(n_313), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_363), .Y(n_387) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_356), .B(n_293), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_346), .B(n_305), .Y(n_389) );
OAI22xp33_ASAP7_75t_L g390 ( .A1(n_369), .A2(n_302), .B1(n_327), .B2(n_322), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_351), .A2(n_348), .B1(n_346), .B2(n_352), .C(n_347), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_344), .A2(n_307), .B(n_327), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_356), .A2(n_282), .B1(n_260), .B2(n_266), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_354), .A2(n_282), .B1(n_275), .B2(n_279), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_366), .B(n_286), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_366), .B(n_286), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_365), .B1(n_364), .B2(n_360), .C(n_281), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_370), .B(n_380), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_390), .A2(n_249), .B(n_250), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_380), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_381), .B(n_367), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_381), .B(n_343), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_376), .A2(n_360), .B(n_363), .C(n_364), .Y(n_404) );
AOI21xp5_ASAP7_75t_SL g405 ( .A1(n_384), .A2(n_354), .B(n_345), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_355), .B1(n_364), .B2(n_343), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_387), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_374), .B(n_343), .Y(n_408) );
AOI33xp33_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_285), .A3(n_215), .B1(n_201), .B2(n_181), .B3(n_220), .Y(n_409) );
NOR2xp33_ASAP7_75t_SL g410 ( .A(n_389), .B(n_363), .Y(n_410) );
OAI31xp33_ASAP7_75t_SL g411 ( .A1(n_375), .A2(n_349), .A3(n_340), .B(n_249), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_395), .B(n_291), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_363), .B1(n_358), .B2(n_349), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_377), .B(n_250), .C(n_358), .D(n_201), .Y(n_414) );
OAI33xp33_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_172), .A3(n_220), .B1(n_215), .B2(n_190), .B3(n_181), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_385), .B(n_363), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_389), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_395), .B(n_291), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_371), .B(n_363), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_396), .B(n_291), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_371), .A2(n_349), .B1(n_358), .B2(n_345), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_382), .B(n_349), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_385), .B(n_291), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_383), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_394), .B(n_345), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g429 ( .A1(n_388), .A2(n_166), .A3(n_172), .B1(n_190), .B2(n_288), .B3(n_15), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_385), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_385), .B(n_291), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_421), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_399), .B(n_412), .Y(n_433) );
INVx4_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_407), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_424), .A2(n_154), .B1(n_144), .B2(n_393), .C(n_388), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_397), .B(n_379), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g438 ( .A1(n_404), .A2(n_340), .A3(n_334), .B(n_321), .Y(n_438) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_411), .A2(n_345), .B(n_340), .C(n_144), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_421), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_401), .B(n_392), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_426), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_417), .B(n_392), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_416), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_412), .B(n_155), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_431), .A2(n_166), .B(n_254), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_417), .B(n_144), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_431), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_398), .A2(n_340), .B1(n_334), .B2(n_274), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_402), .A2(n_9), .A3(n_10), .B1(n_12), .B2(n_13), .B3(n_15), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_419), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_427), .A2(n_274), .B1(n_144), .B2(n_154), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_430), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_410), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_418), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_422), .B(n_274), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_420), .B(n_66), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_409), .B(n_175), .C(n_223), .Y(n_461) );
OAI33xp33_ASAP7_75t_L g462 ( .A1(n_414), .A2(n_12), .A3(n_13), .B1(n_17), .B2(n_228), .B3(n_272), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_425), .B(n_322), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_405), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_405), .Y(n_466) );
NOR3xp33_ASAP7_75t_SL g467 ( .A(n_403), .B(n_18), .C(n_21), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_400), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_413), .B(n_314), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_400), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_428), .B(n_314), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_400), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_408), .B(n_23), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_429), .B(n_26), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_415), .A2(n_314), .B1(n_295), .B2(n_321), .Y(n_476) );
AOI221xp5_ASAP7_75t_SL g477 ( .A1(n_424), .A2(n_175), .B1(n_192), .B2(n_206), .C(n_223), .Y(n_477) );
NAND2xp33_ASAP7_75t_R g478 ( .A(n_467), .B(n_27), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_433), .B(n_295), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_457), .B(n_223), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
INVx5_ASAP7_75t_L g482 ( .A(n_434), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_457), .B(n_223), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_474), .A2(n_262), .B1(n_273), .B2(n_286), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_458), .B(n_29), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_457), .B(n_223), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_439), .B(n_224), .C(n_273), .D(n_278), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_435), .B(n_34), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_448), .B(n_206), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_455), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_435), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_442), .B(n_206), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_434), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_442), .B(n_206), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_434), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_442), .B(n_192), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_452), .B(n_39), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_440), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_434), .Y(n_505) );
NAND2xp33_ASAP7_75t_SL g506 ( .A(n_460), .B(n_450), .Y(n_506) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_460), .B(n_294), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_459), .B(n_40), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_437), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_465), .B(n_224), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_459), .B(n_42), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_437), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_444), .B(n_47), .Y(n_513) );
NOR2xp33_ASAP7_75t_SL g514 ( .A(n_438), .B(n_294), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_441), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_509), .B(n_443), .Y(n_516) );
AOI321xp33_ASAP7_75t_SL g517 ( .A1(n_490), .A2(n_456), .A3(n_452), .B1(n_462), .B2(n_475), .C(n_461), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_501), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_496), .B(n_461), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_512), .B(n_443), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_505), .B(n_449), .Y(n_521) );
AOI31xp33_ASAP7_75t_L g522 ( .A1(n_499), .A2(n_462), .A3(n_436), .B(n_477), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_506), .A2(n_436), .B(n_464), .C(n_466), .Y(n_523) );
NAND4xp25_ASAP7_75t_SL g524 ( .A(n_508), .B(n_477), .C(n_466), .D(n_475), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_501), .B(n_453), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_507), .A2(n_444), .B1(n_449), .B2(n_460), .Y(n_526) );
OAI21xp33_ASAP7_75t_L g527 ( .A1(n_494), .A2(n_463), .B(n_453), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_499), .A2(n_444), .B1(n_449), .B2(n_460), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_482), .A2(n_444), .B1(n_449), .B2(n_473), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_503), .A2(n_463), .B1(n_473), .B2(n_469), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_486), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_503), .A2(n_472), .B1(n_470), .B2(n_468), .C(n_445), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_482), .A2(n_454), .B1(n_469), .B2(n_471), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
AOI222xp33_ASAP7_75t_L g535 ( .A1(n_490), .A2(n_445), .B1(n_472), .B2(n_470), .C1(n_468), .C2(n_471), .Y(n_535) );
OAI222xp33_ASAP7_75t_L g536 ( .A1(n_482), .A2(n_472), .B1(n_470), .B2(n_468), .C1(n_476), .C2(n_446), .Y(n_536) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_514), .A2(n_306), .B(n_446), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_489), .B(n_446), .C(n_306), .Y(n_538) );
AOI211xp5_ASAP7_75t_L g539 ( .A1(n_508), .A2(n_49), .B(n_51), .C(n_54), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_479), .B(n_58), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_498), .B(n_446), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_482), .B(n_61), .Y(n_542) );
AOI211xp5_ASAP7_75t_L g543 ( .A1(n_511), .A2(n_65), .B(n_67), .C(n_68), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_492), .B(n_257), .C(n_270), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_502), .B(n_71), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_515), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_478), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_513), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_531), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_534), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_546), .Y(n_551) );
INVx2_ASAP7_75t_SL g552 ( .A(n_525), .Y(n_552) );
NAND2x1p5_ASAP7_75t_SL g553 ( .A(n_519), .B(n_480), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_516), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_547), .B(n_487), .Y(n_556) );
AOI211x1_ASAP7_75t_L g557 ( .A1(n_522), .A2(n_510), .B(n_495), .C(n_500), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_521), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_518), .B(n_491), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_528), .A2(n_484), .B1(n_488), .B2(n_483), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_535), .B(n_481), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_548), .B(n_485), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_542), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_532), .B(n_480), .C(n_483), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_527), .B(n_485), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_541), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_554), .B(n_532), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_556), .A2(n_524), .B1(n_526), .B2(n_530), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_554), .B(n_523), .Y(n_569) );
XOR2xp5_ASAP7_75t_L g570 ( .A(n_558), .B(n_529), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_555), .B(n_504), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_556), .A2(n_533), .B1(n_540), .B2(n_538), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_561), .Y(n_573) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_552), .B(n_539), .Y(n_574) );
OAI31xp33_ASAP7_75t_L g575 ( .A1(n_563), .A2(n_537), .A3(n_536), .B(n_545), .Y(n_575) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_564), .A2(n_543), .B(n_544), .C(n_517), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_566), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_567), .A2(n_557), .B1(n_553), .B2(n_549), .C(n_550), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_577), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_574), .Y(n_580) );
INVxp33_ASAP7_75t_SL g581 ( .A(n_570), .Y(n_581) );
AND2x2_ASAP7_75t_SL g582 ( .A(n_567), .B(n_565), .Y(n_582) );
AOI211xp5_ASAP7_75t_L g583 ( .A1(n_575), .A2(n_562), .B(n_559), .C(n_551), .Y(n_583) );
INVxp33_ASAP7_75t_SL g584 ( .A(n_568), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_576), .A2(n_497), .B1(n_560), .B2(n_572), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_571), .A2(n_570), .B1(n_573), .B2(n_568), .Y(n_586) );
OA22x2_ASAP7_75t_L g587 ( .A1(n_573), .A2(n_570), .B1(n_568), .B2(n_569), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_579), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_585), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_580), .Y(n_590) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_578), .B(n_582), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_589), .B(n_578), .C(n_583), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_588), .Y(n_593) );
XOR2xp5_ASAP7_75t_L g594 ( .A(n_590), .B(n_581), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_593), .Y(n_595) );
XNOR2xp5_ASAP7_75t_L g596 ( .A(n_594), .B(n_587), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_595), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_597), .A2(n_596), .B1(n_584), .B2(n_592), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_598), .A2(n_591), .B(n_586), .Y(n_599) );
endmodule