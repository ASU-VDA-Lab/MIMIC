module fake_jpeg_28826_n_111 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_SL g11 ( 
.A(n_9),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_2),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_44),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_20),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_54),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_30),
.C(n_24),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_58),
.B(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_10),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_13),
.B1(n_17),
.B2(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_5),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_59),
.B1(n_61),
.B2(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_17),
.B1(n_7),
.B2(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_33),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_67),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_10),
.C(n_33),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_78),
.B(n_83),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_48),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_55),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_62),
.C(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_56),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_71),
.B(n_65),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_92),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_91),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_62),
.B(n_73),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_70),
.B(n_74),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_80),
.C(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_75),
.C(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_77),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_66),
.CI(n_70),
.CON(n_101),
.SN(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_95),
.B(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_99),
.B1(n_66),
.B2(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.C(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_98),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_56),
.B(n_52),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_52),
.Y(n_111)
);


endmodule