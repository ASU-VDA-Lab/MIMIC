module fake_jpeg_1634_n_681 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_681);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_681;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_574;
wire n_542;
wire n_313;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_61),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_66),
.Y(n_225)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_69),
.A2(n_46),
.B1(n_55),
.B2(n_50),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_9),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_79),
.Y(n_136)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_72),
.Y(n_133)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_77),
.Y(n_178)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_10),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_87),
.Y(n_163)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_98),
.Y(n_179)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_10),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_121),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_104),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx5_ASAP7_75t_SL g203 ( 
.A(n_105),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_42),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_20),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_111),
.Y(n_194)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_115),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

HAxp5_ASAP7_75t_SL g125 ( 
.A(n_25),
.B(n_0),
.CON(n_125),
.SN(n_125)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_125),
.B(n_0),
.CON(n_186),
.SN(n_186)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_41),
.Y(n_221)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_39),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_138),
.B(n_147),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_39),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_152),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_66),
.B(n_56),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_157),
.B(n_165),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_52),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_164),
.B(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_48),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_48),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_167),
.B(n_172),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_70),
.A2(n_55),
.B1(n_50),
.B2(n_31),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_170),
.A2(n_213),
.B1(n_1),
.B2(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_86),
.B(n_56),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_72),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_46),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_175),
.B(n_181),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_125),
.A2(n_57),
.B1(n_49),
.B2(n_44),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_180),
.A2(n_191),
.B1(n_196),
.B2(n_226),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_91),
.B(n_44),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_186),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_100),
.B(n_25),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_120),
.A2(n_57),
.B1(n_49),
.B2(n_21),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_130),
.A2(n_57),
.B1(n_49),
.B2(n_21),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_33),
.B1(n_87),
.B2(n_89),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_95),
.B(n_55),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_96),
.B(n_50),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_92),
.B(n_31),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_201),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_97),
.B(n_57),
.C(n_41),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_206),
.B(n_4),
.C(n_5),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_124),
.B(n_13),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_209),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_126),
.B(n_13),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_103),
.A2(n_41),
.B1(n_33),
.B2(n_29),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_76),
.B(n_81),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_73),
.A2(n_33),
.B1(n_29),
.B2(n_12),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_147),
.A2(n_107),
.B1(n_129),
.B2(n_128),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_235),
.Y(n_353)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_175),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_237),
.B(n_303),
.Y(n_316)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_131),
.B1(n_106),
.B2(n_127),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_240),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_334)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_182),
.A2(n_109),
.B1(n_122),
.B2(n_117),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_183),
.A2(n_116),
.B1(n_115),
.B2(n_129),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_193),
.A2(n_107),
.B1(n_69),
.B2(n_87),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_136),
.B(n_160),
.CI(n_186),
.CON(n_246),
.SN(n_246)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_246),
.B(n_173),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_248),
.A2(n_220),
.B1(n_192),
.B2(n_208),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_249),
.A2(n_253),
.B1(n_262),
.B2(n_275),
.Y(n_367)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_156),
.B(n_1),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_252),
.B(n_256),
.Y(n_323)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_151),
.Y(n_254)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_254),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_189),
.A2(n_12),
.B1(n_18),
.B2(n_17),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_255),
.A2(n_267),
.B1(n_279),
.B2(n_283),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_168),
.B(n_1),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_142),
.Y(n_257)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_257),
.Y(n_369)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_150),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_161),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_260),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_191),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_166),
.Y(n_265)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_265),
.Y(n_340)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_194),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_2),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_268),
.B(n_269),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_139),
.B(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_270),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_149),
.Y(n_272)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_274),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_196),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_179),
.Y(n_277)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_195),
.A2(n_218),
.B1(n_178),
.B2(n_169),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_291),
.Y(n_317)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_169),
.Y(n_282)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_282),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_13),
.B1(n_16),
.B2(n_6),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_284),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_226),
.A2(n_8),
.B1(n_13),
.B2(n_15),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_286),
.A2(n_261),
.B1(n_268),
.B2(n_231),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_178),
.A2(n_8),
.B1(n_19),
.B2(n_4),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_133),
.A2(n_5),
.B1(n_19),
.B2(n_146),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_133),
.A2(n_5),
.B1(n_148),
.B2(n_185),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_134),
.A2(n_220),
.B1(n_137),
.B2(n_140),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_204),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_293),
.Y(n_328)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_145),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_295),
.Y(n_342)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_211),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_197),
.A2(n_225),
.B1(n_205),
.B2(n_155),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_296),
.A2(n_297),
.B1(n_210),
.B2(n_203),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_134),
.A2(n_184),
.B1(n_137),
.B2(n_140),
.Y(n_297)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_135),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_307),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_197),
.B(n_214),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_278),
.C(n_248),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_162),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_187),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_270),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_159),
.B(n_190),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_305),
.B(n_306),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_171),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_159),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_314),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_241),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_309),
.B(n_324),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_276),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_230),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_247),
.B(n_225),
.C(n_200),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_327),
.C(n_364),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_321),
.B(n_338),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_263),
.B(n_223),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_247),
.B(n_173),
.C(n_144),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_261),
.A2(n_203),
.B(n_141),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_329),
.A2(n_277),
.B(n_282),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_SL g413 ( 
.A1(n_332),
.A2(n_358),
.B(n_365),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_234),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_333),
.B(n_339),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_250),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g341 ( 
.A1(n_271),
.A2(n_141),
.B(n_190),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_341),
.B(n_347),
.Y(n_410)
);

AO22x1_ASAP7_75t_L g346 ( 
.A1(n_261),
.A2(n_184),
.B1(n_143),
.B2(n_153),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_233),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_229),
.B(n_141),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_361),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_252),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_354),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_299),
.A2(n_143),
.B1(n_153),
.B2(n_154),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_256),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_360),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_285),
.B(n_187),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_154),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_232),
.B(n_192),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_367),
.A2(n_253),
.B1(n_300),
.B2(n_281),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_372),
.A2(n_405),
.B1(n_346),
.B2(n_359),
.Y(n_443)
);

A2O1A1O1Ixp25_ASAP7_75t_L g373 ( 
.A1(n_311),
.A2(n_246),
.B(n_280),
.C(n_269),
.D(n_302),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_373),
.A2(n_392),
.B(n_400),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_321),
.A2(n_300),
.B1(n_281),
.B2(n_249),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_276),
.C(n_264),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_386),
.C(n_397),
.Y(n_422)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_329),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_382),
.B(n_396),
.Y(n_449)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_367),
.A2(n_262),
.B1(n_275),
.B2(n_305),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_404),
.B1(n_414),
.B2(n_308),
.Y(n_424)
);

AO22x1_ASAP7_75t_SL g387 ( 
.A1(n_317),
.A2(n_266),
.B1(n_259),
.B2(n_258),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_399),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_351),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_391),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_353),
.A2(n_246),
.B1(n_291),
.B2(n_295),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_228),
.C(n_265),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_398),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_323),
.B(n_227),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_353),
.A2(n_293),
.B1(n_292),
.B2(n_274),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_401),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_323),
.B(n_236),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_403),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_257),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_360),
.A2(n_284),
.B1(n_301),
.B2(n_307),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_317),
.A2(n_208),
.B1(n_251),
.B2(n_239),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_345),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_406),
.B(n_412),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_228),
.C(n_238),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_407),
.B(n_350),
.C(n_359),
.Y(n_440)
);

OA22x2_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_242),
.B1(n_304),
.B2(n_260),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_409),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_349),
.B(n_254),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_334),
.A2(n_272),
.B1(n_273),
.B2(n_294),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_411),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_337),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_334),
.A2(n_319),
.B1(n_348),
.B2(n_316),
.Y(n_414)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_418),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_349),
.B(n_327),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_339),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_328),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_385),
.A2(n_319),
.B1(n_331),
.B2(n_314),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_419),
.A2(n_413),
.B1(n_377),
.B2(n_375),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_382),
.A2(n_308),
.B(n_315),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_420),
.A2(n_401),
.B(n_373),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_325),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_423),
.B(n_440),
.C(n_397),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_424),
.A2(n_443),
.B1(n_446),
.B2(n_447),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

INVx11_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_384),
.B(n_324),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_441),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_415),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_412),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_436),
.Y(n_490)
);

OAI32xp33_ASAP7_75t_L g437 ( 
.A1(n_410),
.A2(n_344),
.A3(n_325),
.B1(n_357),
.B2(n_346),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_403),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_395),
.B(n_350),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_444),
.B(n_445),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_372),
.A2(n_356),
.B1(n_357),
.B2(n_342),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_377),
.A2(n_356),
.B1(n_342),
.B2(n_363),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_409),
.B(n_340),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_448),
.B(n_453),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_390),
.B(n_342),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_451),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_343),
.Y(n_453)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_391),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_378),
.B(n_380),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_386),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_449),
.B(n_420),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_461),
.A2(n_462),
.B(n_465),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_449),
.A2(n_400),
.B(n_388),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_467),
.B1(n_468),
.B2(n_479),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_428),
.A2(n_441),
.B(n_450),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_428),
.A2(n_388),
.B(n_374),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_466),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_424),
.A2(n_399),
.B1(n_402),
.B2(n_394),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_443),
.A2(n_376),
.B1(n_392),
.B2(n_389),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_475),
.C(n_477),
.Y(n_506)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_473),
.Y(n_503)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_474),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_476),
.A2(n_445),
.B(n_432),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_407),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_478),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_419),
.A2(n_375),
.B1(n_376),
.B2(n_389),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_434),
.B(n_375),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_454),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_482),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_423),
.C(n_422),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_488),
.C(n_440),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_435),
.A2(n_405),
.B1(n_370),
.B2(n_404),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_484),
.A2(n_486),
.B1(n_494),
.B2(n_497),
.Y(n_530)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_447),
.A2(n_371),
.B1(n_406),
.B2(n_408),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_423),
.B(n_387),
.C(n_355),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_435),
.B(n_408),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_489),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_422),
.B(n_387),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_453),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_442),
.A2(n_408),
.B1(n_416),
.B2(n_355),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_457),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_457),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_425),
.A2(n_340),
.B1(n_343),
.B2(n_312),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_490),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_499),
.B(n_500),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_480),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_460),
.A2(n_434),
.B1(n_426),
.B2(n_425),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_501),
.A2(n_519),
.B1(n_479),
.B2(n_502),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_505),
.B(n_529),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_463),
.Y(n_507)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_509),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_448),
.Y(n_510)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_496),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_515),
.B(n_517),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_526),
.C(n_475),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_465),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_426),
.B1(n_446),
.B2(n_454),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_492),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_472),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_451),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_522),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_467),
.A2(n_442),
.B1(n_458),
.B2(n_459),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_523),
.A2(n_312),
.B1(n_368),
.B2(n_352),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_524),
.B(n_506),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_492),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_527),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_483),
.B(n_458),
.C(n_459),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_461),
.Y(n_527)
);

OAI22x1_ASAP7_75t_L g528 ( 
.A1(n_489),
.A2(n_437),
.B1(n_452),
.B2(n_439),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_528),
.A2(n_531),
.B1(n_487),
.B2(n_489),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_470),
.B(n_439),
.Y(n_529)
);

HB1xp67_ASAP7_75t_SL g531 ( 
.A(n_488),
.Y(n_531)
);

FAx1_ASAP7_75t_SL g532 ( 
.A(n_481),
.B(n_433),
.CI(n_436),
.CON(n_532),
.SN(n_532)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_532),
.B(n_474),
.Y(n_558)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_473),
.Y(n_533)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_533),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_477),
.B(n_421),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_534),
.B(n_478),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_535),
.B(n_565),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_539),
.A2(n_551),
.B1(n_554),
.B2(n_563),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_546),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_542),
.B(n_558),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_512),
.A2(n_487),
.B1(n_489),
.B2(n_495),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_543),
.A2(n_567),
.B1(n_513),
.B2(n_518),
.Y(n_591)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_502),
.Y(n_547)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_547),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_516),
.B(n_493),
.C(n_469),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_553),
.C(n_556),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_501),
.A2(n_464),
.B1(n_466),
.B2(n_462),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_506),
.B(n_469),
.C(n_476),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_519),
.A2(n_484),
.B1(n_497),
.B2(n_463),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_427),
.C(n_421),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_557),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_509),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_559),
.B(n_515),
.Y(n_578)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_504),
.Y(n_561)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_561),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_562),
.B(n_524),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_525),
.A2(n_485),
.B1(n_471),
.B2(n_482),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_526),
.B(n_429),
.C(n_471),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_564),
.B(n_527),
.C(n_507),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_529),
.B(n_429),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_504),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_566),
.B(n_533),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_570),
.B(n_556),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_540),
.A2(n_517),
.B(n_512),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_571),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_521),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_573),
.B(n_581),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_574),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g576 ( 
.A(n_549),
.B(n_553),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_576),
.B(n_582),
.Y(n_597)
);

CKINVDCx14_ASAP7_75t_R g611 ( 
.A(n_578),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_538),
.B(n_521),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_550),
.B(n_491),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_538),
.B(n_505),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_583),
.B(n_586),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_498),
.C(n_530),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_588),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_552),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_549),
.B(n_491),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_589),
.B(n_590),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_558),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_591),
.A2(n_539),
.B1(n_554),
.B2(n_551),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_548),
.B(n_523),
.C(n_513),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_593),
.C(n_565),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_535),
.B(n_528),
.C(n_510),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_604),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_537),
.Y(n_596)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_596),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_575),
.A2(n_541),
.B1(n_543),
.B2(n_536),
.Y(n_599)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_573),
.B(n_562),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_601),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_575),
.A2(n_536),
.B1(n_545),
.B2(n_567),
.Y(n_602)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_602),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_603),
.A2(n_577),
.B1(n_571),
.B2(n_587),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_574),
.B(n_563),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_606),
.B(n_544),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_570),
.B(n_540),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_608),
.B(n_393),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_592),
.C(n_569),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_609),
.B(n_610),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_572),
.B(n_545),
.C(n_508),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_532),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_612),
.B(n_579),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_577),
.A2(n_566),
.B1(n_561),
.B2(n_555),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_518),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_569),
.B(n_508),
.C(n_557),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_615),
.B(n_568),
.C(n_585),
.Y(n_622)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_617),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_598),
.A2(n_583),
.B1(n_581),
.B2(n_580),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_619),
.A2(n_621),
.B1(n_631),
.B2(n_632),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_607),
.A2(n_532),
.B(n_580),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_620),
.A2(n_623),
.B(n_597),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_607),
.A2(n_606),
.B1(n_603),
.B2(n_611),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_622),
.B(n_634),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_612),
.A2(n_568),
.B(n_584),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_626),
.B(n_604),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_630),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_613),
.A2(n_560),
.B1(n_514),
.B2(n_579),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_605),
.A2(n_560),
.B1(n_514),
.B2(n_368),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_633),
.B(n_601),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_610),
.B(n_335),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_637),
.A2(n_310),
.B(n_369),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_616),
.B(n_615),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_639),
.B(n_641),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_618),
.B(n_600),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_609),
.C(n_600),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_642),
.B(n_643),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_629),
.B(n_594),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_627),
.B(n_594),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_644),
.B(n_645),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_625),
.B(n_595),
.C(n_608),
.Y(n_645)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_646),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_647),
.B(n_648),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_624),
.B(n_335),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_617),
.B(n_352),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_649),
.B(n_310),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_637),
.A2(n_620),
.B(n_623),
.Y(n_650)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_650),
.B(n_638),
.C(n_646),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_636),
.A2(n_628),
.B1(n_621),
.B2(n_630),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_652),
.B(n_654),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_640),
.B(n_622),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_642),
.B(n_632),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_659),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_635),
.A2(n_619),
.B1(n_631),
.B2(n_633),
.Y(n_659)
);

OAI21x1_ASAP7_75t_SL g667 ( 
.A1(n_660),
.A2(n_661),
.B(n_635),
.Y(n_667)
);

AOI21x1_ASAP7_75t_L g672 ( 
.A1(n_662),
.A2(n_667),
.B(n_653),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_656),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_663),
.B(n_665),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_651),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_655),
.A2(n_638),
.B(n_645),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_666),
.A2(n_668),
.B(n_336),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_650),
.A2(n_369),
.B(n_322),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_664),
.A2(n_658),
.B(n_652),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_671),
.A2(n_672),
.B(n_673),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g673 ( 
.A(n_669),
.B(n_660),
.C(n_659),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_336),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_675),
.A2(n_677),
.B1(n_313),
.B2(n_318),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_670),
.B(n_322),
.Y(n_677)
);

BUFx24_ASAP7_75t_SL g679 ( 
.A(n_678),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_676),
.Y(n_680)
);

XOR2xp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_313),
.Y(n_681)
);


endmodule