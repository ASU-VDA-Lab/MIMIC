module fake_jpeg_29934_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_1),
.C(n_2),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_31),
.B(n_35),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_74),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_41),
.B1(n_52),
.B2(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_47),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_3),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_55),
.B1(n_54),
.B2(n_53),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_51),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_50),
.B1(n_42),
.B2(n_52),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_66),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_2),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_102),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_66),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_100),
.C(n_7),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_21),
.B(n_38),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_19),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_104),
.C(n_13),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_18),
.B1(n_37),
.B2(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_98),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_4),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_110),
.C(n_97),
.Y(n_116)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_11),
.C(n_12),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_106),
.C(n_114),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_96),
.C(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_98),
.C(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_122),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_114),
.B(n_95),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_123),
.A3(n_120),
.B1(n_115),
.B2(n_95),
.C1(n_118),
.C2(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_14),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_15),
.C(n_22),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_26),
.Y(n_128)
);

OAI221xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.C(n_33),
.Y(n_129)
);


endmodule