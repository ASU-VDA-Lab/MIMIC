module real_jpeg_28788_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_71),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_0),
.A2(n_25),
.B1(n_28),
.B2(n_71),
.Y(n_168)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_25),
.B1(n_28),
.B2(n_39),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_25),
.B1(n_28),
.B2(n_56),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_7),
.A2(n_74),
.B1(n_75),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_7),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_83),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_83),
.Y(n_182)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_9),
.B(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_63),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_63),
.B(n_131),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_76),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_9),
.A2(n_25),
.B(n_29),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_9),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_9),
.A2(n_41),
.B1(n_44),
.B2(n_182),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_12),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_25),
.B1(n_28),
.B2(n_69),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_66),
.Y(n_67)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_14),
.Y(n_130)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_103),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_34),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_24),
.A2(n_36),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_24),
.A2(n_36),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_24),
.A2(n_36),
.B1(n_138),
.B2(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_24),
.B(n_76),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_27),
.A2(n_32),
.B(n_76),
.C(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_28),
.B(n_187),
.Y(n_186)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_31),
.A2(n_64),
.A3(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_32),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_54),
.B(n_57),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_36),
.A2(n_139),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_45),
.B(n_47),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_41),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_41),
.A2(n_174),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_42),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_42),
.A2(n_48),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_42),
.A2(n_43),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_43),
.B(n_126),
.Y(n_169)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_43),
.Y(n_183)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_102),
.B(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.C(n_72),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_55),
.B(n_58),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_67),
.B1(n_111),
.B2(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_73),
.B1(n_80),
.B2(n_100),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.CON(n_73),
.SN(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_78),
.Y(n_80)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_76),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_98),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.C(n_109),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_104),
.A2(n_105),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_114),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_200),
.B(n_206),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_150),
.B(n_199),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_140),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_122),
.B(n_140),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_133),
.C(n_136),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_123),
.A2(n_124),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_127),
.Y(n_147)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_147),
.C(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_193),
.B(n_198),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_170),
.B(n_192),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_153),
.B(n_160),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_166),
.C(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_168),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_178),
.B(n_191),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_176),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_190),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_201),
.B(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);


endmodule