module real_jpeg_30655_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_0),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_0),
.A2(n_114),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_0),
.A2(n_114),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_0),
.A2(n_114),
.B1(n_471),
.B2(n_474),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_1),
.Y(n_206)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_1),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_1),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_1),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_3),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_3),
.A2(n_234),
.B1(n_338),
.B2(n_341),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_3),
.A2(n_234),
.B1(n_412),
.B2(n_415),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_3),
.A2(n_234),
.B1(n_539),
.B2(n_540),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_4),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_4),
.A2(n_69),
.B1(n_368),
.B2(n_373),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_4),
.A2(n_69),
.B1(n_187),
.B2(n_495),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_4),
.A2(n_69),
.B1(n_556),
.B2(n_559),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_5),
.A2(n_273),
.B1(n_278),
.B2(n_280),
.Y(n_272)
);

INVx2_ASAP7_75t_R g280 ( 
.A(n_5),
.Y(n_280)
);

AO22x1_ASAP7_75t_L g347 ( 
.A1(n_5),
.A2(n_280),
.B1(n_348),
.B2(n_351),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_5),
.A2(n_280),
.B1(n_423),
.B2(n_427),
.Y(n_422)
);

AO22x1_ASAP7_75t_L g530 ( 
.A1(n_5),
.A2(n_280),
.B1(n_531),
.B2(n_533),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_5),
.A2(n_280),
.B1(n_552),
.B2(n_553),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_6),
.A2(n_251),
.B1(n_253),
.B2(n_256),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_6),
.A2(n_256),
.B1(n_308),
.B2(n_313),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_6),
.A2(n_256),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_6),
.A2(n_256),
.B1(n_488),
.B2(n_490),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_7),
.A2(n_300),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_7),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_7),
.A2(n_325),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_7),
.A2(n_325),
.B1(n_499),
.B2(n_501),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_7),
.A2(n_70),
.B1(n_325),
.B2(n_549),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_8),
.A2(n_146),
.B1(n_148),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_150),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_8),
.A2(n_150),
.B1(n_219),
.B2(n_520),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_9),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_11),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_11),
.Y(n_277)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_11),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_76),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_106),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_12),
.A2(n_106),
.B1(n_435),
.B2(n_437),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_12),
.A2(n_106),
.B1(n_514),
.B2(n_516),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_16),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_14),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_15),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_15),
.A2(n_61),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_15),
.A2(n_61),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_18),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_18),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_19),
.A2(n_208),
.B1(n_250),
.B2(n_257),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_19),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_19),
.B(n_144),
.Y(n_354)
);

OAI32xp33_ASAP7_75t_L g375 ( 
.A1(n_19),
.A2(n_128),
.A3(n_376),
.B1(n_378),
.B2(n_382),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_19),
.A2(n_264),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_19),
.B(n_235),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_19),
.A2(n_464),
.B(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_240),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_238),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_173),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_173),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_151),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_67),
.C(n_109),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_29),
.A2(n_30),
.B1(n_109),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_30),
.B(n_154),
.Y(n_153)
);

AO21x2_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_41),
.B(n_55),
.Y(n_30)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_31),
.A2(n_41),
.B1(n_184),
.B2(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_31),
.B(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_31),
.A2(n_41),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_31),
.A2(n_41),
.B1(n_411),
.B2(n_494),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_31),
.A2(n_41),
.B1(n_494),
.B2(n_513),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_31),
.A2(n_41),
.B1(n_223),
.B2(n_513),
.Y(n_565)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AO21x2_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_42),
.B(n_47),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_36),
.Y(n_218)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_36),
.Y(n_473)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_38),
.Y(n_252)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_41),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_45),
.Y(n_319)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_45),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_46),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_46),
.Y(n_312)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_46),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_47),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_51),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_51),
.Y(n_353)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_55),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_56),
.B(n_264),
.Y(n_382)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_59),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_65),
.Y(n_228)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_65),
.Y(n_414)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_66),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_67),
.B(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_79),
.B1(n_102),
.B2(n_107),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_68),
.A2(n_79),
.B1(n_107),
.B2(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_74),
.Y(n_491)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_75),
.Y(n_489)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_79),
.A2(n_107),
.B1(n_530),
.B2(n_536),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_92),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_80)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_81),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_81),
.Y(n_553)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_82),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_82),
.Y(n_486)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_83),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_84),
.Y(n_535)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_87),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_91),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_98),
.Y(n_462)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_99),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_101),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_101),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_102),
.Y(n_172)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_R g438 ( 
.A(n_108),
.B(n_264),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_108),
.A2(n_171),
.B1(n_483),
.B2(n_487),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_108),
.A2(n_171),
.B1(n_548),
.B2(n_551),
.Y(n_547)
);

OAI22x1_ASAP7_75t_SL g579 ( 
.A1(n_108),
.A2(n_171),
.B1(n_548),
.B2(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_120),
.B1(n_143),
.B2(n_145),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_111),
.A2(n_144),
.B1(n_193),
.B2(n_199),
.Y(n_192)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_118),
.Y(n_402)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_120),
.A2(n_143),
.B1(n_145),
.B2(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_120),
.A2(n_143),
.B1(n_391),
.B2(n_396),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_120),
.A2(n_143),
.B1(n_396),
.B2(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_120),
.A2(n_143),
.B1(n_422),
.B2(n_498),
.Y(n_497)
);

OA22x2_ASAP7_75t_L g537 ( 
.A1(n_120),
.A2(n_143),
.B1(n_498),
.B2(n_538),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_120),
.A2(n_143),
.B1(n_538),
.B2(n_555),
.Y(n_554)
);

AO21x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_128),
.B(n_134),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_130),
.Y(n_393)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_130),
.Y(n_502)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_140),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_135),
.Y(n_496)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22x1_ASAP7_75t_L g581 ( 
.A1(n_144),
.A2(n_193),
.B1(n_199),
.B2(n_582),
.Y(n_581)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2x1_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_163),
.Y(n_152)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g381 ( 
.A(n_162),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_163)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_200),
.Y(n_173)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_174),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_177),
.B(n_200),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_178),
.A2(n_179),
.B(n_192),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_192),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_181),
.A2(n_182),
.B1(n_307),
.B2(n_317),
.Y(n_306)
);

NAND2x1_ASAP7_75t_SL g346 ( 
.A(n_181),
.B(n_347),
.Y(n_346)
);

AOI22x1_ASAP7_75t_L g385 ( 
.A1(n_181),
.A2(n_182),
.B1(n_347),
.B2(n_386),
.Y(n_385)
);

NAND2x1_ASAP7_75t_L g345 ( 
.A(n_182),
.B(n_307),
.Y(n_345)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_203),
.B(n_229),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g594 ( 
.A(n_202),
.B(n_595),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_222),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_203),
.A2(n_573),
.B1(n_574),
.B2(n_575),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_203),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_207),
.B(n_215),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_208),
.A2(n_250),
.B1(n_272),
.B2(n_281),
.Y(n_271)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_208),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_208),
.A2(n_323),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_208),
.A2(n_470),
.B1(n_519),
.B2(n_522),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_208),
.A2(n_257),
.B1(n_519),
.B2(n_564),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_211),
.Y(n_468)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx2_ASAP7_75t_SL g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_213),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_215),
.Y(n_564)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_222),
.Y(n_575)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx4f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g595 ( 
.A(n_229),
.B(n_573),
.Y(n_595)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_230),
.Y(n_580)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_606),
.B(n_613),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_505),
.B(n_601),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_442),
.B(n_504),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_404),
.B(n_441),
.Y(n_243)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_356),
.B(n_403),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_331),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_285),
.B(n_328),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_270),
.B(n_284),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_262),
.Y(n_248)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_261),
.Y(n_335)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_261),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_297),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_264),
.A2(n_296),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_266),
.A2(n_322),
.B1(n_326),
.B2(n_327),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_283),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_283),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_276),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_276),
.Y(n_436)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_321),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_305),
.B1(n_306),
.B2(n_320),
.Y(n_286)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g329 ( 
.A(n_287),
.B(n_305),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_295),
.B1(n_299),
.B2(n_304),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_305),
.B(n_320),
.Y(n_332)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_320),
.Y(n_330)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_329),
.B(n_330),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AO22x1_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_337),
.B1(n_364),
.B2(n_367),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_326),
.A2(n_367),
.B1(n_432),
.B2(n_434),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_326),
.A2(n_434),
.B1(n_466),
.B2(n_469),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_357),
.B(n_358),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_344),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_354),
.C(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B(n_354),
.C(n_355),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_346),
.C(n_354),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_R g360 ( 
.A(n_345),
.B(n_346),
.Y(n_360)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_350),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_353),
.Y(n_517)
);

NOR2x1_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_361),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_383),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_362),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_375),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_363),
.B(n_375),
.Y(n_408)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_SL g395 ( 
.A(n_380),
.Y(n_395)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_381),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_389),
.B2(n_390),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_389),
.C(n_440),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_387),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_397),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_399),
.Y(n_558)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_439),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_405),
.B(n_439),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_419),
.B2(n_420),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_417),
.B2(n_418),
.Y(n_407)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_408),
.Y(n_418)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_409),
.B(n_418),
.C(n_419),
.Y(n_503)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_430),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_421),
.B(n_438),
.C(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_426),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_429),
.Y(n_500)
);

XNOR2x1_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_438),
.Y(n_430)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_503),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_503),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_480),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_478),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_478),
.C(n_480),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_465),
.B1(n_476),
.B2(n_477),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_477),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_446),
.B(n_477),
.Y(n_561)
);

OAI32xp33_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_449),
.A3(n_452),
.B1(n_456),
.B2(n_463),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_SL g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

BUFx2_ASAP7_75t_SL g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_492),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_SL g510 ( 
.A(n_482),
.B(n_493),
.C(n_497),
.Y(n_510)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_SL g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_487),
.Y(n_536)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NAND4xp25_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_541),
.C(n_585),
.D(n_596),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_507),
.B(n_508),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_526),
.Y(n_508)
);

XNOR2x1_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_511),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_510),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_511),
.B(n_526),
.C(n_598),
.Y(n_597)
);

XOR2x2_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_518),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_512),
.B(n_518),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx3_ASAP7_75t_SL g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_528),
.Y(n_526)
);

XNOR2x1_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_537),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_529),
.B(n_537),
.C(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_535),
.Y(n_534)
);

A2O1A1O1Ixp25_ASAP7_75t_L g601 ( 
.A1(n_541),
.A2(n_585),
.B(n_602),
.C(n_604),
.D(n_605),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_566),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_542),
.B(n_566),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_560),
.C(n_562),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_562),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_546),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_568),
.C(n_570),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_554),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_547),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_554),
.Y(n_570)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_555),
.Y(n_582)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_560),
.B(n_600),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_565),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_563),
.B(n_565),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_571),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_567),
.B(n_572),
.C(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_576),
.Y(n_571)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_576),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_577),
.A2(n_578),
.B1(n_583),
.B2(n_584),
.Y(n_576)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_577),
.Y(n_584)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_578),
.Y(n_583)
);

XNOR2x1_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_581),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_579),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_581),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_584),
.B(n_590),
.C(n_591),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_586),
.B(n_588),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_588),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_592),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_589),
.B(n_608),
.C(n_609),
.Y(n_607)
);

XOR2x1_ASAP7_75t_L g592 ( 
.A(n_593),
.B(n_594),
.Y(n_592)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_593),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_594),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_597),
.B(n_599),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_597),
.B(n_599),
.C(n_603),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_610),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_607),
.B(n_610),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_612),
.Y(n_610)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);


endmodule