module fake_jpeg_31556_n_71 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_28;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_43;
wire n_29;
wire n_50;
wire n_37;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_21),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_29),
.B1(n_28),
.B2(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_25),
.A2(n_21),
.B1(n_34),
.B2(n_22),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_30),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_29),
.B1(n_36),
.B2(n_26),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_23),
.A2(n_35),
.B1(n_29),
.B2(n_28),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_47),
.B1(n_42),
.B2(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_51),
.A2(n_47),
.B(n_43),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_58),
.B1(n_52),
.B2(n_53),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_52),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_49),
.B(n_61),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_43),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_48),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_67),
.B1(n_49),
.B2(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_48),
.Y(n_71)
);


endmodule