module fake_jpeg_27732_n_22 (n_3, n_2, n_1, n_0, n_4, n_5, n_22);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_3),
.B(n_2),
.Y(n_6)
);

OAI21xp33_ASAP7_75t_L g7 ( 
.A1(n_1),
.A2(n_5),
.B(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_10),
.B(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_14),
.CI(n_9),
.CON(n_16),
.SN(n_16)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_5),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_13),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_15),
.B(n_18),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_16),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_17),
.C(n_16),
.Y(n_22)
);


endmodule