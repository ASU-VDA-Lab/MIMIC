module fake_jpeg_17850_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_33),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_18),
.B1(n_15),
.B2(n_20),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_13),
.B1(n_18),
.B2(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_42),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_15),
.B1(n_22),
.B2(n_23),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_25),
.B1(n_24),
.B2(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_23),
.B1(n_19),
.B2(n_14),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_21),
.Y(n_68)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_64),
.Y(n_76)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_29),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_67),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_68),
.B(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_67),
.C(n_64),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_35),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_50),
.B1(n_44),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_68),
.B1(n_55),
.B2(n_62),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_21),
.B(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_39),
.B1(n_13),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_82),
.B1(n_26),
.B2(n_66),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_26),
.B1(n_14),
.B2(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_89),
.B1(n_93),
.B2(n_84),
.C(n_81),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_68),
.B1(n_57),
.B2(n_53),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_59),
.B1(n_32),
.B2(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_95),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_76),
.C(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_32),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_47),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_78),
.C(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_104),
.B1(n_100),
.B2(n_103),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_81),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_74),
.B(n_73),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_96),
.B(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_35),
.C(n_70),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_35),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_86),
.B1(n_89),
.B2(n_88),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_97),
.B1(n_47),
.B2(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

OAI321xp33_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_107),
.A3(n_109),
.B1(n_4),
.B2(n_5),
.C(n_3),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_11),
.B(n_7),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_111),
.B(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_117),
.B1(n_118),
.B2(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_123),
.B1(n_127),
.B2(n_2),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_130),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_139),
.C(n_136),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_134),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.C(n_9),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_140),
.A2(n_137),
.B(n_123),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_10),
.C(n_12),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_12),
.Y(n_145)
);


endmodule