module fake_jpeg_29010_n_46 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_16),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_17),
.B1(n_9),
.B2(n_15),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_16),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_33),
.B(n_29),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_17),
.B1(n_11),
.B2(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_26),
.B1(n_20),
.B2(n_5),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_3),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_33),
.C(n_4),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_32),
.B(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.C(n_5),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_35),
.C(n_7),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_6),
.B(n_8),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_43),
.B(n_12),
.Y(n_46)
);


endmodule