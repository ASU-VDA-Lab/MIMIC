module fake_jpeg_27166_n_95 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_0),
.B(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_47),
.B1(n_6),
.B2(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_2),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_36),
.B1(n_34),
.B2(n_37),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_54),
.B1(n_32),
.B2(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_38),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_37),
.B1(n_33),
.B2(n_34),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_5),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_7),
.B(n_8),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_6),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_43),
.B1(n_18),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_77),
.B1(n_59),
.B2(n_58),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_69),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_16),
.C(n_31),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_68),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_75),
.B1(n_76),
.B2(n_26),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_9),
.B(n_10),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_15),
.Y(n_81)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_13),
.B(n_14),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_75),
.B(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_83),
.B1(n_66),
.B2(n_64),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_84),
.C(n_79),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.B(n_65),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_84),
.B1(n_86),
.B2(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_78),
.B1(n_74),
.B2(n_71),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_60),
.B(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_72),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_80),
.Y(n_95)
);


endmodule