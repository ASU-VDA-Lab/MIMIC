module fake_netlist_5_146_n_1676 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1676);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1676;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_26),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_24),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_20),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_65),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_78),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_48),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_50),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_29),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_44),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_38),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_87),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_38),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_56),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_92),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_68),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_82),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_53),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_11),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_36),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_41),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_24),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_104),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_13),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_4),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_52),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_19),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_37),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_58),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_7),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_110),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_60),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_70),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_77),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_46),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_59),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_141),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_39),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_64),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_97),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_74),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_34),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_117),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_6),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_55),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_116),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_103),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_39),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_96),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_8),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_16),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_83),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_34),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_3),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_27),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_69),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_18),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_108),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_0),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_12),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_79),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_101),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_15),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_36),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_113),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_23),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_95),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_54),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_3),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_5),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_106),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_66),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_122),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_91),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_89),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_146),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_43),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_128),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_154),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_144),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_35),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_47),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_76),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_119),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_73),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_17),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_80),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_61),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_98),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_12),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_10),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_86),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_88),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_111),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_142),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_16),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_41),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_140),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_30),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_14),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_132),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_130),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_51),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_256),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_188),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_196),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_203),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_206),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_208),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_157),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_158),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_158),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

BUFx2_ASAP7_75t_SL g322 ( 
.A(n_160),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_155),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_178),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_211),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_190),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_212),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_214),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_197),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_182),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_216),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_218),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_234),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_241),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_204),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_246),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_155),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_156),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_221),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_170),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_226),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_229),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_170),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_171),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_171),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_268),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_172),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_157),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_198),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_163),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_172),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_191),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_163),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_174),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_159),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_175),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_161),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_157),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_165),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_169),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_263),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_175),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_166),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_168),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_177),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_186),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_184),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_187),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_263),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_186),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_189),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_160),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_310),
.A2(n_245),
.B1(n_244),
.B2(n_236),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_371),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

CKINVDCx11_ASAP7_75t_R g390 ( 
.A(n_308),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_257),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_257),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_314),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_309),
.B(n_274),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_340),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_332),
.A2(n_230),
.B1(n_292),
.B2(n_299),
.Y(n_401)
);

BUFx12f_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_199),
.B(n_169),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_274),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_340),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_326),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_361),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_164),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_356),
.A2(n_248),
.B1(n_247),
.B2(n_276),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_164),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_374),
.B(n_199),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_167),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_328),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_322),
.B(n_173),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_322),
.B(n_270),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_311),
.B(n_213),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_377),
.B(n_167),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_321),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_362),
.B(n_213),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_331),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_338),
.A2(n_262),
.B1(n_261),
.B2(n_286),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_325),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_368),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_382),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_312),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_379),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_337),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_346),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_313),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_313),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_364),
.B(n_237),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_315),
.B(n_192),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_359),
.B(n_318),
.Y(n_451)
);

NOR2x1p5_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_347),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_402),
.B(n_342),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_418),
.A2(n_323),
.B1(n_376),
.B2(n_366),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_445),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_409),
.Y(n_458)
);

AND3x2_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_253),
.C(n_237),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_418),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_442),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_387),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_390),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_449),
.B(n_315),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_442),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_388),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_316),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_389),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_449),
.B(n_316),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_390),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_440),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_402),
.B(n_319),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_327),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_437),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_437),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_436),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_389),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_434),
.Y(n_489)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_405),
.A2(n_278),
.B(n_253),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_445),
.B(n_327),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_434),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_451),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_423),
.B(n_329),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g499 ( 
.A(n_385),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_410),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_441),
.B(n_329),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_411),
.A2(n_194),
.B(n_193),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_424),
.B(n_330),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_447),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_441),
.B(n_330),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_441),
.B(n_341),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_440),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_444),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_441),
.B(n_333),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_448),
.B(n_333),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_444),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_410),
.Y(n_519)
);

AND3x2_ASAP7_75t_L g520 ( 
.A(n_431),
.B(n_295),
.C(n_278),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_418),
.B(n_334),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_450),
.B(n_343),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_428),
.B(n_263),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_448),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_410),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_439),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_411),
.B(n_334),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_401),
.A2(n_249),
.B1(n_267),
.B2(n_282),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_448),
.B(n_335),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_418),
.B(n_335),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_444),
.Y(n_531)
);

INVxp33_ASAP7_75t_SL g532 ( 
.A(n_385),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_428),
.B(n_336),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_263),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_448),
.B(n_336),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_440),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

AO21x2_ASAP7_75t_L g539 ( 
.A1(n_415),
.A2(n_200),
.B(n_195),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_408),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_440),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_410),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_414),
.B(n_349),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_383),
.B(n_295),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_414),
.B(n_349),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_440),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_415),
.B(n_351),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_419),
.B(n_351),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_419),
.B(n_372),
.C(n_360),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_410),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_421),
.Y(n_551)
);

NOR2x1p5_ASAP7_75t_L g552 ( 
.A(n_426),
.B(n_360),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_396),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_400),
.B(n_162),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_440),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_421),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_396),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_450),
.B(n_344),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_396),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_443),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_450),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_400),
.B(n_305),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_426),
.B(n_372),
.Y(n_563)
);

INVx8_ASAP7_75t_L g564 ( 
.A(n_396),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_400),
.B(n_202),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_396),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_421),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_383),
.A2(n_323),
.B1(n_339),
.B2(n_357),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_427),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_427),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_400),
.B(n_209),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_R g574 ( 
.A(n_439),
.B(n_381),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_433),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_412),
.Y(n_577)
);

AND3x2_ASAP7_75t_L g578 ( 
.A(n_383),
.B(n_353),
.C(n_317),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_443),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_400),
.B(n_215),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_432),
.A2(n_381),
.B1(n_306),
.B2(n_302),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_435),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_R g583 ( 
.A(n_446),
.B(n_219),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_407),
.B(n_220),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_435),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_384),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_412),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_399),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_432),
.B(n_180),
.Y(n_591)
);

AND2x2_ASAP7_75t_SL g592 ( 
.A(n_399),
.B(n_263),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_384),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_420),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_420),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_392),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_422),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_422),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_429),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_413),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_461),
.B(n_407),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_456),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_524),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_592),
.A2(n_539),
.B1(n_503),
.B2(n_532),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_547),
.A2(n_176),
.B1(n_399),
.B2(n_446),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_592),
.B(n_407),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_524),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_521),
.A2(n_265),
.B1(n_223),
.B2(n_217),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_565),
.A2(n_407),
.B(n_416),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_484),
.B(n_401),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_552),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_425),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_425),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_504),
.B(n_391),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_533),
.B(n_391),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_522),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_527),
.B(n_425),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_589),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_548),
.B(n_413),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_563),
.B(n_413),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_554),
.B(n_417),
.Y(n_623)
);

AO221x1_ASAP7_75t_L g624 ( 
.A1(n_494),
.A2(n_227),
.B1(n_232),
.B2(n_235),
.C(n_239),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_562),
.B(n_417),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_471),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_530),
.B(n_417),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_557),
.B(n_201),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_589),
.B(n_397),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_594),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_594),
.B(n_397),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_597),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_557),
.B(n_205),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_597),
.B(n_397),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_557),
.B(n_210),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_471),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_479),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_598),
.B(n_397),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_495),
.B(n_406),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_598),
.B(n_403),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_599),
.B(n_403),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_457),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_516),
.A2(n_222),
.B1(n_224),
.B2(n_242),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_599),
.B(n_403),
.Y(n_645)
);

NOR2x1p5_ASAP7_75t_L g646 ( 
.A(n_549),
.B(n_247),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_480),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_557),
.B(n_243),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_508),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_457),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_522),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_454),
.A2(n_251),
.B1(n_260),
.B2(n_264),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_557),
.B(n_271),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_508),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_513),
.B(n_529),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_SL g657 ( 
.A(n_577),
.B(n_499),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_566),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_538),
.B(n_403),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_540),
.B(n_398),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_479),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_566),
.B(n_398),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_503),
.A2(n_301),
.B1(n_277),
.B2(n_281),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_600),
.B(n_386),
.Y(n_664)
);

NOR3xp33_ASAP7_75t_L g665 ( 
.A(n_591),
.B(n_406),
.C(n_348),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_503),
.A2(n_539),
.B1(n_532),
.B2(n_544),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_462),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_559),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_458),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_539),
.A2(n_273),
.B1(n_297),
.B2(n_288),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_544),
.A2(n_283),
.B1(n_307),
.B2(n_429),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_513),
.B(n_535),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_464),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_491),
.B(n_430),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_544),
.A2(n_438),
.B1(n_430),
.B2(n_404),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_600),
.B(n_386),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_513),
.B(n_180),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_600),
.B(n_559),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_523),
.A2(n_438),
.B(n_404),
.C(n_352),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_465),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_559),
.B(n_416),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_559),
.B(n_416),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_472),
.B(n_416),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_588),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_522),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_588),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_593),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_510),
.B(n_354),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_595),
.B(n_416),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_561),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_506),
.B(n_392),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_596),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_458),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_502),
.B(n_394),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_543),
.B(n_183),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_574),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_507),
.B(n_394),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_596),
.Y(n_698)
);

INVx8_ASAP7_75t_L g699 ( 
.A(n_577),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_515),
.A2(n_225),
.B1(n_228),
.B2(n_231),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_526),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_595),
.B(n_553),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_595),
.B(n_233),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_544),
.A2(n_276),
.B1(n_248),
.B2(n_275),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_455),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_455),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_465),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_522),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_460),
.B(n_395),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_470),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_558),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_564),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_460),
.B(n_395),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_564),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_491),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_463),
.B(n_238),
.Y(n_716)
);

BUFx8_ASAP7_75t_L g717 ( 
.A(n_577),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_558),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_523),
.A2(n_534),
.B(n_501),
.C(n_545),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_501),
.Y(n_720)
);

BUFx5_ASAP7_75t_L g721 ( 
.A(n_463),
.Y(n_721)
);

OAI221xp5_ASAP7_75t_L g722 ( 
.A1(n_528),
.A2(n_568),
.B1(n_581),
.B2(n_517),
.C(n_486),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_553),
.B(n_240),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_468),
.B(n_183),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_468),
.B(n_469),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_544),
.A2(n_534),
.B1(n_486),
.B2(n_514),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_506),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_469),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_558),
.B(n_355),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_572),
.B(n_185),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_580),
.B(n_185),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_553),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_476),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_476),
.A2(n_255),
.B1(n_286),
.B2(n_266),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_510),
.A2(n_279),
.B1(n_269),
.B2(n_306),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_485),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_467),
.B(n_269),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_584),
.B(n_293),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_514),
.A2(n_255),
.B1(n_275),
.B2(n_304),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_531),
.B(n_285),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_531),
.B(n_285),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_564),
.B(n_289),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_473),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_473),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_564),
.B(n_289),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_560),
.B(n_272),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_558),
.Y(n_747)
);

INVxp33_ASAP7_75t_L g748 ( 
.A(n_583),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_560),
.B(n_272),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_579),
.B(n_290),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_579),
.B(n_290),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_586),
.B(n_279),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_466),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_478),
.B(n_298),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_510),
.A2(n_293),
.B1(n_298),
.B2(n_302),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_586),
.B(n_500),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_492),
.B(n_436),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_500),
.B(n_179),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_705),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_706),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_728),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_606),
.A2(n_510),
.B1(n_483),
.B2(n_541),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_616),
.B(n_587),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_647),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_648),
.B(n_483),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_619),
.B(n_453),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_606),
.A2(n_483),
.B1(n_541),
.B2(n_555),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_650),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_616),
.B(n_587),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_715),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_612),
.A2(n_546),
.B(n_537),
.C(n_474),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_712),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_658),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_612),
.B(n_483),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_604),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_715),
.B(n_585),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_638),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_655),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_601),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_661),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_720),
.B(n_585),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_712),
.B(n_555),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_617),
.A2(n_303),
.B1(n_266),
.B2(n_262),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_720),
.B(n_582),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_640),
.B(n_578),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_551),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_684),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_656),
.B(n_487),
.Y(n_788)
);

AND3x1_ASAP7_75t_SL g789 ( 
.A(n_646),
.B(n_452),
.C(n_722),
.Y(n_789)
);

BUFx4f_ASAP7_75t_L g790 ( 
.A(n_699),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_622),
.B(n_551),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_729),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_686),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_687),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_602),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_605),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_640),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_656),
.B(n_482),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_732),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_658),
.B(n_459),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_727),
.Y(n_801)
);

O2A1O1Ixp5_ASAP7_75t_L g802 ( 
.A1(n_627),
.A2(n_490),
.B(n_474),
.C(n_575),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_620),
.B(n_630),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_609),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_669),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_695),
.A2(n_546),
.B(n_537),
.C(n_525),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_692),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_693),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_698),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_672),
.A2(n_505),
.B1(n_498),
.B2(n_511),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_743),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_672),
.B(n_520),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_744),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_688),
.B(n_358),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_696),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_632),
.Y(n_816)
);

INVx5_ASAP7_75t_L g817 ( 
.A(n_712),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_526),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_613),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_717),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_688),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_674),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_717),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_695),
.B(n_254),
.C(n_261),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_SL g825 ( 
.A(n_701),
.B(n_753),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_733),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_R g827 ( 
.A(n_657),
.B(n_466),
.Y(n_827)
);

AND2x6_ASAP7_75t_SL g828 ( 
.A(n_757),
.B(n_481),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_618),
.B(n_498),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_677),
.B(n_481),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_663),
.A2(n_582),
.B1(n_576),
.B2(n_575),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_736),
.Y(n_832)
);

OR2x6_ASAP7_75t_L g833 ( 
.A(n_699),
.B(n_556),
.Y(n_833)
);

INVx5_ASAP7_75t_L g834 ( 
.A(n_712),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_643),
.Y(n_835)
);

AND2x6_ASAP7_75t_SL g836 ( 
.A(n_737),
.B(n_249),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_652),
.B(n_498),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_690),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_651),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_614),
.B(n_556),
.Y(n_840)
);

OR2x2_ASAP7_75t_SL g841 ( 
.A(n_615),
.B(n_249),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_691),
.B(n_482),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_694),
.B(n_567),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_699),
.B(n_567),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_697),
.B(n_576),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_708),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_603),
.B(n_721),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_667),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_737),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_675),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_665),
.B(n_254),
.C(n_304),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_663),
.A2(n_573),
.B1(n_571),
.B2(n_570),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_662),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_711),
.B(n_505),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_718),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_SL g857 ( 
.A(n_748),
.B(n_179),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_747),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_675),
.B(n_482),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_751),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_607),
.B(n_303),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_725),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_603),
.B(n_573),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_660),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_713),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_754),
.Y(n_867)
);

AND2x2_ASAP7_75t_SL g868 ( 
.A(n_666),
.B(n_670),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_714),
.Y(n_869)
);

BUFx4f_ASAP7_75t_L g870 ( 
.A(n_674),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_754),
.B(n_571),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_703),
.B(n_570),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_668),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_674),
.Y(n_874)
);

NOR2x1p5_ASAP7_75t_L g875 ( 
.A(n_730),
.B(n_282),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_751),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_674),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_732),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_721),
.B(n_569),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_673),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_721),
.B(n_569),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_740),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_724),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_721),
.B(n_497),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_721),
.B(n_497),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_702),
.B(n_505),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_703),
.B(n_489),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_674),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_680),
.Y(n_889)
);

AND2x2_ASAP7_75t_SL g890 ( 
.A(n_666),
.B(n_670),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_707),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_721),
.B(n_496),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_710),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_758),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_700),
.B(n_550),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_734),
.B(n_739),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_702),
.B(n_489),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_756),
.Y(n_898)
);

OR2x2_ASAP7_75t_SL g899 ( 
.A(n_731),
.B(n_738),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_758),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_726),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_608),
.A2(n_550),
.B(n_542),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_608),
.B(n_496),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_741),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_723),
.B(n_542),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_653),
.A2(n_704),
.B1(n_624),
.B2(n_671),
.Y(n_906)
);

INVx3_ASAP7_75t_SL g907 ( 
.A(n_723),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_756),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_704),
.B(n_512),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_746),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_626),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_629),
.B(n_493),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_634),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_734),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_637),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_678),
.B(n_536),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_742),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_745),
.Y(n_918)
);

AND2x2_ASAP7_75t_SL g919 ( 
.A(n_671),
.B(n_726),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_749),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_735),
.B(n_536),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_659),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_628),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_631),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_635),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_639),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_641),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_642),
.B(n_493),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_689),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_645),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_679),
.Y(n_931)
);

AND3x1_ASAP7_75t_L g932 ( 
.A(n_739),
.B(n_267),
.C(n_282),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_623),
.B(n_519),
.Y(n_933)
);

AOI22x1_ASAP7_75t_L g934 ( 
.A1(n_611),
.A2(n_519),
.B1(n_518),
.B2(n_477),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_681),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_755),
.B(n_512),
.Y(n_936)
);

AO22x1_ASAP7_75t_L g937 ( 
.A1(n_850),
.A2(n_610),
.B1(n_750),
.B2(n_752),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_759),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_774),
.A2(n_719),
.B(n_683),
.C(n_636),
.Y(n_939)
);

INVx8_ASAP7_75t_L g940 ( 
.A(n_817),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_797),
.B(n_689),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_851),
.A2(n_682),
.B(n_676),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_816),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_817),
.B(n_628),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_826),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_786),
.A2(n_664),
.B(n_625),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_797),
.B(n_716),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_867),
.B(n_644),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_791),
.A2(n_654),
.B(n_649),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_775),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_832),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_780),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_SL g953 ( 
.A(n_824),
.B(n_654),
.C(n_649),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_777),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_838),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_770),
.B(n_636),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_792),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_869),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_791),
.A2(n_633),
.B(n_512),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_811),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_879),
.A2(n_512),
.B(n_488),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_815),
.B(n_490),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_862),
.B(n_865),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_866),
.B(n_475),
.Y(n_964)
);

AND3x1_ASAP7_75t_SL g965 ( 
.A(n_875),
.B(n_267),
.C(n_284),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_SL g966 ( 
.A(n_824),
.B(n_284),
.C(n_207),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_801),
.B(n_284),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_868),
.A2(n_890),
.B1(n_914),
.B2(n_896),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_805),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_881),
.A2(n_848),
.B(n_884),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_868),
.A2(n_890),
.B1(n_919),
.B2(n_901),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_910),
.B(n_207),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_SL g973 ( 
.A1(n_932),
.A2(n_207),
.B1(n_179),
.B2(n_10),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_817),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_766),
.A2(n_910),
.B(n_861),
.C(n_900),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_854),
.B(n_901),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_798),
.A2(n_139),
.B(n_137),
.C(n_134),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_861),
.A2(n_2),
.B1(n_9),
.B2(n_14),
.C(n_15),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_881),
.A2(n_131),
.B(n_129),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_835),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_848),
.A2(n_127),
.B(n_126),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_900),
.A2(n_9),
.B(n_17),
.C(n_18),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_884),
.A2(n_125),
.B(n_112),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_869),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_919),
.B(n_93),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_821),
.B(n_84),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_814),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_808),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_819),
.B(n_85),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_883),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_920),
.B(n_75),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_SL g992 ( 
.A1(n_771),
.A2(n_72),
.B(n_49),
.C(n_45),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_929),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_864),
.B(n_22),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_860),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_839),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_800),
.B(n_25),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_902),
.A2(n_28),
.B(n_29),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_929),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_999)
);

OAI33xp33_ASAP7_75t_L g1000 ( 
.A1(n_783),
.A2(n_31),
.A3(n_32),
.B1(n_33),
.B2(n_37),
.B3(n_40),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_818),
.B(n_33),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_885),
.A2(n_40),
.B(n_42),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_790),
.B(n_42),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_849),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_882),
.B(n_904),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_925),
.B(n_43),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_760),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_R g1008 ( 
.A(n_790),
.B(n_825),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_926),
.B(n_927),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_830),
.B(n_814),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_869),
.B(n_823),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_761),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_800),
.B(n_765),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_858),
.Y(n_1014)
);

CKINVDCx6p67_ASAP7_75t_R g1015 ( 
.A(n_820),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_828),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_921),
.A2(n_906),
.B1(n_876),
.B2(n_918),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_833),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_785),
.A2(n_783),
.B(n_907),
.C(n_788),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_785),
.A2(n_789),
.B1(n_894),
.B2(n_918),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_802),
.A2(n_902),
.B(n_806),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_924),
.B(n_922),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_907),
.B(n_857),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_917),
.B(n_918),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_899),
.B(n_812),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_873),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_847),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_906),
.A2(n_769),
.B1(n_763),
.B2(n_803),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_763),
.A2(n_769),
.B1(n_877),
.B2(n_871),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_845),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_SL g1031 ( 
.A(n_812),
.B(n_852),
.C(n_827),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_803),
.B(n_871),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_917),
.B(n_773),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_930),
.B(n_935),
.Y(n_1034)
);

OAI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_779),
.A2(n_795),
.B1(n_804),
.B2(n_796),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_765),
.B(n_762),
.C(n_773),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_892),
.A2(n_933),
.B(n_859),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_873),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_789),
.A2(n_917),
.B1(n_921),
.B2(n_936),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_817),
.A2(n_834),
.B(n_781),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_764),
.B(n_768),
.Y(n_1041)
);

INVx5_ASAP7_75t_L g1042 ( 
.A(n_834),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_877),
.A2(n_799),
.B1(n_870),
.B2(n_936),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_L g1044 ( 
.A(n_833),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_877),
.A2(n_799),
.B1(n_870),
.B2(n_843),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_778),
.B(n_856),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_843),
.B(n_846),
.Y(n_1047)
);

AO22x1_ASAP7_75t_L g1048 ( 
.A1(n_829),
.A2(n_855),
.B1(n_837),
.B2(n_886),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_834),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_889),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_802),
.A2(n_909),
.B(n_903),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_923),
.B(n_793),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_834),
.B(n_923),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_787),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_776),
.A2(n_784),
.B(n_781),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_923),
.B(n_878),
.Y(n_1056)
);

INVx6_ASAP7_75t_L g1057 ( 
.A(n_833),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_767),
.A2(n_794),
.B(n_809),
.C(n_807),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_846),
.B(n_840),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_776),
.A2(n_784),
.B1(n_853),
.B2(n_831),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_912),
.A2(n_928),
.B(n_840),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_842),
.B(n_872),
.C(n_887),
.Y(n_1062)
);

CKINVDCx16_ASAP7_75t_R g1063 ( 
.A(n_827),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_813),
.A2(n_931),
.B(n_872),
.C(n_887),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_878),
.B(n_888),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_905),
.A2(n_898),
.B1(n_908),
.B2(n_886),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_897),
.A2(n_905),
.B(n_895),
.C(n_874),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_880),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_897),
.A2(n_822),
.B(n_874),
.C(n_913),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_829),
.B(n_855),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_844),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_772),
.B(n_844),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_822),
.A2(n_915),
.B(n_911),
.C(n_893),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_916),
.B(n_837),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_836),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_891),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_990),
.B(n_841),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_939),
.A2(n_863),
.B(n_853),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_1042),
.B(n_772),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1055),
.A2(n_1061),
.B(n_946),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_969),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_SL g1082 ( 
.A1(n_1060),
.A2(n_888),
.B(n_782),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_978),
.B(n_810),
.C(n_831),
.Y(n_1083)
);

AOI21x1_ASAP7_75t_SL g1084 ( 
.A1(n_1006),
.A2(n_941),
.B(n_994),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_958),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_963),
.B(n_916),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_988),
.Y(n_1087)
);

CKINVDCx11_ASAP7_75t_R g1088 ( 
.A(n_1015),
.Y(n_1088)
);

AOI221xp5_ASAP7_75t_SL g1089 ( 
.A1(n_971),
.A2(n_1028),
.B1(n_982),
.B2(n_968),
.C(n_999),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_943),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_990),
.B(n_1001),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1013),
.B(n_1070),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1032),
.B(n_1009),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1022),
.B(n_976),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_947),
.B(n_1047),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_937),
.A2(n_948),
.B(n_1025),
.C(n_1028),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_955),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_945),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1059),
.B(n_975),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_951),
.Y(n_1100)
);

BUFx5_ASAP7_75t_L g1101 ( 
.A(n_1026),
.Y(n_1101)
);

AO31x2_ASAP7_75t_L g1102 ( 
.A1(n_1069),
.A2(n_971),
.A3(n_1060),
.B(n_1067),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1037),
.A2(n_1029),
.B(n_949),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_1021),
.A2(n_1051),
.B(n_998),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1063),
.Y(n_1105)
);

AOI221xp5_ASAP7_75t_L g1106 ( 
.A1(n_973),
.A2(n_1019),
.B1(n_1023),
.B2(n_1000),
.C(n_993),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_R g1107 ( 
.A(n_1030),
.B(n_1016),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1021),
.A2(n_1051),
.B(n_970),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_R g1109 ( 
.A1(n_1075),
.A2(n_1003),
.B1(n_966),
.B2(n_965),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1017),
.A2(n_1039),
.B1(n_1020),
.B2(n_1066),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1041),
.B(n_1052),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1073),
.A2(n_1045),
.A3(n_959),
.B(n_1043),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1007),
.Y(n_1113)
);

AO21x1_ASAP7_75t_L g1114 ( 
.A1(n_985),
.A2(n_1064),
.B(n_1062),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_953),
.A2(n_1058),
.B(n_985),
.C(n_1036),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1012),
.B(n_938),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_956),
.A2(n_1054),
.B1(n_1044),
.B2(n_1034),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1005),
.B(n_1038),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1068),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_1003),
.B(n_974),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_SL g1121 ( 
.A1(n_974),
.A2(n_1049),
.B(n_1040),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_1011),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1008),
.Y(n_1123)
);

AOI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1056),
.A2(n_1048),
.B(n_1065),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_995),
.A2(n_1002),
.A3(n_981),
.B(n_979),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_960),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_L g1127 ( 
.A(n_1031),
.B(n_972),
.C(n_991),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1042),
.A2(n_1049),
.B(n_940),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1024),
.B(n_1046),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_977),
.A2(n_983),
.B(n_964),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1076),
.A2(n_1074),
.A3(n_1050),
.B(n_980),
.Y(n_1131)
);

AO32x2_ASAP7_75t_L g1132 ( 
.A1(n_987),
.A2(n_992),
.A3(n_1027),
.B1(n_962),
.B2(n_1035),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_1053),
.A2(n_1033),
.B(n_1044),
.C(n_986),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_955),
.B(n_952),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_958),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_940),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_940),
.A2(n_944),
.B(n_1072),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_996),
.A2(n_1004),
.B(n_1014),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_958),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1013),
.B(n_986),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_957),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_954),
.A2(n_967),
.A3(n_1057),
.B(n_1071),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_989),
.A2(n_984),
.B(n_1018),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_950),
.B(n_997),
.Y(n_1144)
);

AO21x1_ASAP7_75t_L g1145 ( 
.A1(n_997),
.A2(n_967),
.B(n_1057),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1018),
.A2(n_1071),
.B(n_984),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_967),
.A2(n_939),
.B(n_1061),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_942),
.A2(n_934),
.B(n_961),
.Y(n_1148)
);

INVx3_ASAP7_75t_SL g1149 ( 
.A(n_1015),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_943),
.Y(n_1150)
);

AND3x4_ASAP7_75t_L g1151 ( 
.A(n_1013),
.B(n_808),
.C(n_805),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_942),
.A2(n_934),
.B(n_961),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_939),
.A2(n_1061),
.B(n_1037),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_963),
.B(n_797),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_963),
.B(n_797),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_943),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_952),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_963),
.B(n_797),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_940),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_963),
.B(n_797),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1032),
.A2(n_850),
.B1(n_867),
.B2(n_868),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_963),
.B(n_797),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_975),
.A2(n_612),
.B(n_766),
.C(n_824),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_955),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_942),
.A2(n_934),
.B(n_961),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_963),
.B(n_797),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_R g1167 ( 
.A(n_1063),
.B(n_669),
.Y(n_1167)
);

INVxp67_ASAP7_75t_SL g1168 ( 
.A(n_1032),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_943),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_939),
.A2(n_1061),
.B(n_1037),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_942),
.A2(n_934),
.B(n_961),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_990),
.B(n_456),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_939),
.A2(n_806),
.A3(n_771),
.B(n_1069),
.Y(n_1173)
);

AOI221x1_ASAP7_75t_L g1174 ( 
.A1(n_1062),
.A2(n_1028),
.B1(n_939),
.B2(n_1036),
.C(n_774),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_939),
.A2(n_806),
.A3(n_771),
.B(n_1069),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_942),
.A2(n_934),
.B(n_961),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_SL g1177 ( 
.A(n_985),
.B(n_868),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1015),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1032),
.A2(n_850),
.B1(n_867),
.B2(n_868),
.Y(n_1179)
);

CKINVDCx11_ASAP7_75t_R g1180 ( 
.A(n_1015),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1015),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_969),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_975),
.A2(n_612),
.B(n_766),
.C(n_824),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_971),
.A2(n_896),
.B1(n_824),
.B2(n_993),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_963),
.B(n_797),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_990),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_963),
.B(n_797),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_942),
.A2(n_934),
.B(n_961),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_SL g1189 ( 
.A1(n_978),
.A2(n_653),
.B1(n_896),
.B2(n_612),
.C(n_971),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_SL g1190 ( 
.A1(n_1067),
.A2(n_1069),
.B(n_941),
.C(n_991),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_975),
.A2(n_612),
.B(n_766),
.C(n_824),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_939),
.A2(n_806),
.A3(n_771),
.B(n_1069),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_SL g1193 ( 
.A1(n_976),
.A2(n_1058),
.B(n_1039),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_952),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1013),
.B(n_1070),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_990),
.B(n_456),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1055),
.A2(n_851),
.B(n_1061),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_963),
.B(n_797),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1021),
.A2(n_1051),
.B(n_998),
.Y(n_1199)
);

NAND2x1_ASAP7_75t_L g1200 ( 
.A(n_974),
.B(n_1049),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1010),
.B(n_990),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_963),
.B(n_797),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_L g1203 ( 
.A(n_978),
.B(n_612),
.C(n_850),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1152),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1171),
.A2(n_1188),
.B(n_1176),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1081),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1172),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1167),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1091),
.B(n_1201),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1174),
.A2(n_1114),
.A3(n_1080),
.B(n_1197),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1182),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1177),
.A2(n_1203),
.B1(n_1120),
.B2(n_1111),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1196),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1177),
.A2(n_1203),
.B1(n_1120),
.B2(n_1161),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1088),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1106),
.A2(n_1095),
.B(n_1093),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1153),
.A2(n_1170),
.B(n_1147),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1100),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1179),
.A2(n_1184),
.B1(n_1083),
.B2(n_1110),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1150),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1103),
.A2(n_1084),
.B(n_1078),
.Y(n_1221)
);

AND2x4_ASAP7_75t_SL g1222 ( 
.A(n_1122),
.B(n_1159),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1131),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_SL g1224 ( 
.A1(n_1193),
.A2(n_1145),
.B(n_1124),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1186),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1163),
.B(n_1191),
.C(n_1183),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1096),
.A2(n_1115),
.B(n_1099),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1103),
.A2(n_1078),
.B(n_1104),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1168),
.B(n_1154),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1090),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1155),
.B(n_1158),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1184),
.A2(n_1083),
.B1(n_1127),
.B2(n_1109),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1089),
.A2(n_1189),
.B(n_1094),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1199),
.A2(n_1108),
.B(n_1137),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1180),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1202),
.A2(n_1166),
.B1(n_1198),
.B2(n_1185),
.Y(n_1236)
);

BUFx2_ASAP7_75t_SL g1237 ( 
.A(n_1087),
.Y(n_1237)
);

AOI221xp5_ASAP7_75t_L g1238 ( 
.A1(n_1189),
.A2(n_1089),
.B1(n_1187),
.B2(n_1160),
.C(n_1162),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1097),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1131),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1117),
.A2(n_1132),
.A3(n_1108),
.B(n_1119),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_SL g1242 ( 
.A1(n_1151),
.A2(n_1123),
.B1(n_1077),
.B2(n_1105),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1133),
.A2(n_1190),
.B(n_1129),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1086),
.A2(n_1164),
.B1(n_1126),
.B2(n_1138),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1082),
.A2(n_1130),
.B(n_1121),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1136),
.Y(n_1246)
);

NOR3xp33_ASAP7_75t_SL g1247 ( 
.A(n_1178),
.B(n_1181),
.C(n_1144),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1113),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1156),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1130),
.A2(n_1128),
.B(n_1146),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1143),
.A2(n_1200),
.B(n_1116),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1157),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1085),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1169),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1092),
.B(n_1195),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1194),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1140),
.A2(n_1079),
.B(n_1139),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1134),
.B(n_1118),
.C(n_1141),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1131),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1092),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1173),
.A2(n_1192),
.B(n_1175),
.Y(n_1261)
);

NAND2x1p5_ASAP7_75t_L g1262 ( 
.A(n_1135),
.B(n_1101),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1132),
.A2(n_1192),
.B(n_1175),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1142),
.B(n_1135),
.Y(n_1264)
);

BUFx4f_ASAP7_75t_L g1265 ( 
.A(n_1149),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1101),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1142),
.B(n_1102),
.Y(n_1267)
);

INVx6_ASAP7_75t_L g1268 ( 
.A(n_1142),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1102),
.B(n_1125),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1102),
.B(n_1125),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1132),
.A2(n_1125),
.B1(n_1112),
.B2(n_1173),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1173),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1175),
.A2(n_1192),
.B(n_1112),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1112),
.B(n_1107),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1107),
.A2(n_850),
.B1(n_867),
.B2(n_1203),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_SL g1276 ( 
.A(n_1203),
.B(n_727),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1095),
.B(n_1093),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_SL g1278 ( 
.A1(n_1115),
.A2(n_982),
.B(n_995),
.C(n_1067),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1140),
.B(n_1039),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1131),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1091),
.B(n_1201),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1152),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1098),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1177),
.A2(n_850),
.B1(n_867),
.B2(n_532),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1203),
.A2(n_850),
.B1(n_867),
.B2(n_1111),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1152),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1177),
.A2(n_850),
.B1(n_867),
.B2(n_532),
.Y(n_1287)
);

AO21x1_ASAP7_75t_L g1288 ( 
.A1(n_1177),
.A2(n_1183),
.B(n_1163),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1140),
.B(n_1039),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1203),
.A2(n_978),
.B1(n_612),
.B2(n_973),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1088),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1203),
.A2(n_978),
.B1(n_612),
.B2(n_973),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1152),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1174),
.A2(n_1170),
.B(n_1153),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_R g1295 ( 
.A(n_1159),
.B(n_402),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1172),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1203),
.A2(n_978),
.B1(n_612),
.B2(n_973),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1098),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1095),
.B(n_1093),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1161),
.B(n_1179),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1174),
.A2(n_1170),
.B(n_1153),
.Y(n_1301)
);

AOI221x1_ASAP7_75t_L g1302 ( 
.A1(n_1203),
.A2(n_1115),
.B1(n_1147),
.B2(n_1184),
.C(n_1179),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1203),
.A2(n_850),
.B1(n_867),
.B2(n_1111),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1095),
.B(n_1093),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1131),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1081),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1098),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1082),
.B(n_1137),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1157),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1152),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1252),
.Y(n_1312)
);

OAI211xp5_ASAP7_75t_L g1313 ( 
.A1(n_1290),
.A2(n_1297),
.B(n_1292),
.C(n_1232),
.Y(n_1313)
);

O2A1O1Ixp5_ASAP7_75t_L g1314 ( 
.A1(n_1288),
.A2(n_1227),
.B(n_1300),
.C(n_1226),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_SL g1315 ( 
.A1(n_1274),
.A2(n_1270),
.B(n_1269),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1223),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1209),
.B(n_1281),
.Y(n_1317)
);

OAI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1285),
.A2(n_1303),
.B1(n_1302),
.B2(n_1212),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1290),
.A2(n_1292),
.B(n_1297),
.C(n_1300),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1236),
.B(n_1277),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1231),
.B(n_1232),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_SL g1322 ( 
.A1(n_1264),
.A2(n_1267),
.B(n_1305),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1255),
.B(n_1225),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1219),
.A2(n_1243),
.B(n_1216),
.C(n_1214),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1299),
.B(n_1304),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1284),
.A2(n_1287),
.B1(n_1219),
.B2(n_1275),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1296),
.B(n_1207),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1258),
.A2(n_1212),
.B1(n_1244),
.B2(n_1239),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1278),
.A2(n_1224),
.B(n_1238),
.C(n_1213),
.Y(n_1329)
);

BUFx2_ASAP7_75t_SL g1330 ( 
.A(n_1235),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1244),
.A2(n_1247),
.B1(n_1279),
.B2(n_1289),
.Y(n_1331)
);

BUFx8_ASAP7_75t_SL g1332 ( 
.A(n_1235),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1276),
.B(n_1218),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1278),
.A2(n_1271),
.B(n_1230),
.C(n_1248),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1252),
.B(n_1206),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1249),
.A2(n_1254),
.B(n_1220),
.C(n_1283),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1206),
.B(n_1306),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1256),
.B(n_1309),
.Y(n_1338)
);

AND2x4_ASAP7_75t_SL g1339 ( 
.A(n_1291),
.B(n_1211),
.Y(n_1339)
);

AND2x6_ASAP7_75t_L g1340 ( 
.A(n_1279),
.B(n_1289),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1240),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1208),
.B(n_1298),
.Y(n_1342)
);

NOR2xp67_ASAP7_75t_L g1343 ( 
.A(n_1208),
.B(n_1307),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1294),
.B(n_1301),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1233),
.B(n_1294),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1237),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1242),
.A2(n_1265),
.B1(n_1222),
.B2(n_1308),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1294),
.B(n_1301),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1272),
.A2(n_1301),
.B(n_1305),
.C(n_1240),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1265),
.A2(n_1222),
.B1(n_1268),
.B2(n_1217),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1259),
.A2(n_1280),
.B(n_1295),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1215),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1246),
.B(n_1253),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1262),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1233),
.B(n_1262),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1266),
.A2(n_1280),
.B1(n_1260),
.B2(n_1210),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1221),
.B(n_1261),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1221),
.B(n_1261),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1257),
.B(n_1251),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1260),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1257),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1210),
.A2(n_1241),
.B1(n_1273),
.B2(n_1263),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1210),
.A2(n_1241),
.B1(n_1273),
.B2(n_1263),
.Y(n_1363)
);

AND2x2_ASAP7_75t_SL g1364 ( 
.A(n_1245),
.B(n_1228),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1241),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1250),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1228),
.B(n_1234),
.Y(n_1367)
);

INVx5_ASAP7_75t_L g1368 ( 
.A(n_1245),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1204),
.B(n_1205),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1282),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1286),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1293),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1310),
.B(n_1264),
.Y(n_1373)
);

AOI221x1_ASAP7_75t_SL g1374 ( 
.A1(n_1285),
.A2(n_612),
.B1(n_783),
.B2(n_1203),
.C(n_1303),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1290),
.A2(n_1203),
.B(n_1115),
.C(n_1292),
.Y(n_1375)
);

OAI31xp33_ASAP7_75t_L g1376 ( 
.A1(n_1290),
.A2(n_1203),
.A3(n_612),
.B(n_973),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1277),
.A2(n_1168),
.B(n_867),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1208),
.B(n_1258),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1223),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1311),
.B(n_1377),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1373),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1320),
.B(n_1318),
.Y(n_1385)
);

BUFx2_ASAP7_75t_SL g1386 ( 
.A(n_1342),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1316),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1373),
.B(n_1359),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1380),
.B(n_1382),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1316),
.Y(n_1390)
);

BUFx8_ASAP7_75t_SL g1391 ( 
.A(n_1332),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1359),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1344),
.B(n_1348),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1364),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1321),
.B(n_1325),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1355),
.B(n_1367),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1365),
.B(n_1345),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1332),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1352),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1361),
.Y(n_1402)
);

NAND2x1p5_ASAP7_75t_L g1403 ( 
.A(n_1368),
.B(n_1366),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1341),
.B(n_1381),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1370),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1371),
.A2(n_1356),
.B(n_1369),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1336),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1336),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1372),
.A2(n_1322),
.B(n_1351),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1334),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1334),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1349),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1340),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1319),
.A2(n_1324),
.B(n_1350),
.Y(n_1414)
);

INVxp33_ASAP7_75t_L g1415 ( 
.A(n_1378),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1376),
.A2(n_1326),
.B1(n_1328),
.B2(n_1331),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1327),
.B(n_1338),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1314),
.B(n_1317),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1319),
.B(n_1313),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1314),
.A2(n_1324),
.B(n_1333),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1393),
.B(n_1312),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1413),
.B(n_1375),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1387),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1405),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1405),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1392),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1388),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1387),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1394),
.B(n_1323),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1388),
.Y(n_1430)
);

NAND2x1p5_ASAP7_75t_L g1431 ( 
.A(n_1413),
.B(n_1354),
.Y(n_1431)
);

AND2x2_ASAP7_75t_SL g1432 ( 
.A(n_1413),
.B(n_1322),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1402),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1390),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1383),
.B(n_1374),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1397),
.B(n_1335),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1397),
.B(n_1353),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1390),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1403),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1404),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1414),
.B(n_1379),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1412),
.B(n_1346),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1384),
.B(n_1315),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1424),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1435),
.A2(n_1419),
.B1(n_1385),
.B2(n_1415),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1435),
.A2(n_1416),
.B1(n_1419),
.B2(n_1313),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1427),
.B(n_1384),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1424),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1427),
.B(n_1384),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1427),
.B(n_1384),
.Y(n_1450)
);

AOI211x1_ASAP7_75t_L g1451 ( 
.A1(n_1443),
.A2(n_1396),
.B(n_1383),
.C(n_1389),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1441),
.A2(n_1414),
.B(n_1416),
.Y(n_1452)
);

AOI211xp5_ASAP7_75t_L g1453 ( 
.A1(n_1442),
.A2(n_1385),
.B(n_1375),
.C(n_1415),
.Y(n_1453)
);

AND2x4_ASAP7_75t_SL g1454 ( 
.A(n_1422),
.B(n_1413),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1441),
.B(n_1420),
.C(n_1329),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1427),
.B(n_1401),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1422),
.A2(n_1420),
.B1(n_1396),
.B2(n_1389),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1425),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1440),
.B(n_1412),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1433),
.A2(n_1406),
.B(n_1409),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1430),
.B(n_1395),
.Y(n_1462)
);

OAI33xp33_ASAP7_75t_L g1463 ( 
.A1(n_1442),
.A2(n_1410),
.A3(n_1411),
.B1(n_1407),
.B2(n_1408),
.B3(n_1417),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_SL g1464 ( 
.A(n_1442),
.B(n_1329),
.C(n_1399),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1426),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1428),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1422),
.A2(n_1414),
.B1(n_1420),
.B2(n_1418),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1422),
.A2(n_1420),
.B1(n_1411),
.B2(n_1410),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1440),
.B(n_1398),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1430),
.B(n_1436),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1431),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1429),
.B(n_1418),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1421),
.Y(n_1473)
);

NOR5xp2_ASAP7_75t_SL g1474 ( 
.A(n_1422),
.B(n_1347),
.C(n_1414),
.D(n_1420),
.E(n_1386),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1438),
.B(n_1398),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1426),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1439),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1444),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1452),
.B(n_1432),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1452),
.A2(n_1422),
.B(n_1407),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1444),
.Y(n_1481)
);

CKINVDCx16_ASAP7_75t_R g1482 ( 
.A(n_1464),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1461),
.A2(n_1455),
.B(n_1467),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1472),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1471),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1448),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1465),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1445),
.A2(n_1464),
.B(n_1446),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1465),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1476),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1471),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1457),
.B(n_1422),
.Y(n_1492)
);

INVx4_ASAP7_75t_SL g1493 ( 
.A(n_1471),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1476),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1459),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1456),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1460),
.B(n_1434),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1460),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1459),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1454),
.B(n_1439),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1466),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1502)
);

AOI33xp33_ASAP7_75t_L g1503 ( 
.A1(n_1482),
.A2(n_1445),
.A3(n_1453),
.B1(n_1418),
.B2(n_1401),
.B3(n_1443),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_SL g1504 ( 
.A(n_1488),
.B(n_1453),
.C(n_1457),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1488),
.B(n_1451),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_SL g1507 ( 
.A(n_1480),
.B(n_1446),
.C(n_1468),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1490),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1490),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1496),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1482),
.Y(n_1511)
);

INVxp67_ASAP7_75t_SL g1512 ( 
.A(n_1477),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1498),
.B(n_1451),
.Y(n_1513)
);

INVx6_ASAP7_75t_L g1514 ( 
.A(n_1490),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1497),
.B(n_1475),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1478),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1496),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1498),
.B(n_1429),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1490),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1484),
.B(n_1447),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1479),
.A2(n_1468),
.B1(n_1432),
.B2(n_1473),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1498),
.B(n_1429),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

NAND4xp25_ASAP7_75t_L g1527 ( 
.A(n_1480),
.B(n_1343),
.C(n_1417),
.D(n_1443),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1496),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1481),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1479),
.B(n_1437),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1493),
.B(n_1447),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1499),
.Y(n_1532)
);

AND2x2_ASAP7_75t_SL g1533 ( 
.A(n_1483),
.B(n_1432),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1493),
.B(n_1449),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1485),
.B(n_1391),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1493),
.B(n_1449),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1493),
.B(n_1450),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1497),
.B(n_1437),
.Y(n_1541)
);

NAND2x1_ASAP7_75t_L g1542 ( 
.A(n_1477),
.B(n_1462),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1493),
.B(n_1454),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1503),
.B(n_1487),
.Y(n_1544)
);

AO21x1_ASAP7_75t_L g1545 ( 
.A1(n_1512),
.A2(n_1499),
.B(n_1495),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1511),
.A2(n_1492),
.B1(n_1483),
.B2(n_1500),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1511),
.B(n_1493),
.Y(n_1547)
);

AOI211xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1504),
.A2(n_1474),
.B(n_1501),
.C(n_1495),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1506),
.B(n_1487),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1511),
.B(n_1491),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1541),
.B(n_1502),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_1489),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1511),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1536),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1543),
.B(n_1491),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1532),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1510),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1483),
.C(n_1492),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1516),
.Y(n_1559)
);

OAI21xp33_ASAP7_75t_L g1560 ( 
.A1(n_1507),
.A2(n_1492),
.B(n_1494),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1513),
.B(n_1489),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1516),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1535),
.B(n_1501),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1517),
.B(n_1502),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1517),
.B(n_1502),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1543),
.B(n_1490),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1518),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1535),
.B(n_1437),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1485),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1510),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1505),
.B(n_1490),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1530),
.B(n_1436),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1518),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1519),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1519),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1522),
.Y(n_1576)
);

NAND2xp67_ASAP7_75t_L g1577 ( 
.A(n_1528),
.B(n_1339),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1527),
.B(n_1330),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1559),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1554),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1562),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1556),
.B(n_1520),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1547),
.B(n_1505),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1558),
.A2(n_1533),
.B1(n_1492),
.B2(n_1483),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1555),
.B(n_1515),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1567),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1555),
.B(n_1533),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1550),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1573),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1569),
.B(n_1550),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1553),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1569),
.B(n_1523),
.Y(n_1593)
);

AND2x2_ASAP7_75t_SL g1594 ( 
.A(n_1544),
.B(n_1483),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1548),
.B(n_1525),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1578),
.B(n_1400),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1566),
.B(n_1571),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1576),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1549),
.B(n_1528),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1566),
.B(n_1490),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1561),
.B(n_1523),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1552),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1557),
.Y(n_1603)
);

AOI32xp33_ASAP7_75t_L g1604 ( 
.A1(n_1585),
.A2(n_1560),
.A3(n_1546),
.B1(n_1578),
.B2(n_1571),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1601),
.B(n_1563),
.Y(n_1605)
);

NAND2x1_ASAP7_75t_L g1606 ( 
.A(n_1583),
.B(n_1566),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1603),
.Y(n_1607)
);

AOI31xp33_ASAP7_75t_L g1608 ( 
.A1(n_1589),
.A2(n_1545),
.A3(n_1571),
.B(n_1574),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1603),
.Y(n_1609)
);

AOI322xp5_ASAP7_75t_L g1610 ( 
.A1(n_1580),
.A2(n_1542),
.A3(n_1568),
.B1(n_1545),
.B2(n_1574),
.C1(n_1557),
.C2(n_1570),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1592),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1570),
.Y(n_1612)
);

AOI322xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1588),
.A2(n_1474),
.A3(n_1542),
.B1(n_1463),
.B2(n_1539),
.C1(n_1538),
.C2(n_1531),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1579),
.Y(n_1614)
);

A2O1A1Ixp33_ASAP7_75t_SL g1615 ( 
.A1(n_1595),
.A2(n_1575),
.B(n_1508),
.C(n_1526),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1579),
.Y(n_1616)
);

O2A1O1Ixp5_ASAP7_75t_L g1617 ( 
.A1(n_1600),
.A2(n_1526),
.B(n_1508),
.C(n_1575),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1583),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1602),
.B(n_1591),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1596),
.A2(n_1526),
.B(n_1508),
.Y(n_1620)
);

OAI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1594),
.A2(n_1492),
.B(n_1577),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1531),
.Y(n_1622)
);

AOI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1594),
.A2(n_1509),
.B(n_1564),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1618),
.B(n_1586),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1611),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1622),
.B(n_1593),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1606),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1608),
.A2(n_1584),
.B(n_1583),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1619),
.B(n_1593),
.Y(n_1629)
);

INVxp67_ASAP7_75t_SL g1630 ( 
.A(n_1619),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1612),
.B(n_1586),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1584),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1610),
.B(n_1584),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1607),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1628),
.A2(n_1615),
.B(n_1617),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1630),
.A2(n_1588),
.B1(n_1621),
.B2(n_1597),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1633),
.B(n_1604),
.C(n_1620),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_SL g1638 ( 
.A(n_1629),
.B(n_1620),
.C(n_1613),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1626),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1614),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1631),
.A2(n_1599),
.B(n_1597),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1626),
.Y(n_1642)
);

XNOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1632),
.B(n_1605),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1637),
.A2(n_1632),
.B(n_1624),
.Y(n_1644)
);

AOI222xp33_ASAP7_75t_L g1645 ( 
.A1(n_1638),
.A2(n_1625),
.B1(n_1634),
.B2(n_1616),
.C1(n_1627),
.C2(n_1609),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1636),
.A2(n_1627),
.B1(n_1582),
.B2(n_1514),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1635),
.A2(n_1639),
.B1(n_1642),
.B2(n_1641),
.C(n_1587),
.Y(n_1647)
);

OAI311xp33_ASAP7_75t_L g1648 ( 
.A1(n_1643),
.A2(n_1598),
.A3(n_1587),
.B1(n_1581),
.C1(n_1590),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1645),
.B(n_1640),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1644),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1647),
.B(n_1581),
.Y(n_1651)
);

BUFx4f_ASAP7_75t_SL g1652 ( 
.A(n_1646),
.Y(n_1652)
);

XOR2xp5_ASAP7_75t_L g1653 ( 
.A(n_1648),
.B(n_1360),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1646),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1652),
.Y(n_1655)
);

XOR2xp5_ASAP7_75t_L g1656 ( 
.A(n_1653),
.B(n_1590),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1650),
.A2(n_1598),
.B1(n_1514),
.B2(n_1521),
.Y(n_1657)
);

AND4x1_ASAP7_75t_L g1658 ( 
.A(n_1649),
.B(n_1534),
.C(n_1539),
.D(n_1538),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1654),
.Y(n_1659)
);

XNOR2xp5_ASAP7_75t_L g1660 ( 
.A(n_1658),
.B(n_1651),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1659),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1655),
.B(n_1509),
.C(n_1564),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1661),
.B(n_1656),
.Y(n_1663)
);

OAI221xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1663),
.A2(n_1657),
.B1(n_1660),
.B2(n_1662),
.C(n_1565),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1664),
.Y(n_1665)
);

OR3x1_ASAP7_75t_L g1666 ( 
.A(n_1664),
.B(n_1463),
.C(n_1522),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1665),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1666),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1667),
.A2(n_1565),
.B1(n_1514),
.B2(n_1521),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1668),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1670),
.Y(n_1671)
);

AOI22x1_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1669),
.B1(n_1337),
.B2(n_1551),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_SL g1673 ( 
.A(n_1672),
.B(n_1572),
.C(n_1537),
.Y(n_1673)
);

OAI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1673),
.A2(n_1521),
.B1(n_1514),
.B2(n_1551),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1521),
.B1(n_1534),
.B2(n_1529),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1540),
.B1(n_1537),
.B2(n_1529),
.Y(n_1676)
);


endmodule