module fake_jpeg_1595_n_127 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_127);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_16),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_44),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_13),
.B(n_14),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_17),
.A3(n_25),
.B1(n_19),
.B2(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_25),
.B1(n_19),
.B2(n_15),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_31),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_9),
.B1(n_11),
.B2(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_32),
.B1(n_38),
.B2(n_64),
.Y(n_75)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_28),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_55),
.B1(n_66),
.B2(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_55),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_52),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_84),
.C(n_81),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_60),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_47),
.Y(n_85)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_76),
.B(n_70),
.C(n_84),
.D(n_80),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_82),
.B(n_69),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_61),
.C(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_84),
.C(n_71),
.Y(n_99)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_88),
.B1(n_95),
.B2(n_91),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_105),
.B(n_94),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

AOI21x1_ASAP7_75t_L g113 ( 
.A1(n_108),
.A2(n_111),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_70),
.B1(n_85),
.B2(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_97),
.B1(n_83),
.B2(n_100),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_93),
.B(n_95),
.C(n_77),
.D(n_63),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_116),
.B(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_98),
.C(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_100),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_65),
.A3(n_68),
.B1(n_90),
.B2(n_100),
.C1(n_114),
.C2(n_117),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_122),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_114),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_90),
.Y(n_127)
);


endmodule