module fake_netlist_6_4718_n_1565 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1565);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1565;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

BUFx10_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_48),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_51),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_46),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_1),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_87),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_30),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_70),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_78),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_41),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_41),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_52),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_40),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_23),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_31),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_73),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_24),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_1),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_115),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_91),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_26),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_72),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_26),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_23),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_49),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_92),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_105),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_122),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_135),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_7),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_16),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_106),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_64),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_8),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_3),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_101),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_42),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_53),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_54),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_74),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_18),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_47),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_2),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_50),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_44),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_139),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_119),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_60),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_38),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_28),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_22),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_125),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_100),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_142),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_62),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_63),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_16),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_114),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_19),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_104),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_38),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_89),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_137),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_18),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_75),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_103),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_99),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_33),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_27),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_128),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_35),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_57),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_111),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_35),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_71),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_97),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_6),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_82),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_15),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_124),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_45),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_76),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_69),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_94),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_13),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_68),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_116),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_61),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_31),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_56),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_15),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_79),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_39),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_17),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_12),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_34),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_123),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_9),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_43),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_6),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_81),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_19),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_107),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_229),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_187),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_274),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_274),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_R g306 ( 
.A(n_242),
.B(n_55),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_265),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_178),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_172),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_172),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_195),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_201),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_205),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_169),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_256),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_178),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_189),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_178),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_188),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_209),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_178),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_222),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_178),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_196),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_211),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_214),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_213),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_278),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_183),
.B(n_3),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_197),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_198),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_199),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_233),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_173),
.B(n_4),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_200),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_234),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_202),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_154),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_185),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_235),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_186),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_190),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_238),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_203),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_204),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_206),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_246),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_173),
.B(n_5),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_166),
.B(n_8),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_255),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_162),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_239),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_248),
.B(n_10),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_192),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_224),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_162),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_255),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_151),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_151),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_251),
.Y(n_370)
);

NAND2xp33_ASAP7_75t_R g371 ( 
.A(n_153),
.B(n_11),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_207),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_228),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_208),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_R g376 ( 
.A(n_320),
.B(n_212),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_308),
.B(n_153),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_323),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_315),
.B(n_155),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_326),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_307),
.B(n_170),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_366),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_337),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_308),
.B(n_155),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_339),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_157),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_340),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_325),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_344),
.B(n_216),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_333),
.B(n_157),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_245),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_302),
.B(n_158),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_346),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_243),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_354),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_355),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_373),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_316),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_375),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_368),
.B(n_158),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_R g425 ( 
.A(n_312),
.B(n_219),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_313),
.B(n_161),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_367),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_332),
.B(n_213),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_301),
.B(n_161),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_313),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_336),
.B(n_151),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_314),
.B(n_164),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_314),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_321),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_360),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_374),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_318),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_304),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_309),
.B(n_215),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_310),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_388),
.Y(n_448)
);

BUFx4f_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_321),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_389),
.B(n_366),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_305),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_407),
.B(n_327),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_404),
.Y(n_456)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_435),
.B(n_359),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_434),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_327),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_435),
.B(n_166),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_407),
.B(n_329),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_329),
.Y(n_466)
);

BUFx4f_ASAP7_75t_L g467 ( 
.A(n_400),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_415),
.B(n_369),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_407),
.B(n_341),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_430),
.B(n_184),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_381),
.B(n_184),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_381),
.B(n_217),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_407),
.B(n_341),
.Y(n_474)
);

AND3x2_ASAP7_75t_L g475 ( 
.A(n_415),
.B(n_356),
.C(n_218),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_433),
.B(n_180),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_402),
.B(n_345),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_392),
.B(n_345),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_405),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_446),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_442),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_420),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_392),
.B(n_349),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_437),
.B(n_217),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_426),
.A2(n_370),
.B1(n_362),
.B2(n_353),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_402),
.B(n_349),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_389),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_445),
.B(n_218),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_445),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_446),
.B(n_362),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_259),
.B1(n_292),
.B2(n_294),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_403),
.B(n_311),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_419),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_445),
.B(n_259),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_436),
.B(n_324),
.Y(n_499)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

OR2x2_ASAP7_75t_SL g502 ( 
.A(n_396),
.B(n_250),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_425),
.B(n_245),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_431),
.B(n_328),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_378),
.B(n_215),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_377),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_403),
.B(n_330),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_377),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_431),
.B(n_347),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_363),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_379),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_378),
.B(n_280),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_376),
.B(n_306),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_422),
.B(n_280),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_421),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_378),
.B(n_293),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_406),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_422),
.B(n_293),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_385),
.B(n_348),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_382),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_406),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_401),
.B(n_245),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_406),
.Y(n_527)
);

XNOR2x2_ASAP7_75t_L g528 ( 
.A(n_423),
.B(n_295),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_379),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_380),
.B(n_386),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_391),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_443),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_386),
.B(n_350),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_387),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_378),
.B(n_252),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_390),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_439),
.B(n_351),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_SL g540 ( 
.A1(n_393),
.A2(n_279),
.B(n_257),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_429),
.B(n_364),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_439),
.A2(n_299),
.B1(n_284),
.B2(n_286),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_394),
.Y(n_543)
);

BUFx10_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_393),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_398),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_439),
.B(n_365),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_406),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_414),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_406),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_296),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_441),
.A2(n_289),
.B1(n_245),
.B2(n_262),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_427),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_411),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_441),
.B(n_165),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_441),
.B(n_262),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_383),
.B(n_384),
.Y(n_560)
);

HAxp5_ASAP7_75t_SL g561 ( 
.A(n_413),
.B(n_152),
.CON(n_561),
.SN(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_410),
.B(n_262),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_410),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_429),
.A2(n_262),
.B1(n_300),
.B2(n_232),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_416),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_SL g567 ( 
.A(n_418),
.B(n_371),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_432),
.A2(n_262),
.B1(n_237),
.B2(n_231),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_432),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_432),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_383),
.B(n_223),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_428),
.B(n_254),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_383),
.B(n_230),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_428),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_409),
.A2(n_179),
.B1(n_156),
.B2(n_160),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_417),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_448),
.B(n_399),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_450),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_448),
.B(n_159),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_456),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_488),
.B(n_163),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_457),
.A2(n_487),
.B1(n_480),
.B2(n_455),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_452),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_399),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_451),
.A2(n_478),
.B1(n_460),
.B2(n_457),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_490),
.A2(n_194),
.B1(n_221),
.B2(n_220),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_488),
.B(n_165),
.Y(n_587)
);

AND2x6_ASAP7_75t_SL g588 ( 
.A(n_468),
.B(n_168),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_460),
.B(n_175),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_478),
.B(n_399),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_494),
.B(n_175),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_459),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_465),
.B(n_176),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_491),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_510),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_523),
.B(n_181),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_576),
.B(n_384),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_466),
.B(n_193),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_499),
.A2(n_236),
.B1(n_258),
.B2(n_240),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_561),
.A2(n_288),
.B1(n_225),
.B2(n_297),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_517),
.B(n_181),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_461),
.B(n_182),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_513),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_512),
.B(n_384),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_538),
.B(n_182),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_532),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_479),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_505),
.B(n_410),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_410),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_483),
.Y(n_613)
);

OAI22x1_ASAP7_75t_SL g614 ( 
.A1(n_533),
.A2(n_177),
.B1(n_174),
.B2(n_297),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_482),
.B(n_167),
.Y(n_615)
);

BUFx8_ASAP7_75t_L g616 ( 
.A(n_566),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_447),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_501),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_499),
.A2(n_253),
.B1(n_241),
.B2(n_249),
.Y(n_619)
);

NOR2x1_ASAP7_75t_L g620 ( 
.A(n_469),
.B(n_210),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_461),
.B(n_226),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_503),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_449),
.B(n_226),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_523),
.B(n_268),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_496),
.B(n_167),
.Y(n_625)
);

NOR2x1p5_ASAP7_75t_L g626 ( 
.A(n_482),
.B(n_171),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_244),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_558),
.B(n_264),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_569),
.B(n_273),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_456),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_554),
.B(n_271),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_508),
.B(n_271),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_507),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_570),
.B(n_275),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_509),
.B(n_267),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_453),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g637 ( 
.A(n_489),
.B(n_247),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_515),
.B(n_287),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_529),
.B(n_534),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_471),
.A2(n_417),
.B(n_298),
.C(n_270),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_531),
.B(n_417),
.Y(n_641)
);

BUFx8_ASAP7_75t_L g642 ( 
.A(n_518),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_449),
.B(n_270),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_474),
.B(n_276),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_567),
.A2(n_514),
.B1(n_470),
.B2(n_572),
.Y(n_645)
);

AND2x6_ASAP7_75t_SL g646 ( 
.A(n_468),
.B(n_291),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_506),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_453),
.B(n_276),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_467),
.B(n_291),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_555),
.A2(n_266),
.B1(n_283),
.B2(n_174),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_467),
.B(n_277),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_514),
.B(n_285),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_555),
.A2(n_269),
.B1(n_283),
.B2(n_177),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_458),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_458),
.Y(n_655)
);

OAI221xp5_ASAP7_75t_L g656 ( 
.A1(n_495),
.A2(n_269),
.B1(n_225),
.B2(n_260),
.C(n_261),
.Y(n_656)
);

NOR3xp33_ASAP7_75t_L g657 ( 
.A(n_463),
.B(n_272),
.C(n_260),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_463),
.B(n_272),
.C(n_261),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_497),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_454),
.B(n_285),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_471),
.A2(n_472),
.B(n_504),
.C(n_559),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_526),
.B(n_282),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_518),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_520),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_539),
.B(n_281),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_541),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_484),
.B(n_266),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_484),
.B(n_263),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_526),
.B(n_263),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_171),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_545),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_504),
.B(n_11),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_537),
.B(n_12),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_502),
.B(n_13),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_486),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_560),
.B(n_83),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_546),
.B(n_148),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_519),
.B(n_20),
.C(n_21),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_528),
.B(n_20),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_536),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_547),
.B(n_548),
.Y(n_682)
);

BUFx12f_ASAP7_75t_L g683 ( 
.A(n_524),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_550),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_522),
.B(n_93),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_552),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_470),
.A2(n_66),
.B1(n_146),
.B2(n_141),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_468),
.B(n_21),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_470),
.A2(n_58),
.B1(n_140),
.B2(n_136),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_553),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_462),
.B(n_147),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_541),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_556),
.Y(n_693)
);

AOI221xp5_ASAP7_75t_L g694 ( 
.A1(n_495),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.C(n_29),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_477),
.B(n_25),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_542),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_696)
);

OAI221xp5_ASAP7_75t_L g697 ( 
.A1(n_542),
.A2(n_32),
.B1(n_37),
.B2(n_40),
.C(n_43),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_470),
.A2(n_109),
.B1(n_130),
.B2(n_95),
.Y(n_698)
);

CKINVDCx11_ASAP7_75t_R g699 ( 
.A(n_524),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_571),
.B(n_96),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_565),
.B(n_98),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_565),
.A2(n_113),
.B1(n_126),
.B2(n_134),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_475),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_37),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_535),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_563),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_535),
.A2(n_540),
.B1(n_500),
.B2(n_498),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_544),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_481),
.B(n_568),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_477),
.B(n_543),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_568),
.B(n_500),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_475),
.B(n_500),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_544),
.B(n_557),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_574),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_521),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_SL g717 ( 
.A1(n_680),
.A2(n_557),
.B1(n_575),
.B2(n_473),
.Y(n_717)
);

CKINVDCx8_ASAP7_75t_R g718 ( 
.A(n_646),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_583),
.B(n_493),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_681),
.B(n_549),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_580),
.B(n_527),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_579),
.A2(n_492),
.B1(n_575),
.B2(n_562),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_696),
.A2(n_562),
.B1(n_485),
.B2(n_511),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_582),
.A2(n_549),
.B1(n_564),
.B2(n_521),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_594),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_577),
.B(n_521),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_630),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_692),
.B(n_525),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_578),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_589),
.B(n_530),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_592),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_595),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_632),
.B(n_530),
.Y(n_733)
);

OAI321xp33_ASAP7_75t_L g734 ( 
.A1(n_680),
.A2(n_551),
.A3(n_697),
.B1(n_602),
.B2(n_696),
.C(n_694),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_716),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_625),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_676),
.Y(n_737)
);

AND2x2_ASAP7_75t_SL g738 ( 
.A(n_623),
.B(n_643),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_655),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_682),
.A2(n_590),
.B(n_584),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_636),
.B(n_667),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_581),
.A2(n_674),
.B(n_673),
.C(n_628),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_615),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_607),
.A2(n_708),
.B(n_581),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_603),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_716),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_671),
.B(n_587),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_692),
.B(n_664),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_645),
.A2(n_663),
.B1(n_647),
.B2(n_665),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_671),
.B(n_652),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_652),
.B(n_649),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_713),
.A2(n_621),
.B(n_604),
.C(n_610),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_669),
.B(n_597),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_641),
.A2(n_598),
.B(n_639),
.Y(n_754)
);

O2A1O1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_586),
.A2(n_660),
.B(n_644),
.C(n_666),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_613),
.B(n_618),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_622),
.B(n_633),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_627),
.A2(n_599),
.B(n_593),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_672),
.B(n_684),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_659),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_686),
.B(n_648),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_701),
.A2(n_620),
.B(n_700),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_690),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_604),
.B(n_621),
.C(n_657),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_677),
.A2(n_660),
.B(n_685),
.Y(n_765)
);

OAI321xp33_ASAP7_75t_L g766 ( 
.A1(n_675),
.A2(n_656),
.A3(n_650),
.B1(n_653),
.B2(n_668),
.C(n_624),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_648),
.B(n_715),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_690),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_693),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_676),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_635),
.B(n_638),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_707),
.A2(n_705),
.B(n_617),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_596),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_629),
.B(n_634),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_591),
.B(n_608),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_667),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_608),
.B(n_695),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_605),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_606),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_651),
.B(n_704),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_601),
.B(n_619),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_667),
.B(n_626),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_609),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_640),
.A2(n_691),
.B(n_702),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_662),
.B(n_713),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_658),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_667),
.B(n_637),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_678),
.A2(n_688),
.B(n_711),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_687),
.A2(n_698),
.B(n_689),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_670),
.A2(n_675),
.B(n_714),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_614),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_653),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_679),
.A2(n_642),
.B(n_588),
.C(n_616),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_642),
.B(n_683),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_709),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_585),
.A2(n_448),
.B(n_661),
.C(n_460),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_585),
.A2(n_448),
.B(n_661),
.C(n_460),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_585),
.B(n_488),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_654),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_R g800 ( 
.A(n_699),
.B(n_538),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_585),
.B(n_488),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_706),
.B(n_448),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_585),
.A2(n_696),
.B1(n_706),
.B2(n_448),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_SL g804 ( 
.A(n_681),
.B(n_538),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_654),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_585),
.A2(n_696),
.B1(n_706),
.B2(n_448),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_706),
.B(n_448),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_582),
.A2(n_710),
.B(n_661),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_632),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_683),
.B(n_538),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_706),
.B(n_448),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_699),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_585),
.B(n_488),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_706),
.B(n_448),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_706),
.B(n_448),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_654),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_578),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_582),
.A2(n_710),
.B(n_661),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_582),
.A2(n_710),
.B(n_661),
.Y(n_822)
);

INVx5_ASAP7_75t_L g823 ( 
.A(n_716),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_585),
.A2(n_696),
.B1(n_706),
.B2(n_448),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_706),
.B(n_448),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_585),
.B(n_448),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_631),
.B(n_494),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_626),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_667),
.Y(n_831)
);

OA22x2_ASAP7_75t_L g832 ( 
.A1(n_585),
.A2(n_602),
.B1(n_579),
.B2(n_706),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_585),
.B(n_448),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_699),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_585),
.A2(n_696),
.B1(n_706),
.B2(n_448),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_582),
.A2(n_710),
.B(n_661),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_578),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_630),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_585),
.B(n_488),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_585),
.B(n_448),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_585),
.A2(n_448),
.B(n_661),
.C(n_460),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_667),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_585),
.B(n_448),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_667),
.Y(n_848)
);

CKINVDCx10_ASAP7_75t_R g849 ( 
.A(n_699),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_582),
.A2(n_710),
.B(n_661),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_626),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_582),
.A2(n_710),
.B(n_661),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_594),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_706),
.B(n_448),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_712),
.A2(n_612),
.B(n_611),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_706),
.B(n_448),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_585),
.B(n_488),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_765),
.A2(n_813),
.B(n_807),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_827),
.B(n_833),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_818),
.A2(n_828),
.B(n_825),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_842),
.B(n_847),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_802),
.B(n_808),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_751),
.A2(n_781),
.B1(n_750),
.B2(n_747),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_829),
.B(n_736),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_737),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_812),
.B(n_816),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_796),
.A2(n_844),
.B(n_797),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_803),
.A2(n_836),
.B(n_824),
.C(n_806),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_817),
.B(n_826),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_770),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_721),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_795),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_854),
.A2(n_856),
.B(n_804),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_777),
.B(n_810),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_803),
.A2(n_806),
.B(n_824),
.C(n_836),
.Y(n_875)
);

OA22x2_ASAP7_75t_L g876 ( 
.A1(n_792),
.A2(n_798),
.B1(n_801),
.B2(n_815),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_738),
.B(n_761),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_729),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_776),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_764),
.A2(n_766),
.B(n_755),
.C(n_742),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_795),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_841),
.A2(n_857),
.B(n_784),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_725),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_800),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_795),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_782),
.B(n_748),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_743),
.B(n_745),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_752),
.A2(n_749),
.B(n_753),
.C(n_789),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_717),
.B(n_767),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_835),
.A2(n_855),
.B(n_845),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_853),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_775),
.B(n_720),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_733),
.B(n_771),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_840),
.A2(n_843),
.B(n_758),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_754),
.B(n_774),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_776),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_740),
.A2(n_726),
.B(n_762),
.Y(n_897)
);

AOI21xp33_ASAP7_75t_L g898 ( 
.A1(n_832),
.A2(n_734),
.B(n_850),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_776),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_832),
.A2(n_722),
.B1(n_850),
.B2(n_809),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_780),
.B(n_744),
.C(n_790),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_748),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_809),
.A2(n_852),
.B(n_837),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_785),
.A2(n_786),
.B1(n_787),
.B2(n_719),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_830),
.Y(n_905)
);

AO31x2_ASAP7_75t_L g906 ( 
.A1(n_723),
.A2(n_730),
.A3(n_772),
.B(n_768),
.Y(n_906)
);

AND3x4_ASAP7_75t_L g907 ( 
.A(n_811),
.B(n_728),
.C(n_718),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_821),
.A2(n_852),
.B(n_837),
.Y(n_908)
);

INVx8_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_821),
.A2(n_822),
.B1(n_723),
.B2(n_756),
.Y(n_910)
);

NOR2x1_ASAP7_75t_SL g911 ( 
.A(n_823),
.B(n_848),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_757),
.B(n_759),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_731),
.B(n_820),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_839),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_732),
.B(n_838),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_724),
.A2(n_778),
.B(n_769),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_799),
.B(n_819),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_851),
.B(n_728),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_741),
.A2(n_846),
.B1(n_831),
.B2(n_848),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_831),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_846),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_846),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_823),
.A2(n_746),
.B(n_735),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_848),
.B(n_823),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_739),
.B(n_760),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_773),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_779),
.B(n_783),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_823),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_805),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_788),
.B(n_791),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_793),
.A2(n_794),
.B(n_814),
.C(n_834),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_849),
.B(n_827),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_827),
.B(n_833),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_827),
.A2(n_842),
.B1(n_847),
.B2(n_833),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_796),
.A2(n_844),
.B(n_797),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_776),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_829),
.B(n_631),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_776),
.B(n_831),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_782),
.B(n_580),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_725),
.Y(n_940)
);

O2A1O1Ixp5_ASAP7_75t_L g941 ( 
.A1(n_827),
.A2(n_579),
.B(n_842),
.C(n_833),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_827),
.A2(n_842),
.B1(n_847),
.B2(n_833),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_725),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_827),
.A2(n_842),
.B(n_847),
.C(n_833),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_765),
.A2(n_712),
.B(n_807),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_827),
.B(n_833),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_827),
.B(n_833),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_827),
.B(n_833),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_827),
.B(n_833),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_729),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_827),
.B(n_833),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_721),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_829),
.B(n_631),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_829),
.B(n_631),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_829),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_827),
.A2(n_842),
.B(n_847),
.C(n_833),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_796),
.A2(n_844),
.B(n_797),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_737),
.Y(n_958)
);

NAND2x1_ASAP7_75t_L g959 ( 
.A(n_727),
.B(n_716),
.Y(n_959)
);

AO31x2_ASAP7_75t_L g960 ( 
.A1(n_796),
.A2(n_797),
.A3(n_844),
.B(n_813),
.Y(n_960)
);

AOI221x1_ASAP7_75t_L g961 ( 
.A1(n_796),
.A2(n_797),
.B1(n_844),
.B2(n_842),
.C(n_833),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_725),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_725),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_796),
.A2(n_797),
.A3(n_844),
.B(n_813),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_L g965 ( 
.A(n_803),
.B(n_806),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_796),
.A2(n_844),
.B(n_797),
.Y(n_966)
);

AO21x1_ASAP7_75t_L g967 ( 
.A1(n_827),
.A2(n_842),
.B(n_833),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_765),
.A2(n_712),
.B(n_807),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_721),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_827),
.B(n_833),
.Y(n_970)
);

OAI22x1_ASAP7_75t_L g971 ( 
.A1(n_750),
.A2(n_585),
.B1(n_833),
.B2(n_827),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_765),
.A2(n_712),
.B(n_807),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_738),
.B(n_585),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_859),
.B(n_861),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_L g975 ( 
.A(n_863),
.B(n_965),
.C(n_956),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_884),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_950),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_SL g978 ( 
.A(n_934),
.B(n_942),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_L g979 ( 
.A(n_944),
.B(n_941),
.C(n_875),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_918),
.B(n_902),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_946),
.B(n_947),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_913),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_948),
.B(n_949),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_934),
.A2(n_942),
.B1(n_970),
.B2(n_951),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_915),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_933),
.B(n_967),
.Y(n_986)
);

AO21x2_ASAP7_75t_L g987 ( 
.A1(n_867),
.A2(n_935),
.B(n_957),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_862),
.A2(n_869),
.B1(n_888),
.B2(n_868),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_891),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_873),
.B(n_892),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_881),
.Y(n_991)
);

AOI222xp33_ASAP7_75t_L g992 ( 
.A1(n_971),
.A2(n_903),
.B1(n_908),
.B2(n_973),
.C1(n_900),
.C2(n_889),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_880),
.A2(n_898),
.B(n_903),
.C(n_908),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_879),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_858),
.A2(n_894),
.B(n_897),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_963),
.Y(n_996)
);

AOI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_877),
.A2(n_866),
.B(n_930),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_926),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_955),
.B(n_874),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_937),
.B(n_953),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_883),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_945),
.A2(n_972),
.B(n_968),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_954),
.B(n_864),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_958),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_883),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_909),
.B(n_924),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_909),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_879),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_955),
.B(n_912),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_887),
.B(n_870),
.Y(n_1010)
);

AOI221xp5_ASAP7_75t_L g1011 ( 
.A1(n_910),
.A2(n_935),
.B1(n_966),
.B2(n_957),
.C(n_867),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_893),
.A2(n_904),
.B1(n_901),
.B2(n_966),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_870),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_961),
.B(n_882),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_865),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_940),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_871),
.B(n_969),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_865),
.B(n_943),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_952),
.B(n_969),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_909),
.B(n_924),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_962),
.B(n_932),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_925),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_876),
.A2(n_905),
.B(n_916),
.Y(n_1023)
);

AOI21xp33_ASAP7_75t_SL g1024 ( 
.A1(n_907),
.A2(n_876),
.B(n_931),
.Y(n_1024)
);

INVx8_ASAP7_75t_L g1025 ( 
.A(n_896),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_922),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_927),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_920),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_899),
.B(n_929),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_872),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_921),
.B(n_919),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_914),
.B(n_921),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_960),
.B(n_964),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_938),
.B(n_964),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_917),
.B(n_906),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_896),
.A2(n_936),
.B1(n_959),
.B2(n_923),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_936),
.B(n_906),
.Y(n_1037)
);

AND2x2_ASAP7_75t_SL g1038 ( 
.A(n_911),
.B(n_885),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_937),
.B(n_953),
.Y(n_1039)
);

NOR2xp67_ASAP7_75t_L g1040 ( 
.A(n_904),
.B(n_764),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_886),
.B(n_939),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_859),
.B(n_861),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_937),
.B(n_953),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_859),
.B(n_861),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_SL g1045 ( 
.A1(n_934),
.A2(n_750),
.B1(n_476),
.B2(n_448),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_859),
.B(n_861),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_879),
.Y(n_1047)
);

BUFx4_ASAP7_75t_SL g1048 ( 
.A(n_881),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_884),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_909),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_859),
.B(n_861),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_909),
.B(n_958),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_958),
.Y(n_1053)
);

BUFx8_ASAP7_75t_L g1054 ( 
.A(n_872),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_881),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_958),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_859),
.B(n_861),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_891),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_859),
.B(n_861),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_879),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_859),
.B(n_861),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_884),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_928),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_872),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_934),
.A2(n_942),
.B1(n_833),
.B2(n_842),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_937),
.B(n_953),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_944),
.A2(n_956),
.B(n_448),
.C(n_942),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_867),
.A2(n_957),
.B(n_935),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_895),
.A2(n_890),
.B(n_860),
.Y(n_1069)
);

CKINVDCx16_ASAP7_75t_R g1070 ( 
.A(n_872),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_886),
.B(n_939),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_937),
.B(n_953),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_963),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_881),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_859),
.B(n_861),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_958),
.Y(n_1076)
);

OR2x6_ASAP7_75t_SL g1077 ( 
.A(n_884),
.B(n_538),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_863),
.A2(n_833),
.B(n_842),
.C(n_827),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_883),
.Y(n_1079)
);

NOR2xp67_ASAP7_75t_SL g1080 ( 
.A(n_872),
.B(n_683),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_963),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_859),
.B(n_861),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_878),
.Y(n_1083)
);

OR2x6_ASAP7_75t_L g1084 ( 
.A(n_909),
.B(n_958),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_859),
.B(n_861),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_863),
.B(n_449),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_878),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1000),
.B(n_1039),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_991),
.Y(n_1089)
);

INVx5_ASAP7_75t_L g1090 ( 
.A(n_1006),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1083),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1065),
.A2(n_1045),
.B1(n_1078),
.B2(n_1085),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1001),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1065),
.A2(n_981),
.B1(n_1082),
.B2(n_974),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_SL g1095 ( 
.A1(n_978),
.A2(n_975),
.B1(n_984),
.B2(n_979),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_978),
.A2(n_983),
.B1(n_1061),
.B2(n_1042),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_1034),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_1001),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_1054),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1048),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1087),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1044),
.B(n_1046),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_998),
.Y(n_1103)
);

AO21x2_ASAP7_75t_L g1104 ( 
.A1(n_995),
.A2(n_1002),
.B(n_1069),
.Y(n_1104)
);

INVxp33_ASAP7_75t_L g1105 ( 
.A(n_1010),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1017),
.B(n_1019),
.Y(n_1106)
);

BUFx4_ASAP7_75t_SL g1107 ( 
.A(n_1049),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1043),
.B(n_1066),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_SL g1109 ( 
.A1(n_975),
.A2(n_984),
.B1(n_979),
.B2(n_986),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_992),
.A2(n_1011),
.B1(n_988),
.B2(n_1040),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_982),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_1055),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_992),
.A2(n_1040),
.B1(n_1086),
.B2(n_987),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1075),
.A2(n_1059),
.B1(n_1051),
.B2(n_1057),
.Y(n_1115)
);

CKINVDCx11_ASAP7_75t_R g1116 ( 
.A(n_1077),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1006),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1013),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1022),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1027),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1009),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_1007),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1029),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_1054),
.Y(n_1124)
);

BUFx2_ASAP7_75t_SL g1125 ( 
.A(n_1062),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1006),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1068),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_999),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_1007),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_R g1130 ( 
.A(n_1068),
.B(n_1024),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_SL g1131 ( 
.A(n_976),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1067),
.A2(n_990),
.B1(n_1015),
.B2(n_993),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1004),
.Y(n_1133)
);

CKINVDCx16_ASAP7_75t_R g1134 ( 
.A(n_1070),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_987),
.A2(n_1012),
.B1(n_1023),
.B2(n_999),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1033),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1024),
.B(n_997),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1007),
.B(n_1050),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1005),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_994),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1079),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1025),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1053),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1037),
.Y(n_1144)
);

CKINVDCx6p67_ASAP7_75t_R g1145 ( 
.A(n_1064),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1035),
.A2(n_1014),
.B(n_1036),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1072),
.A2(n_1003),
.B1(n_1081),
.B2(n_1079),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1015),
.B(n_1018),
.Y(n_1148)
);

AO21x1_ASAP7_75t_L g1149 ( 
.A1(n_997),
.A2(n_1031),
.B(n_1032),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1023),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_1017),
.B(n_1019),
.Y(n_1151)
);

BUFx2_ASAP7_75t_R g1152 ( 
.A(n_1074),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1056),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1021),
.A2(n_1076),
.B1(n_996),
.B2(n_1073),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1063),
.A2(n_1031),
.B(n_1020),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1028),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1038),
.A2(n_1071),
.B1(n_1041),
.B2(n_980),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_994),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1020),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_1025),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1041),
.A2(n_1084),
.B1(n_1052),
.B2(n_1016),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1008),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1080),
.A2(n_989),
.B1(n_1058),
.B2(n_1030),
.Y(n_1163)
);

AO21x1_ASAP7_75t_SL g1164 ( 
.A1(n_1052),
.A2(n_1084),
.B(n_1025),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1052),
.A2(n_1084),
.B1(n_1050),
.B2(n_1026),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1047),
.A2(n_863),
.B1(n_585),
.B2(n_1065),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1060),
.B(n_1000),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1060),
.A2(n_827),
.B1(n_842),
.B2(n_833),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1060),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_977),
.Y(n_1170)
);

INVx6_ASAP7_75t_L g1171 ( 
.A(n_1007),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1067),
.A2(n_585),
.B(n_448),
.Y(n_1172)
);

INVx6_ASAP7_75t_L g1173 ( 
.A(n_1007),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1064),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1034),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1000),
.B(n_1039),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_978),
.A2(n_827),
.B1(n_842),
.B2(n_833),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1017),
.B(n_1019),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_1049),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1085),
.B(n_974),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1000),
.B(n_1039),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1034),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_978),
.A2(n_827),
.B1(n_842),
.B2(n_833),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1065),
.A2(n_863),
.B1(n_585),
.B2(n_1045),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_1064),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_978),
.A2(n_827),
.B1(n_842),
.B2(n_833),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1127),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1127),
.B(n_1136),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1090),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1146),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1097),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1144),
.B(n_1097),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1097),
.B(n_1175),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1175),
.B(n_1182),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1172),
.A2(n_1092),
.B(n_1184),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1117),
.B(n_1126),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1104),
.Y(n_1197)
);

CKINVDCx11_ASAP7_75t_R g1198 ( 
.A(n_1099),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1109),
.B(n_1095),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1104),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1130),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1135),
.B(n_1110),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1110),
.A2(n_1186),
.B(n_1177),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1130),
.Y(n_1204)
);

AO21x1_ASAP7_75t_SL g1205 ( 
.A1(n_1114),
.A2(n_1150),
.B(n_1135),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1141),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1149),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1155),
.B(n_1159),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1118),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1120),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1120),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1101),
.Y(n_1213)
);

INVxp33_ASAP7_75t_SL g1214 ( 
.A(n_1107),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1117),
.B(n_1126),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1121),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1132),
.A2(n_1096),
.B(n_1166),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1137),
.A2(n_1186),
.B(n_1177),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1137),
.A2(n_1183),
.B(n_1103),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1183),
.A2(n_1094),
.B(n_1180),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1139),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1090),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1111),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1112),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1102),
.A2(n_1168),
.B(n_1115),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1091),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1090),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1099),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1148),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1170),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1128),
.B(n_1123),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1090),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1165),
.A2(n_1161),
.B(n_1138),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1105),
.B(n_1168),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1133),
.Y(n_1235)
);

AO21x1_ASAP7_75t_SL g1236 ( 
.A1(n_1165),
.A2(n_1161),
.B(n_1162),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1143),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1106),
.B(n_1151),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1129),
.B(n_1173),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1129),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1187),
.B(n_1088),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1188),
.B(n_1176),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1195),
.A2(n_1105),
.B1(n_1181),
.B2(n_1108),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1188),
.Y(n_1244)
);

NOR2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1222),
.B(n_1124),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1188),
.B(n_1167),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1189),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1201),
.B(n_1147),
.Y(n_1248)
);

NOR2x1_ASAP7_75t_SL g1249 ( 
.A(n_1217),
.B(n_1164),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1223),
.Y(n_1250)
);

NOR2x1_ASAP7_75t_L g1251 ( 
.A(n_1207),
.B(n_1129),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1208),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1195),
.A2(n_1116),
.B1(n_1156),
.B2(n_1154),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1201),
.B(n_1093),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1208),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1204),
.B(n_1098),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1204),
.B(n_1178),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1208),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1223),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1224),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1219),
.B(n_1190),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1219),
.B(n_1178),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1219),
.B(n_1178),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1219),
.B(n_1106),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1199),
.B(n_1153),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1219),
.B(n_1106),
.Y(n_1266)
);

OAI221xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1199),
.A2(n_1163),
.B1(n_1145),
.B2(n_1157),
.C(n_1153),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1197),
.B(n_1134),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1215),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1213),
.Y(n_1270)
);

OAI221xp5_ASAP7_75t_L g1271 ( 
.A1(n_1203),
.A2(n_1138),
.B1(n_1122),
.B2(n_1171),
.C(n_1173),
.Y(n_1271)
);

OAI221xp5_ASAP7_75t_L g1272 ( 
.A1(n_1253),
.A2(n_1220),
.B1(n_1203),
.B2(n_1243),
.C(n_1225),
.Y(n_1272)
);

OAI221xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1253),
.A2(n_1199),
.B1(n_1243),
.B2(n_1234),
.C(n_1202),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1262),
.B(n_1193),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1268),
.B(n_1225),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1262),
.B(n_1193),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1248),
.A2(n_1220),
.B(n_1202),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1254),
.B(n_1256),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1254),
.B(n_1229),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1267),
.A2(n_1218),
.B1(n_1265),
.B2(n_1202),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1261),
.A2(n_1197),
.B(n_1200),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1271),
.A2(n_1217),
.B(n_1218),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1254),
.B(n_1229),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1262),
.B(n_1194),
.Y(n_1285)
);

NAND3xp33_ASAP7_75t_L g1286 ( 
.A(n_1267),
.B(n_1234),
.C(n_1218),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1256),
.B(n_1206),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1256),
.B(n_1206),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1241),
.B(n_1210),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1265),
.A2(n_1218),
.B1(n_1156),
.B2(n_1235),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1241),
.B(n_1210),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1241),
.B(n_1221),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1241),
.B(n_1221),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1249),
.A2(n_1217),
.B1(n_1218),
.B2(n_1233),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1246),
.B(n_1216),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1268),
.B(n_1224),
.C(n_1216),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1246),
.B(n_1242),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1263),
.B(n_1194),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1268),
.B(n_1226),
.C(n_1230),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1271),
.A2(n_1237),
.B1(n_1235),
.B2(n_1152),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1246),
.B(n_1217),
.Y(n_1301)
);

AND4x1_ASAP7_75t_L g1302 ( 
.A(n_1251),
.B(n_1198),
.C(n_1232),
.D(n_1116),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1263),
.B(n_1208),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1263),
.B(n_1208),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1246),
.B(n_1209),
.Y(n_1305)
);

AOI221xp5_ASAP7_75t_L g1306 ( 
.A1(n_1248),
.A2(n_1237),
.B1(n_1231),
.B2(n_1230),
.C(n_1226),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1242),
.B(n_1268),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1251),
.B(n_1238),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1264),
.B(n_1191),
.Y(n_1309)
);

OAI221xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1271),
.A2(n_1209),
.B1(n_1145),
.B2(n_1239),
.C(n_1215),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1242),
.B(n_1209),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1248),
.A2(n_1205),
.B1(n_1236),
.B2(n_1196),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1248),
.A2(n_1214),
.B(n_1238),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_SL g1314 ( 
.A1(n_1249),
.A2(n_1239),
.B(n_1227),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1270),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1251),
.B(n_1232),
.C(n_1211),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1250),
.B(n_1212),
.C(n_1211),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1257),
.B(n_1192),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1315),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1303),
.B(n_1266),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1303),
.B(n_1266),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1304),
.B(n_1266),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1301),
.B(n_1311),
.Y(n_1323)
);

NAND2x1_ASAP7_75t_SL g1324 ( 
.A(n_1304),
.B(n_1255),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1274),
.B(n_1252),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1287),
.B(n_1250),
.Y(n_1326)
);

AND2x2_ASAP7_75t_SL g1327 ( 
.A(n_1302),
.B(n_1252),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1315),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1274),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1276),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1282),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1276),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1285),
.B(n_1252),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1278),
.B(n_1244),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1282),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1285),
.B(n_1261),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1282),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1279),
.B(n_1244),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1288),
.B(n_1259),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1305),
.B(n_1259),
.Y(n_1340)
);

AND3x1_ASAP7_75t_L g1341 ( 
.A(n_1277),
.B(n_1198),
.C(n_1228),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1298),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1309),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1297),
.B(n_1255),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1308),
.B(n_1258),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1294),
.B(n_1258),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1280),
.B(n_1260),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1292),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1293),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1317),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1282),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1316),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1289),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1291),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1341),
.A2(n_1272),
.B1(n_1286),
.B2(n_1300),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1329),
.B(n_1269),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1350),
.B(n_1307),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1350),
.B(n_1284),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1335),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1323),
.B(n_1295),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1332),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1335),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1335),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1332),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1319),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1319),
.Y(n_1366)
);

INVxp33_ASAP7_75t_L g1367 ( 
.A(n_1324),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1335),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1335),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1348),
.B(n_1275),
.Y(n_1370)
);

NOR2xp67_ASAP7_75t_L g1371 ( 
.A(n_1352),
.B(n_1296),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1348),
.B(n_1306),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1328),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1323),
.B(n_1318),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_L g1375 ( 
.A(n_1347),
.B(n_1283),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1352),
.B(n_1296),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1328),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1329),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1347),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1341),
.A2(n_1286),
.B1(n_1273),
.B2(n_1327),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1342),
.B(n_1269),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1326),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1343),
.B(n_1244),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1326),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1349),
.B(n_1257),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1339),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1349),
.B(n_1353),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1342),
.Y(n_1388)
);

NAND2x1_ASAP7_75t_L g1389 ( 
.A(n_1351),
.B(n_1314),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1339),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1320),
.B(n_1269),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1320),
.B(n_1269),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1365),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1388),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1357),
.B(n_1340),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1366),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1391),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1356),
.B(n_1327),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1371),
.B(n_1327),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1373),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1379),
.B(n_1353),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1378),
.B(n_1345),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1355),
.A2(n_1283),
.B1(n_1281),
.B2(n_1310),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1360),
.B(n_1340),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1377),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_L g1407 ( 
.A1(n_1375),
.A2(n_1346),
.B(n_1312),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1356),
.B(n_1325),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1382),
.B(n_1354),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1360),
.B(n_1354),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1380),
.B(n_1376),
.C(n_1372),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1384),
.B(n_1336),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1370),
.B(n_1228),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1381),
.B(n_1325),
.Y(n_1414)
);

OAI32xp33_ASAP7_75t_L g1415 ( 
.A1(n_1376),
.A2(n_1346),
.A3(n_1343),
.B1(n_1351),
.B2(n_1290),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1386),
.A2(n_1313),
.B1(n_1346),
.B2(n_1345),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1390),
.B(n_1124),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1381),
.B(n_1325),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1378),
.B(n_1345),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1361),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1364),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1387),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1383),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1383),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_1359),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1374),
.Y(n_1427)
);

OAI21xp33_ASAP7_75t_L g1428 ( 
.A1(n_1367),
.A2(n_1302),
.B(n_1314),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1389),
.Y(n_1429)
);

NAND2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1389),
.B(n_1247),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1374),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1367),
.B(n_1185),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1391),
.B(n_1333),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1392),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1362),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1393),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1432),
.B(n_1411),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1396),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1430),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1399),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1401),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1394),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1406),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1394),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1420),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1404),
.A2(n_1345),
.B1(n_1392),
.B2(n_1269),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1435),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1398),
.B(n_1320),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1417),
.Y(n_1449)
);

AOI222xp33_ASAP7_75t_L g1450 ( 
.A1(n_1407),
.A2(n_1331),
.B1(n_1299),
.B2(n_1249),
.C1(n_1345),
.C2(n_1351),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1399),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1435),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1421),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1413),
.B(n_1185),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1408),
.B(n_1321),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1403),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1404),
.A2(n_1331),
.B1(n_1258),
.B2(n_1351),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1400),
.B(n_1334),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1427),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1403),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1428),
.B(n_1359),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1431),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1413),
.B(n_1179),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1416),
.A2(n_1245),
.B1(n_1257),
.B2(n_1258),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1429),
.B(n_1359),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1419),
.B(n_1362),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1422),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1419),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1397),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1395),
.B(n_1334),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1415),
.B(n_1179),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1471),
.A2(n_1409),
.B(n_1402),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1471),
.A2(n_1425),
.B1(n_1429),
.B2(n_1351),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_1468),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1440),
.Y(n_1475)
);

NAND4xp25_ASAP7_75t_L g1476 ( 
.A(n_1437),
.B(n_1409),
.C(n_1402),
.D(n_1405),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1437),
.A2(n_1461),
.B(n_1444),
.C(n_1442),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1442),
.Y(n_1479)
);

OAI21xp33_ASAP7_75t_L g1480 ( 
.A1(n_1457),
.A2(n_1426),
.B(n_1434),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1451),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1447),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1458),
.B(n_1410),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1459),
.B(n_1414),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1454),
.B(n_1100),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1447),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1452),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1461),
.A2(n_1462),
.B1(n_1467),
.B2(n_1436),
.C(n_1453),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1449),
.A2(n_1425),
.B(n_1113),
.C(n_1089),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1452),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1438),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1441),
.B(n_1443),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1460),
.A2(n_1424),
.B1(n_1423),
.B2(n_1412),
.Y(n_1493)
);

OAI21xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1450),
.A2(n_1418),
.B(n_1412),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1445),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1446),
.A2(n_1430),
.B1(n_1330),
.B2(n_1433),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1469),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1475),
.B(n_1481),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1474),
.B(n_1478),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1488),
.B(n_1456),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1487),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1477),
.B(n_1469),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1477),
.B(n_1464),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1485),
.B(n_1454),
.Y(n_1504)
);

NAND2x1_ASAP7_75t_SL g1505 ( 
.A(n_1493),
.B(n_1439),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1479),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1482),
.B(n_1448),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1486),
.B(n_1463),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1490),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1484),
.B(n_1463),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1476),
.B(n_1439),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1473),
.B(n_1465),
.C(n_1439),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1483),
.B(n_1455),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1472),
.B(n_1497),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1473),
.A2(n_1465),
.B1(n_1466),
.B2(n_1205),
.Y(n_1515)
);

NAND4xp25_ASAP7_75t_L g1516 ( 
.A(n_1498),
.B(n_1492),
.C(n_1489),
.D(n_1491),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1502),
.A2(n_1494),
.B1(n_1496),
.B2(n_1495),
.Y(n_1517)
);

NOR3xp33_ASAP7_75t_L g1518 ( 
.A(n_1503),
.B(n_1489),
.C(n_1480),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1505),
.A2(n_1470),
.B1(n_1324),
.B2(n_1363),
.C(n_1369),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1513),
.B(n_1466),
.Y(n_1520)
);

AO22x1_ASAP7_75t_L g1521 ( 
.A1(n_1501),
.A2(n_1174),
.B1(n_1100),
.B2(n_1466),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1499),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1512),
.B(n_1174),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1511),
.A2(n_1369),
.B1(n_1368),
.B2(n_1363),
.Y(n_1524)
);

AND2x4_ASAP7_75t_SL g1525 ( 
.A(n_1510),
.B(n_1131),
.Y(n_1525)
);

NOR2x1_ASAP7_75t_L g1526 ( 
.A(n_1516),
.B(n_1504),
.Y(n_1526)
);

AND5x1_ASAP7_75t_L g1527 ( 
.A(n_1518),
.B(n_1511),
.C(n_1504),
.D(n_1500),
.E(n_1514),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1517),
.A2(n_1515),
.B1(n_1508),
.B2(n_1507),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1520),
.Y(n_1529)
);

NOR3xp33_ASAP7_75t_L g1530 ( 
.A(n_1523),
.B(n_1506),
.C(n_1509),
.Y(n_1530)
);

NOR4xp25_ASAP7_75t_L g1531 ( 
.A(n_1522),
.B(n_1515),
.C(n_1368),
.D(n_1363),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1525),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1521),
.B(n_1321),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1519),
.A2(n_1089),
.B(n_1113),
.C(n_1337),
.Y(n_1534)
);

NAND4xp75_ASAP7_75t_L g1535 ( 
.A(n_1526),
.B(n_1174),
.C(n_1524),
.D(n_1125),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1529),
.B(n_1344),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1527),
.A2(n_1239),
.B1(n_1337),
.B2(n_1330),
.C(n_1338),
.Y(n_1537)
);

NOR3xp33_ASAP7_75t_L g1538 ( 
.A(n_1532),
.B(n_1160),
.C(n_1142),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1528),
.B(n_1330),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1536),
.Y(n_1540)
);

NOR2x2_ASAP7_75t_L g1541 ( 
.A(n_1535),
.B(n_1530),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1539),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1538),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1537),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1539),
.A2(n_1533),
.B1(n_1531),
.B2(n_1245),
.Y(n_1545)
);

OAI311xp33_ASAP7_75t_L g1546 ( 
.A1(n_1545),
.A2(n_1534),
.A3(n_1299),
.B1(n_1338),
.C1(n_1322),
.Y(n_1546)
);

NOR2x1_ASAP7_75t_L g1547 ( 
.A(n_1542),
.B(n_1142),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1543),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1540),
.Y(n_1549)
);

NOR2xp67_ASAP7_75t_L g1550 ( 
.A(n_1541),
.B(n_1544),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1547),
.Y(n_1551)
);

XNOR2xp5_ASAP7_75t_L g1552 ( 
.A(n_1550),
.B(n_1245),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1548),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1553),
.Y(n_1554)
);

O2A1O1Ixp5_ASAP7_75t_L g1555 ( 
.A1(n_1554),
.A2(n_1549),
.B(n_1546),
.C(n_1552),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1555),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1555),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1556),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1557),
.A2(n_1554),
.B1(n_1551),
.B2(n_1169),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1559),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1558),
.A2(n_1169),
.B(n_1160),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1560),
.B(n_1344),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1562),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_R g1564 ( 
.A1(n_1563),
.A2(n_1561),
.B1(n_1173),
.B2(n_1171),
.C(n_1337),
.Y(n_1564)
);

AOI211xp5_ASAP7_75t_L g1565 ( 
.A1(n_1564),
.A2(n_1140),
.B(n_1158),
.C(n_1240),
.Y(n_1565)
);


endmodule