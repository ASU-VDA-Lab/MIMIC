module real_jpeg_12301_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_312, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_312;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_38),
.B1(n_44),
.B2(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_38),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_2),
.A2(n_38),
.B1(n_149),
.B2(n_150),
.Y(n_162)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_3),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_4),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_46),
.B1(n_101),
.B2(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_46),
.B1(n_149),
.B2(n_150),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_29),
.C(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_31),
.B1(n_44),
.B2(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_7),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_7),
.B(n_48),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_31),
.B1(n_101),
.B2(n_102),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_58),
.B(n_102),
.C(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_7),
.B(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_31),
.B1(n_149),
.B2(n_150),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_10),
.A2(n_44),
.B1(n_47),
.B2(n_155),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_10),
.A2(n_101),
.B1(n_102),
.B2(n_155),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_10),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.Y(n_286)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_304),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_296),
.B(n_303),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_258),
.B(n_293),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_239),
.B(n_257),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_218),
.B(n_238),
.Y(n_16)
);

AOI321xp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_178),
.A3(n_211),
.B1(n_216),
.B2(n_217),
.C(n_312),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_140),
.B(n_177),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_117),
.B(n_139),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_94),
.B(n_116),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_72),
.B(n_93),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_63),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_63),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_25),
.B(n_90),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_36),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_47),
.B(n_59),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_31),
.B(n_102),
.C(n_130),
.Y(n_148)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_33),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_33),
.A2(n_90),
.B(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_35),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_83),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_36),
.A2(n_154),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_51),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_42),
.B(n_69),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_42),
.A2(n_175),
.B(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_43),
.B(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_48),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_48),
.Y(n_176)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_51),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_52),
.Y(n_175)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_60),
.C(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_56),
.B(n_107),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_56),
.A2(n_104),
.B(n_107),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_56),
.A2(n_171),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_134),
.Y(n_133)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_59),
.B1(n_101),
.B2(n_102),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_71),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_86),
.B(n_92),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_80),
.B(n_85),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_84),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_82),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_110),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_108),
.C(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_102),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_103),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_105),
.B(n_134),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_105),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_109),
.A2(n_176),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_109),
.B(n_121),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_111),
.A2(n_112),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_111),
.A2(n_112),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_112),
.B(n_235),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_112),
.A2(n_246),
.B(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_138),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_138),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_137),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_123),
.C(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_126),
.B(n_145),
.C(n_157),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.CI(n_132),
.CON(n_126),
.SN(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_129),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_131),
.B1(n_149),
.B2(n_150),
.Y(n_166)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_133),
.B(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_133),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_157),
.B2(n_158),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_153),
.B2(n_156),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_168),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_170),
.C(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_163),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_164),
.A2(n_167),
.B(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_164),
.A2(n_182),
.B(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_165),
.B(n_183),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_171),
.B(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_173),
.A2(n_174),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_173),
.A2(n_174),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_174),
.B(n_266),
.C(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_174),
.B(n_290),
.C(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_205),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_205),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_190),
.C(n_201),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_185),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_182),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_186),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_198),
.C(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_194),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_197),
.A2(n_250),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_197),
.B(n_228),
.Y(n_306)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_198),
.A2(n_200),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_198),
.B(n_301),
.C(n_302),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_203),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.C(n_210),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_207),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_210),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_215),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_233),
.B2(n_234),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_234),
.C(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_226),
.C(n_231),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_230),
.B2(n_231),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_241),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_244),
.C(n_252),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_251),
.B2(n_252),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B(n_256),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_264),
.B1(n_265),
.B2(n_275),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_256),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_262),
.C(n_264),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_261),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_267),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_279),
.C(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_271),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_278),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_287),
.B1(n_288),
.B2(n_292),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);


endmodule