module fake_jpeg_1139_n_680 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_543;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_548;
wire n_266;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_16),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_61),
.Y(n_180)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_63),
.B(n_76),
.Y(n_152)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_65),
.B(n_96),
.Y(n_147)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_69),
.Y(n_195)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_20),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_71),
.A2(n_127),
.B1(n_32),
.B2(n_48),
.Y(n_173)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_85),
.B(n_87),
.Y(n_161)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_88),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_56),
.Y(n_93)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_94),
.Y(n_219)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_8),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_58),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_118),
.Y(n_167)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_40),
.Y(n_162)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_47),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_51),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_127)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_34),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_34),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_41),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_133),
.B(n_139),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_69),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g237 ( 
.A(n_140),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_63),
.B(n_40),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_162),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_73),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_165),
.B(n_166),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_61),
.B(n_52),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_48),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_197),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_173),
.A2(n_28),
.B1(n_35),
.B2(n_42),
.Y(n_250)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_93),
.Y(n_175)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

NAND3xp33_ASAP7_75t_SL g179 ( 
.A(n_104),
.B(n_30),
.C(n_32),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_28),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_66),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_187),
.A2(n_105),
.B1(n_62),
.B2(n_111),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_80),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_190),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_64),
.B(n_36),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_191),
.Y(n_291)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_129),
.B(n_24),
.Y(n_197)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_83),
.A2(n_91),
.B1(n_126),
.B2(n_125),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_203),
.A2(n_223),
.B1(n_164),
.B2(n_145),
.Y(n_299)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_205),
.Y(n_287)
);

INVx6_ASAP7_75t_SL g206 ( 
.A(n_78),
.Y(n_206)
);

CKINVDCx9p33_ASAP7_75t_R g259 ( 
.A(n_206),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_117),
.B(n_57),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_60),
.B(n_43),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_209),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_211),
.Y(n_303)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_88),
.Y(n_214)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_89),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_218),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_90),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_100),
.B(n_43),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_113),
.Y(n_249)
);

INVx6_ASAP7_75t_SL g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx9p33_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g315 ( 
.A(n_225),
.Y(n_315)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_227),
.Y(n_317)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_228),
.Y(n_333)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_229),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_167),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_230),
.B(n_251),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_152),
.A2(n_36),
.B1(n_42),
.B2(n_38),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_233),
.A2(n_246),
.B1(n_201),
.B2(n_176),
.Y(n_346)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_179),
.A2(n_128),
.B(n_103),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_239),
.A2(n_258),
.B(n_215),
.Y(n_320)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_131),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_243),
.A2(n_249),
.B(n_282),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_244),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_134),
.Y(n_245)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_245),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_250),
.A2(n_292),
.B1(n_299),
.B2(n_220),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_147),
.B(n_35),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_159),
.B(n_51),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_252),
.B(n_254),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_253),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_14),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_173),
.A2(n_123),
.B1(n_122),
.B2(n_112),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_255),
.A2(n_272),
.B1(n_290),
.B2(n_213),
.Y(n_351)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

CKINVDCx12_ASAP7_75t_R g257 ( 
.A(n_195),
.Y(n_257)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_257),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_184),
.A2(n_23),
.B(n_11),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx3_ASAP7_75t_SL g262 ( 
.A(n_212),
.Y(n_262)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_182),
.Y(n_263)
);

INVx11_ASAP7_75t_L g310 ( 
.A(n_263),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_188),
.B(n_106),
.Y(n_267)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_267),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_199),
.B(n_98),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_269),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_161),
.B(n_99),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_172),
.Y(n_270)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_146),
.Y(n_271)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_190),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_272)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_178),
.Y(n_274)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_6),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_276),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_163),
.B(n_137),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_277),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_180),
.B(n_0),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_278),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_178),
.Y(n_279)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_279),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_136),
.B(n_10),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_286),
.Y(n_314)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_150),
.Y(n_281)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_180),
.B(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_143),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_138),
.Y(n_285)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_144),
.B(n_157),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_215),
.B(n_10),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_294),
.Y(n_332)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_148),
.Y(n_289)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_160),
.A2(n_203),
.B1(n_219),
.B2(n_135),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_155),
.B(n_10),
.Y(n_294)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_182),
.Y(n_296)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_200),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_156),
.Y(n_301)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_174),
.B(n_11),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_194),
.Y(n_355)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_132),
.Y(n_354)
);

OAI21xp33_ASAP7_75t_L g394 ( 
.A1(n_320),
.A2(n_355),
.B(n_364),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_235),
.B(n_195),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_151),
.C(n_183),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_340),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_250),
.A2(n_150),
.B1(n_185),
.B2(n_220),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_336),
.B1(n_351),
.B2(n_360),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_258),
.A2(n_153),
.B(n_181),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_335),
.B(n_260),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_278),
.B(n_181),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_345),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_237),
.Y(n_340)
);

OA22x2_ASAP7_75t_L g342 ( 
.A1(n_255),
.A2(n_164),
.B1(n_145),
.B2(n_132),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_SL g397 ( 
.A1(n_342),
.A2(n_260),
.B(n_303),
.C(n_225),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_241),
.B(n_169),
.C(n_182),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_361),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_278),
.B(n_223),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_346),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_239),
.A2(n_213),
.B1(n_194),
.B2(n_198),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_357),
.B1(n_336),
.B2(n_246),
.Y(n_384)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

AOI22x1_ASAP7_75t_L g357 ( 
.A1(n_243),
.A2(n_169),
.B1(n_135),
.B2(n_221),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_240),
.B(n_201),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_364),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_290),
.A2(n_192),
.B1(n_186),
.B2(n_149),
.Y(n_360)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_232),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_282),
.B(n_201),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_259),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_370),
.B(n_391),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_243),
.B1(n_292),
.B2(n_231),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_372),
.A2(n_386),
.B1(n_406),
.B2(n_354),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_309),
.B(n_272),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_373),
.B(n_392),
.Y(n_416)
);

NOR2x1_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_335),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_374),
.A2(n_313),
.B(n_362),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_349),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_376),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_333),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_326),
.B(n_229),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_378),
.B(n_388),
.Y(n_426)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_308),
.Y(n_383)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_384),
.A2(n_397),
.B1(n_402),
.B2(n_405),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_320),
.A2(n_355),
.B1(n_357),
.B2(n_345),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_385),
.A2(n_393),
.B1(n_407),
.B2(n_412),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_311),
.A2(n_264),
.B1(n_246),
.B2(n_304),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_306),
.Y(n_387)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_328),
.B(n_282),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_310),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_305),
.B(n_334),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_396),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_307),
.B(n_259),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_314),
.B(n_237),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_343),
.A2(n_246),
.B1(n_192),
.B2(n_186),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_410),
.B(n_413),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_305),
.B(n_312),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_338),
.B(n_297),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_398),
.B(n_401),
.Y(n_443)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_297),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_403),
.A2(n_352),
.B(n_296),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_329),
.B(n_228),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_316),
.Y(n_444)
);

INVx11_ASAP7_75t_L g405 ( 
.A(n_310),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_360),
.A2(n_262),
.B1(n_295),
.B2(n_287),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_342),
.A2(n_242),
.B1(n_274),
.B2(n_279),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_408),
.B(n_409),
.Y(n_420)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_344),
.A2(n_303),
.B(n_293),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_333),
.Y(n_411)
);

INVx13_ASAP7_75t_L g415 ( 
.A(n_411),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_342),
.A2(n_354),
.B1(n_359),
.B2(n_339),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_353),
.A2(n_352),
.B(n_317),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_414),
.A2(n_374),
.B(n_371),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_390),
.Y(n_418)
);

INVx13_ASAP7_75t_L g471 ( 
.A(n_418),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_388),
.B(n_398),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_422),
.B(n_432),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_385),
.A2(n_342),
.B1(n_356),
.B2(n_321),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_428),
.A2(n_436),
.B1(n_383),
.B2(n_387),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_439),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_322),
.C(n_318),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_434),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_413),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_319),
.C(n_324),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_384),
.A2(n_356),
.B1(n_321),
.B2(n_315),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_353),
.C(n_316),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_438),
.B(n_449),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_392),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_368),
.A2(n_323),
.B1(n_350),
.B2(n_298),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_440),
.A2(n_446),
.B1(n_452),
.B2(n_406),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_378),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_381),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_444),
.B(n_453),
.Y(n_470)
);

OAI22x1_ASAP7_75t_L g446 ( 
.A1(n_395),
.A2(n_289),
.B1(n_227),
.B2(n_317),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_367),
.B(n_362),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_448),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_367),
.B(n_337),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_377),
.B(n_295),
.C(n_284),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_450),
.A2(n_414),
.B(n_403),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_380),
.B(n_337),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_454),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_368),
.A2(n_323),
.B1(n_350),
.B2(n_244),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_373),
.B(n_348),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_325),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_456),
.B(n_467),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_432),
.A2(n_395),
.B1(n_393),
.B2(n_407),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_457),
.A2(n_480),
.B1(n_426),
.B2(n_449),
.Y(n_504)
);

AOI32xp33_ASAP7_75t_L g459 ( 
.A1(n_445),
.A2(n_377),
.A3(n_370),
.B1(n_396),
.B2(n_391),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_459),
.B(n_488),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_425),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_460),
.A2(n_463),
.B1(n_468),
.B2(n_469),
.Y(n_505)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_461),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_425),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_462),
.B(n_473),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_424),
.Y(n_463)
);

HAxp5_ASAP7_75t_SL g464 ( 
.A(n_427),
.B(n_374),
.CON(n_464),
.SN(n_464)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_416),
.C(n_426),
.Y(n_498)
);

INVx8_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_465),
.Y(n_509)
);

OA22x2_ASAP7_75t_L g467 ( 
.A1(n_437),
.A2(n_386),
.B1(n_397),
.B2(n_372),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_424),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_420),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_454),
.Y(n_472)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_375),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_476),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_SL g475 ( 
.A(n_430),
.B(n_412),
.C(n_410),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_475),
.B(n_429),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_401),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_421),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_419),
.Y(n_479)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_479),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_403),
.Y(n_482)
);

AND2x2_ASAP7_75t_SL g511 ( 
.A(n_482),
.B(n_423),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

AO22x1_ASAP7_75t_L g485 ( 
.A1(n_450),
.A2(n_397),
.B1(n_371),
.B2(n_405),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_490),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_487),
.A2(n_441),
.B1(n_417),
.B2(n_428),
.Y(n_495)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_489),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_443),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_447),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_431),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_495),
.A2(n_500),
.B1(n_507),
.B2(n_477),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_473),
.B(n_431),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_496),
.B(n_421),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_498),
.B(n_489),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_456),
.A2(n_446),
.B(n_417),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_499),
.A2(n_484),
.B(n_482),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_466),
.A2(n_452),
.B1(n_440),
.B2(n_436),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_501),
.B(n_510),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_438),
.C(n_434),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_528),
.C(n_462),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_504),
.A2(n_460),
.B1(n_487),
.B2(n_481),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_465),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_506),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_466),
.A2(n_416),
.B1(n_443),
.B2(n_422),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_476),
.B(n_409),
.Y(n_510)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_463),
.B(n_408),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_512),
.B(n_520),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_483),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_514),
.B(n_470),
.Y(n_531)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_516),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_469),
.B(n_429),
.Y(n_519)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_519),
.Y(n_542)
);

NOR4xp25_ASAP7_75t_L g522 ( 
.A(n_461),
.B(n_423),
.C(n_399),
.D(n_433),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_522),
.B(n_524),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_466),
.B(n_446),
.Y(n_523)
);

XNOR2x1_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_366),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_478),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_433),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_526),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_482),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_527),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_475),
.B(n_400),
.C(n_402),
.Y(n_528)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_530),
.B(n_545),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_531),
.B(n_543),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_478),
.C(n_468),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_560),
.C(n_511),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_495),
.A2(n_472),
.B1(n_491),
.B2(n_481),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_534),
.A2(n_535),
.B1(n_540),
.B2(n_546),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_494),
.Y(n_537)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_537),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_515),
.A2(n_490),
.B(n_455),
.C(n_458),
.Y(n_539)
);

AOI21xp33_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_541),
.B(n_547),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_492),
.A2(n_458),
.B1(n_455),
.B2(n_474),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_471),
.B(n_467),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_467),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_519),
.Y(n_544)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_544),
.Y(n_567)
);

XNOR2x2_ASAP7_75t_SL g545 ( 
.A(n_516),
.B(n_471),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_492),
.A2(n_480),
.B1(n_467),
.B2(n_479),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_550),
.A2(n_499),
.B1(n_515),
.B2(n_526),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_525),
.A2(n_411),
.B(n_376),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_555),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_517),
.B(n_369),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_552),
.B(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_502),
.Y(n_554)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_554),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_556),
.B(n_509),
.Y(n_585)
);

XOR2x2_ASAP7_75t_L g558 ( 
.A(n_507),
.B(n_415),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_558),
.B(n_509),
.Y(n_582)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_508),
.Y(n_559)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_559),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_528),
.B(n_497),
.C(n_511),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_562),
.A2(n_588),
.B1(n_532),
.B2(n_536),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_554),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_550),
.A2(n_513),
.B1(n_526),
.B2(n_493),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_565),
.A2(n_576),
.B1(n_578),
.B2(n_585),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_530),
.B(n_513),
.C(n_493),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_566),
.B(n_572),
.Y(n_603)
);

FAx1_ASAP7_75t_SL g572 ( 
.A(n_561),
.B(n_496),
.CI(n_527),
.CON(n_572),
.SN(n_572)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_540),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_575),
.A2(n_577),
.B1(n_586),
.B2(n_587),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_546),
.A2(n_513),
.B1(n_527),
.B2(n_497),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_559),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_534),
.A2(n_500),
.B1(n_506),
.B2(n_523),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_521),
.C(n_518),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_580),
.C(n_558),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_531),
.B(n_521),
.C(n_509),
.Y(n_580)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_560),
.Y(n_591)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_537),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_535),
.A2(n_435),
.B1(n_415),
.B2(n_366),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_SL g589 ( 
.A(n_570),
.B(n_543),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_589),
.B(n_592),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_591),
.B(n_607),
.Y(n_625)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_593),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_SL g615 ( 
.A(n_594),
.B(n_600),
.Y(n_615)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_574),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_595),
.B(n_596),
.Y(n_627)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_568),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_584),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_597),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_588),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_598),
.B(n_601),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_580),
.B(n_556),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_599),
.B(n_602),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_549),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_564),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_541),
.Y(n_602)
);

INVx13_ASAP7_75t_L g604 ( 
.A(n_572),
.Y(n_604)
);

INVx11_ASAP7_75t_L g621 ( 
.A(n_604),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_553),
.C(n_538),
.Y(n_605)
);

BUFx24_ASAP7_75t_SL g616 ( 
.A(n_605),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_569),
.A2(n_551),
.B(n_536),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_608),
.C(n_611),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_583),
.B(n_555),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_SL g608 ( 
.A(n_570),
.B(n_538),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_SL g611 ( 
.A(n_566),
.B(n_529),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_590),
.A2(n_571),
.B1(n_532),
.B2(n_561),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_612),
.A2(n_363),
.B1(n_330),
.B2(n_273),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_591),
.B(n_582),
.C(n_565),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_613),
.B(n_618),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_603),
.A2(n_544),
.B(n_542),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_617),
.A2(n_624),
.B(n_389),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_597),
.A2(n_571),
.B1(n_567),
.B2(n_542),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_600),
.A2(n_572),
.B1(n_545),
.B2(n_578),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_620),
.B(n_630),
.Y(n_646)
);

NOR3xp33_ASAP7_75t_SL g622 ( 
.A(n_604),
.B(n_539),
.C(n_576),
.Y(n_622)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_622),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_602),
.A2(n_573),
.B(n_562),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_611),
.A2(n_548),
.B1(n_573),
.B2(n_435),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_629),
.B(n_610),
.Y(n_631)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_631),
.A2(n_638),
.B(n_639),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_613),
.B(n_594),
.C(n_592),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_633),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_627),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_623),
.B(n_599),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_634),
.B(n_640),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_609),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_636),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_L g637 ( 
.A1(n_616),
.A2(n_593),
.B1(n_608),
.B2(n_548),
.C(n_589),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_637),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_614),
.B(n_607),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_615),
.B(n_415),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_628),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_643),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_628),
.B(n_325),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_619),
.B(n_348),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_644),
.A2(n_626),
.B(n_625),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_645),
.B(n_330),
.C(n_363),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_635),
.A2(n_617),
.B(n_612),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_648),
.B(n_655),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_649),
.B(n_657),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_654),
.A2(n_650),
.B1(n_651),
.B2(n_647),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_641),
.A2(n_621),
.B(n_622),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_632),
.B(n_636),
.C(n_634),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_631),
.B(n_625),
.C(n_621),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_658),
.B(n_653),
.Y(n_666)
);

AOI322xp5_ASAP7_75t_L g659 ( 
.A1(n_652),
.A2(n_646),
.A3(n_640),
.B1(n_638),
.B2(n_642),
.C1(n_645),
.C2(n_271),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_659),
.B(n_660),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_651),
.A2(n_245),
.B1(n_248),
.B2(n_281),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_661),
.B(n_663),
.Y(n_670)
);

AOI322xp5_ASAP7_75t_L g663 ( 
.A1(n_652),
.A2(n_221),
.A3(n_365),
.B1(n_176),
.B2(n_198),
.C1(n_263),
.C2(n_265),
.Y(n_663)
);

AOI322xp5_ASAP7_75t_L g665 ( 
.A1(n_656),
.A2(n_221),
.A3(n_365),
.B1(n_265),
.B2(n_287),
.C1(n_284),
.C2(n_234),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_665),
.B(n_666),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g668 ( 
.A1(n_662),
.A2(n_291),
.B(n_238),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_668),
.B(n_671),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_664),
.A2(n_234),
.B(n_266),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_SL g672 ( 
.A1(n_667),
.A2(n_660),
.B(n_266),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_672),
.A2(n_5),
.B(n_18),
.Y(n_675)
);

AOI322xp5_ASAP7_75t_L g674 ( 
.A1(n_669),
.A2(n_670),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_13),
.C2(n_15),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_674),
.B(n_18),
.C(n_5),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_675),
.B(n_676),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_677),
.A2(n_673),
.B1(n_18),
.B2(n_1),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_18),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_SL g680 ( 
.A(n_679),
.B(n_1),
.C(n_677),
.Y(n_680)
);


endmodule