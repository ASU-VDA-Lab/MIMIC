module fake_jpeg_27422_n_344 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_68),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2x1_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_33),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_36),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_51),
.B1(n_27),
.B2(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_87),
.B1(n_33),
.B2(n_32),
.Y(n_131)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_51),
.B1(n_27),
.B2(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_98),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_48),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_94),
.B(n_47),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_23),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_99),
.Y(n_106)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_28),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_101),
.Y(n_132)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_65),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_112),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_45),
.B(n_48),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_124),
.B(n_127),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_27),
.B1(n_57),
.B2(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_114),
.B1(n_117),
.B2(n_85),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_21),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_61),
.B1(n_69),
.B2(n_54),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

XNOR2x2_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_23),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_25),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_66),
.B1(n_41),
.B2(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_130),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_47),
.B(n_46),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_46),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_55),
.B1(n_41),
.B2(n_32),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_77),
.B1(n_97),
.B2(n_99),
.Y(n_141)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_131),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_142),
.Y(n_163)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_146),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_84),
.B(n_75),
.C(n_93),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_109),
.B(n_106),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_153),
.C(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_112),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_148),
.Y(n_173)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_152),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_90),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_156),
.Y(n_178)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_105),
.A2(n_98),
.B1(n_77),
.B2(n_83),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_114),
.B1(n_123),
.B2(n_106),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_83),
.B1(n_21),
.B2(n_26),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_132),
.B1(n_25),
.B2(n_2),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_74),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_17),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_25),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_101),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_111),
.B(n_126),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_160),
.A2(n_172),
.B(n_175),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_186),
.B(n_149),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_168),
.B1(n_170),
.B2(n_185),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_132),
.B1(n_130),
.B2(n_125),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_132),
.B1(n_125),
.B2(n_110),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_184),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_133),
.B(n_128),
.C(n_26),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_121),
.B(n_119),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_183),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_158),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_46),
.C(n_43),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_136),
.C(n_147),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_101),
.B1(n_70),
.B2(n_82),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_96),
.B(n_107),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_193),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_207),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_147),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_143),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_163),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_146),
.B1(n_135),
.B2(n_152),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_135),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_189),
.B(n_212),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_43),
.C(n_107),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_43),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_37),
.A3(n_31),
.B1(n_20),
.B2(n_19),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_215),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_19),
.B1(n_37),
.B2(n_31),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_214),
.A2(n_167),
.B1(n_182),
.B2(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_96),
.B1(n_24),
.B2(n_29),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_174),
.B1(n_185),
.B2(n_184),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_237),
.B1(n_195),
.B2(n_214),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_181),
.CI(n_163),
.CON(n_224),
.SN(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_175),
.B(n_167),
.C(n_2),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_230),
.B(n_212),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_37),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_96),
.B1(n_20),
.B2(n_24),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_24),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_30),
.Y(n_261)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_199),
.Y(n_251)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_234),
.A2(n_195),
.B(n_198),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_263),
.B(n_230),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_197),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_239),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_209),
.C(n_193),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_228),
.C(n_238),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_217),
.B1(n_226),
.B2(n_240),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_210),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_0),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_262),
.B1(n_265),
.B2(n_237),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_239),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

HAxp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_30),
.CON(n_263),
.SN(n_263)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_279),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_269),
.A2(n_247),
.B1(n_246),
.B2(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_274),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_220),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_277),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_224),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_254),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_261),
.C(n_263),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_218),
.C(n_225),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_258),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_243),
.C(n_219),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_251),
.C(n_219),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_250),
.B(n_224),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_275),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_294),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_247),
.B1(n_257),
.B2(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_298),
.B1(n_280),
.B2(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_227),
.Y(n_294)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_4),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_283),
.A2(n_252),
.B1(n_262),
.B2(n_259),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_29),
.C(n_28),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_277),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_303),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_304),
.B(n_308),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_271),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_313),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_312),
.B1(n_311),
.B2(n_7),
.Y(n_323)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_307),
.B1(n_302),
.B2(n_299),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_284),
.B(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_295),
.B(n_291),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_296),
.C(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_6),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_300),
.B1(n_303),
.B2(n_306),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_328),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_315),
.A2(n_319),
.B1(n_318),
.B2(n_317),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_325),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_326),
.B(n_316),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_8),
.C(n_11),
.Y(n_336)
);

AOI322xp5_ASAP7_75t_L g339 ( 
.A1(n_337),
.A2(n_335),
.A3(n_336),
.B1(n_327),
.B2(n_324),
.C1(n_12),
.C2(n_15),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_336),
.B(n_14),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_13),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_341),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_338),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_15),
.C(n_16),
.Y(n_344)
);


endmodule