module real_jpeg_33993_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_0),
.Y(n_120)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_1),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_1),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_1),
.B(n_177),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_1),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_1),
.B(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_2),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_4),
.Y(n_117)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_5),
.Y(n_127)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_5),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_6),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_6),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_6),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_6),
.B(n_93),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_6),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_7),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_7),
.B(n_77),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_8),
.B(n_126),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_8),
.B(n_114),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_8),
.B(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_11),
.Y(n_325)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_12),
.B(n_33),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_L g149 ( 
.A(n_12),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_12),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_12),
.B(n_272),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_12),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_12),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_13),
.B(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_14),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_14),
.B(n_39),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_14),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_14),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_14),
.B(n_93),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_15),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_202),
.Y(n_201)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_16),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_16),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_16),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_16),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_16),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_16),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_17),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_212),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_160),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.C(n_136),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_21),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_69),
.B2(n_70),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_50),
.B2(n_51),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_24),
.Y(n_164)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_30),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_31),
.B(n_35),
.C(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.C(n_47),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_40),
.Y(n_274)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_42),
.B(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_48),
.Y(n_203)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_49),
.Y(n_278)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_51),
.B(n_69),
.C(n_164),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_53),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_58),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_60),
.B(n_65),
.Y(n_183)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_61),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_65),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_68),
.Y(n_172)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_85),
.C(n_96),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_71),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_74),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_76),
.A2(n_83),
.B(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_80),
.A2(n_82),
.B(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_85),
.A2(n_96),
.B1(n_97),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_85),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_234)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_95),
.Y(n_331)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_102),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_103),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_104),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_108),
.B(n_137),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_122),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_109),
.B(n_112),
.Y(n_217)
);

OA21x2_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_118),
.B(n_121),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_118),
.Y(n_121)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_154),
.B1(n_155),
.B2(n_159),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_122),
.B(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.C(n_132),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_123),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_249)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_127),
.Y(n_257)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_127),
.Y(n_285)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_262)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_153),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_148),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_139),
.B(n_148),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_SL g205 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_205)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_159),
.C(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_196),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_179),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_184),
.B1(n_194),
.B2(n_195),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_210),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_208),
.B2(n_209),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_204),
.Y(n_206)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_241),
.B(n_348),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_239),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_215),
.B(n_239),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_235),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_236),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.C(n_234),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_230),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_223),
.B(n_230),
.Y(n_297)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_226),
.B(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_265),
.B(n_347),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_263),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_245),
.B(n_263),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.C(n_261),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_246),
.B(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_248),
.B(n_261),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.C(n_254),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_250),
.Y(n_291)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

AO22x1_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_342),
.B(n_346),
.Y(n_265)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_299),
.B(n_341),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_288),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_288),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_281),
.C(n_287),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_269),
.A2(n_270),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_275),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_294),
.C(n_295),
.Y(n_293)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_282),
.B1(n_287),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_286),
.Y(n_317)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_287),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_298),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_293),
.C(n_296),
.Y(n_343)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_292),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_334),
.B(n_340),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_318),
.B(n_333),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_310),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_302),
.B(n_310),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_307),
.Y(n_326)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_317),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_316),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_316),
.C(n_317),
.Y(n_335)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_327),
.B(n_332),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_326),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_344),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);


endmodule