module fake_jpeg_4245_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_30),
.Y(n_65)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_17),
.B1(n_36),
.B2(n_25),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_57),
.B1(n_66),
.B2(n_69),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_58),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_45),
.B1(n_44),
.B2(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_24),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_72),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_79),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_83),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_87),
.Y(n_103)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_34),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_97),
.Y(n_127)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_63),
.B1(n_61),
.B2(n_55),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_40),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_43),
.Y(n_150)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_111),
.Y(n_143)
);

AND2x4_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_41),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_126),
.B(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_67),
.B1(n_53),
.B2(n_48),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_82),
.B1(n_90),
.B2(n_99),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_37),
.B(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_123),
.Y(n_131)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_124),
.B1(n_128),
.B2(n_82),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_54),
.B(n_37),
.C(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_107),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_135),
.B1(n_140),
.B2(n_148),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_151),
.B1(n_119),
.B2(n_124),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_79),
.B1(n_89),
.B2(n_70),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_136),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_76),
.B1(n_87),
.B2(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_147),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_74),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_78),
.B1(n_72),
.B2(n_84),
.Y(n_148)
);

CKINVDCx6p67_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_47),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_99),
.B1(n_62),
.B2(n_41),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_47),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_62),
.B1(n_43),
.B2(n_77),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_62),
.B1(n_77),
.B2(n_22),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_104),
.B1(n_106),
.B2(n_112),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_24),
.B1(n_30),
.B2(n_35),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_106),
.B(n_35),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_163),
.B(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_174),
.C(n_146),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_116),
.B1(n_123),
.B2(n_103),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_189),
.B(n_31),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_111),
.C(n_116),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_126),
.A3(n_121),
.B1(n_36),
.B2(n_27),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_127),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_186),
.B1(n_191),
.B2(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_139),
.A2(n_128),
.B1(n_119),
.B2(n_27),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_31),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_199),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_197),
.A2(n_202),
.B1(n_217),
.B2(n_218),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_132),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_201),
.C(n_206),
.Y(n_225)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_150),
.B1(n_137),
.B2(n_129),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_131),
.B1(n_158),
.B2(n_155),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_221),
.B1(n_191),
.B2(n_187),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_157),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_214),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_47),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_219),
.C(n_220),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_153),
.B1(n_102),
.B2(n_96),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_102),
.B1(n_96),
.B2(n_36),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_142),
.C(n_31),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_31),
.C(n_23),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_224),
.B(n_228),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_160),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_234),
.C(n_239),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_160),
.B(n_181),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_26),
.B(n_23),
.Y(n_270)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

AOI22x1_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_176),
.B1(n_191),
.B2(n_190),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_245),
.B(n_243),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_233),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_195),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_163),
.C(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_237),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_218),
.B(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_189),
.C(n_168),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_188),
.B1(n_169),
.B2(n_167),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_205),
.B1(n_203),
.B2(n_199),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_165),
.C(n_178),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_246),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_207),
.A2(n_188),
.B(n_164),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_220),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_192),
.C(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_171),
.Y(n_248)
);

XOR2x1_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_212),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_255),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_263),
.B(n_10),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_246),
.B(n_229),
.C(n_2),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_270),
.B1(n_254),
.B2(n_262),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_194),
.B1(n_193),
.B2(n_200),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_254),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_285)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_216),
.B1(n_33),
.B2(n_27),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_261),
.B1(n_268),
.B2(n_230),
.Y(n_274)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_33),
.B1(n_23),
.B2(n_26),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_236),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_270),
.B(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_272),
.B(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_263),
.B(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_225),
.C(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_276),
.C(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_225),
.C(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_12),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_259),
.B1(n_250),
.B2(n_266),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_285),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_256),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_291),
.C(n_295),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_252),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_275),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_256),
.C(n_4),
.Y(n_291)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_11),
.C(n_6),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_11),
.B(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_272),
.B(n_11),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_16),
.C(n_6),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_15),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_10),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_302),
.B1(n_278),
.B2(n_284),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_305),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_287),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_309),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_279),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_294),
.B(n_291),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_288),
.A2(n_275),
.B1(n_283),
.B2(n_279),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_274),
.B1(n_0),
.B2(n_8),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_297),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_315)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_298),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_318),
.A2(n_320),
.B(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_290),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_289),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_312),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_313),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_328),
.B(n_330),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_331),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_312),
.C(n_8),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_7),
.B(n_12),
.Y(n_329)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_7),
.Y(n_330)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_316),
.A2(n_13),
.B(n_14),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_330),
.B(n_326),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_317),
.B(n_334),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_333),
.B(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_322),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_15),
.Y(n_340)
);


endmodule