module real_aes_1515_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_832, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_831, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_832;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_831;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_503;
wire n_357;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_782;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_754;
wire n_607;
wire n_417;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_0), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_1), .B(n_644), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_2), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_3), .B(n_695), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_4), .A2(n_241), .B1(n_446), .B2(n_447), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_5), .A2(n_261), .B1(n_408), .B2(n_412), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_6), .A2(n_138), .B1(n_433), .B2(n_434), .Y(n_432) );
AO22x2_ASAP7_75t_L g324 ( .A1(n_7), .A2(n_196), .B1(n_314), .B2(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g758 ( .A(n_7), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_8), .A2(n_129), .B1(n_436), .B2(n_437), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_9), .A2(n_252), .B1(n_395), .B2(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_10), .A2(n_14), .B1(n_631), .B2(n_671), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_11), .A2(n_245), .B1(n_621), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_12), .A2(n_270), .B1(n_444), .B2(n_462), .Y(n_563) );
AO22x1_ASAP7_75t_L g628 ( .A1(n_13), .A2(n_202), .B1(n_629), .B2(n_631), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_15), .A2(n_74), .B1(n_441), .B2(n_447), .Y(n_464) );
OA22x2_ASAP7_75t_L g465 ( .A1(n_16), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_16), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_17), .A2(n_199), .B1(n_358), .B2(n_359), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_18), .A2(n_28), .B1(n_441), .B2(n_444), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_19), .A2(n_100), .B1(n_446), .B2(n_447), .Y(n_445) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_20), .A2(n_73), .B1(n_314), .B2(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_20), .B(n_757), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_21), .A2(n_54), .B1(n_444), .B2(n_446), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_22), .A2(n_159), .B1(n_441), .B2(n_447), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_23), .A2(n_177), .B1(n_364), .B2(n_403), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_24), .A2(n_51), .B1(n_395), .B2(n_396), .Y(n_394) );
AO222x2_ASAP7_75t_SL g497 ( .A1(n_25), .A2(n_155), .B1(n_269), .B2(n_332), .C1(n_388), .C2(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_26), .A2(n_214), .B1(n_358), .B2(n_359), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_27), .A2(n_70), .B1(n_362), .B2(n_364), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_29), .A2(n_143), .B1(n_592), .B2(n_594), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_30), .A2(n_284), .B1(n_362), .B2(n_364), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_31), .A2(n_174), .B1(n_412), .B2(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_32), .A2(n_154), .B1(n_677), .B2(n_807), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_33), .A2(n_68), .B1(n_440), .B2(n_462), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g470 ( .A1(n_34), .A2(n_239), .B1(n_277), .B2(n_428), .C1(n_471), .C2(n_472), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_35), .A2(n_183), .B1(n_364), .B2(n_538), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_36), .A2(n_217), .B1(n_358), .B2(n_359), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_37), .A2(n_90), .B1(n_635), .B2(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_38), .A2(n_246), .B1(n_444), .B2(n_446), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_39), .A2(n_250), .B1(n_408), .B2(n_412), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_40), .A2(n_121), .B1(n_446), .B2(n_447), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_41), .A2(n_170), .B1(n_338), .B2(n_342), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_42), .A2(n_194), .B1(n_362), .B2(n_419), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_43), .A2(n_45), .B1(n_491), .B2(n_625), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_44), .A2(n_115), .B1(n_434), .B2(n_472), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_46), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_47), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_48), .A2(n_186), .B1(n_436), .B2(n_437), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g745 ( .A1(n_49), .A2(n_57), .B1(n_513), .B2(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_50), .A2(n_267), .B1(n_416), .B2(n_418), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_52), .A2(n_151), .B1(n_604), .B2(n_605), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_53), .A2(n_107), .B1(n_368), .B2(n_371), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_55), .B(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_56), .A2(n_281), .B1(n_430), .B2(n_476), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_58), .A2(n_92), .B1(n_390), .B2(n_392), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_59), .A2(n_203), .B1(n_662), .B2(n_664), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_60), .A2(n_171), .B1(n_390), .B2(n_613), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_61), .A2(n_219), .B1(n_440), .B2(n_441), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_62), .A2(n_110), .B1(n_648), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_63), .A2(n_220), .B1(n_496), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_64), .A2(n_153), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_65), .A2(n_78), .B1(n_414), .B2(n_505), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_66), .A2(n_137), .B1(n_378), .B2(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_67), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_69), .A2(n_135), .B1(n_406), .B2(n_440), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_71), .A2(n_88), .B1(n_430), .B2(n_431), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_72), .A2(n_114), .B1(n_433), .B2(n_434), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_75), .A2(n_104), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_76), .A2(n_280), .B1(n_358), .B2(n_359), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_77), .A2(n_263), .B1(n_430), .B2(n_431), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_79), .A2(n_287), .B1(n_297), .B2(n_760), .C(n_763), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_80), .A2(n_167), .B1(n_506), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_81), .A2(n_108), .B1(n_347), .B2(n_351), .Y(n_346) );
INVx3_ASAP7_75t_L g314 ( .A(n_82), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_83), .A2(n_283), .B1(n_491), .B2(n_493), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_84), .A2(n_127), .B1(n_365), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_85), .A2(n_119), .B1(n_640), .B2(n_641), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_86), .A2(n_161), .B1(n_351), .B2(n_391), .Y(n_690) );
AO22x2_ASAP7_75t_L g687 ( .A1(n_87), .A2(n_688), .B1(n_702), .B2(n_703), .Y(n_687) );
INVx1_ASAP7_75t_L g702 ( .A(n_87), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_89), .A2(n_140), .B1(n_505), .B2(n_506), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_91), .A2(n_215), .B1(n_391), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_93), .A2(n_182), .B1(n_440), .B2(n_462), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_94), .B(n_622), .Y(n_728) );
XOR2x2_ASAP7_75t_L g424 ( .A(n_95), .B(n_425), .Y(n_424) );
OA22x2_ASAP7_75t_L g582 ( .A1(n_96), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_96), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_97), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_98), .A2(n_218), .B1(n_430), .B2(n_431), .Y(n_429) );
OA22x2_ASAP7_75t_L g800 ( .A1(n_99), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_99), .Y(n_801) );
INVx1_ASAP7_75t_SL g315 ( .A(n_101), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_101), .B(n_130), .Y(n_759) );
INVx1_ASAP7_75t_L g522 ( .A(n_102), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_103), .A2(n_124), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx2_ASAP7_75t_L g296 ( .A(n_105), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_106), .A2(n_282), .B1(n_440), .B2(n_443), .Y(n_552) );
XOR2x2_ASAP7_75t_L g705 ( .A(n_109), .B(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_111), .A2(n_128), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_112), .A2(n_126), .B1(n_447), .B2(n_635), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_113), .A2(n_227), .B1(n_362), .B2(n_364), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_116), .A2(n_165), .B1(n_647), .B2(n_648), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_117), .A2(n_253), .B1(n_436), .B2(n_437), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_118), .A2(n_230), .B1(n_503), .B2(n_538), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_120), .B(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_122), .A2(n_276), .B1(n_327), .B2(n_397), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_123), .A2(n_237), .B1(n_440), .B2(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_125), .B(n_600), .Y(n_675) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_130), .A2(n_205), .B1(n_314), .B2(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_131), .B(n_428), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_132), .A2(n_201), .B1(n_327), .B2(n_622), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_133), .B(n_428), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_134), .B(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_136), .A2(n_266), .B1(n_342), .B2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_139), .A2(n_152), .B1(n_505), .B2(n_506), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_141), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_142), .B(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_144), .A2(n_247), .B1(n_378), .B2(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_145), .A2(n_223), .B1(n_393), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_146), .A2(n_264), .B1(n_677), .B2(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g316 ( .A(n_147), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_148), .A2(n_180), .B1(n_607), .B2(n_609), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_149), .A2(n_262), .B1(n_400), .B2(n_604), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_150), .A2(n_176), .B1(n_595), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_156), .A2(n_278), .B1(n_371), .B2(n_640), .Y(n_672) );
XNOR2xp5_ASAP7_75t_L g721 ( .A(n_157), .B(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_158), .A2(n_191), .B1(n_358), .B2(n_359), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_160), .A2(n_243), .B1(n_437), .B2(n_491), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_162), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_163), .B(n_529), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_164), .Y(n_817) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_166), .A2(n_765), .B1(n_795), .B2(n_796), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_166), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_168), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_169), .A2(n_231), .B1(n_373), .B2(n_375), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_172), .A2(n_207), .B1(n_358), .B2(n_359), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_173), .A2(n_195), .B1(n_358), .B2(n_359), .Y(n_709) );
AO22x2_ASAP7_75t_L g487 ( .A1(n_175), .A2(n_488), .B1(n_514), .B2(n_515), .Y(n_487) );
INVx1_ASAP7_75t_L g515 ( .A(n_175), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_178), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_179), .A2(n_251), .B1(n_611), .B2(n_613), .Y(n_610) );
XNOR2x1_ASAP7_75t_L g452 ( .A(n_181), .B(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_184), .A2(n_209), .B1(n_375), .B2(n_378), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_185), .A2(n_272), .B1(n_663), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_187), .A2(n_222), .B1(n_512), .B2(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_188), .A2(n_221), .B1(n_436), .B2(n_474), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_189), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_190), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_192), .A2(n_265), .B1(n_436), .B2(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_193), .A2(n_212), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_197), .A2(n_240), .B1(n_399), .B2(n_400), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_198), .A2(n_256), .B1(n_397), .B2(n_498), .Y(n_713) );
INVx1_ASAP7_75t_L g556 ( .A(n_200), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_204), .B(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_206), .A2(n_244), .B1(n_512), .B2(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_208), .A2(n_255), .B1(n_430), .B2(n_476), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_210), .B(n_529), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_211), .A2(n_254), .B1(n_502), .B2(n_590), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_213), .B(n_308), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_216), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_224), .Y(n_793) );
AO22x2_ASAP7_75t_L g558 ( .A1(n_225), .A2(n_559), .B1(n_570), .B2(n_571), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_225), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_226), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g754 ( .A(n_226), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_228), .A2(n_257), .B1(n_471), .B2(n_472), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_229), .A2(n_268), .B1(n_327), .B2(n_332), .Y(n_326) );
INVx1_ASAP7_75t_L g293 ( .A(n_232), .Y(n_293) );
AND2x2_ASAP7_75t_R g798 ( .A(n_232), .B(n_754), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_233), .A2(n_236), .B1(n_666), .B2(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g627 ( .A(n_234), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_234), .A2(n_619), .B1(n_650), .B2(n_831), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_234), .A2(n_633), .B1(n_642), .B2(n_832), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_234), .B(n_628), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_235), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_238), .A2(n_383), .B1(n_384), .B2(n_420), .Y(n_382) );
INVx1_ASAP7_75t_L g420 ( .A(n_238), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_242), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_248), .B(n_295), .Y(n_294) );
XNOR2x1_ASAP7_75t_L g304 ( .A(n_249), .B(n_305), .Y(n_304) );
XOR2xp5_ASAP7_75t_L g449 ( .A(n_249), .B(n_305), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_258), .B(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_259), .A2(n_273), .B1(n_399), .B2(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_260), .A2(n_271), .B1(n_446), .B2(n_447), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_274), .A2(n_279), .B1(n_433), .B2(n_471), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_275), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_285), .Y(n_778) );
CKINVDCx6p67_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g829 ( .A(n_292), .B(n_294), .Y(n_829) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_293), .B(n_754), .Y(n_753) );
AOI21xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_577), .B(n_751), .Y(n_297) );
INVx1_ASAP7_75t_L g762 ( .A(n_298), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_484), .B1(n_485), .B2(n_576), .Y(n_298) );
INVx1_ASAP7_75t_L g576 ( .A(n_299), .Y(n_576) );
XNOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_451), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_381), .B2(n_450), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_304), .A2(n_423), .B1(n_424), .B2(n_449), .Y(n_422) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_356), .Y(n_305) );
NAND4xp25_ASAP7_75t_L g306 ( .A(n_307), .B(n_326), .C(n_337), .D(n_346), .Y(n_306) );
INVx4_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx3_ASAP7_75t_L g388 ( .A(n_309), .Y(n_388) );
INVx4_ASAP7_75t_SL g529 ( .A(n_309), .Y(n_529) );
INVx3_ASAP7_75t_SL g602 ( .A(n_309), .Y(n_602) );
BUFx2_ASAP7_75t_L g645 ( .A(n_309), .Y(n_645) );
INVx3_ASAP7_75t_L g695 ( .A(n_309), .Y(n_695) );
INVx6_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_319), .Y(n_310) );
AND2x4_ASAP7_75t_L g344 ( .A(n_311), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g353 ( .A(n_311), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g428 ( .A(n_311), .B(n_319), .Y(n_428) );
AND2x2_ASAP7_75t_L g434 ( .A(n_311), .B(n_345), .Y(n_434) );
AND2x2_ASAP7_75t_L g437 ( .A(n_311), .B(n_354), .Y(n_437) );
AND2x2_ASAP7_75t_L g471 ( .A(n_311), .B(n_345), .Y(n_471) );
AND2x2_ASAP7_75t_L g474 ( .A(n_311), .B(n_354), .Y(n_474) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_317), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_312), .B(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_312), .Y(n_336) );
INVx2_ASAP7_75t_L g341 ( .A(n_312), .Y(n_341) );
OAI22x1_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_315), .B2(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g318 ( .A(n_314), .Y(n_318) );
INVx2_ASAP7_75t_L g322 ( .A(n_314), .Y(n_322) );
INVx1_ASAP7_75t_L g325 ( .A(n_314), .Y(n_325) );
INVx2_ASAP7_75t_L g331 ( .A(n_317), .Y(n_331) );
AND2x2_ASAP7_75t_L g340 ( .A(n_317), .B(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g360 ( .A(n_317), .Y(n_360) );
AND2x4_ASAP7_75t_L g363 ( .A(n_319), .B(n_330), .Y(n_363) );
AND2x2_ASAP7_75t_L g370 ( .A(n_319), .B(n_340), .Y(n_370) );
AND2x4_ASAP7_75t_L g377 ( .A(n_319), .B(n_366), .Y(n_377) );
AND2x2_ASAP7_75t_L g441 ( .A(n_319), .B(n_366), .Y(n_441) );
AND2x2_ASAP7_75t_L g443 ( .A(n_319), .B(n_330), .Y(n_443) );
AND2x6_ASAP7_75t_L g446 ( .A(n_319), .B(n_340), .Y(n_446) );
AND2x2_ASAP7_75t_L g462 ( .A(n_319), .B(n_330), .Y(n_462) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g329 ( .A(n_321), .B(n_323), .Y(n_329) );
AND2x2_ASAP7_75t_L g335 ( .A(n_321), .B(n_324), .Y(n_335) );
INVx1_ASAP7_75t_L g350 ( .A(n_321), .Y(n_350) );
INVxp67_ASAP7_75t_L g345 ( .A(n_323), .Y(n_345) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g349 ( .A(n_324), .B(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_327), .Y(n_395) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g499 ( .A(n_328), .Y(n_499) );
BUFx3_ASAP7_75t_L g608 ( .A(n_328), .Y(n_608) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g339 ( .A(n_329), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g373 ( .A(n_329), .B(n_366), .Y(n_373) );
AND2x4_ASAP7_75t_L g430 ( .A(n_329), .B(n_330), .Y(n_430) );
AND2x2_ASAP7_75t_L g433 ( .A(n_329), .B(n_340), .Y(n_433) );
AND2x2_ASAP7_75t_L g444 ( .A(n_329), .B(n_366), .Y(n_444) );
AND2x2_ASAP7_75t_L g472 ( .A(n_329), .B(n_340), .Y(n_472) );
AND2x2_ASAP7_75t_L g348 ( .A(n_330), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g436 ( .A(n_330), .B(n_349), .Y(n_436) );
AND2x4_ASAP7_75t_L g366 ( .A(n_331), .B(n_341), .Y(n_366) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_332), .Y(n_609) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g397 ( .A(n_333), .Y(n_397) );
INVx2_ASAP7_75t_L g807 ( .A(n_333), .Y(n_807) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx12f_ASAP7_75t_L g622 ( .A(n_334), .Y(n_622) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
AND2x4_ASAP7_75t_L g359 ( .A(n_335), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g365 ( .A(n_335), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g414 ( .A(n_335), .B(n_360), .Y(n_414) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_335), .B(n_336), .Y(n_431) );
AND2x4_ASAP7_75t_L g440 ( .A(n_335), .B(n_366), .Y(n_440) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_335), .B(n_336), .Y(n_476) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_339), .Y(n_399) );
BUFx3_ASAP7_75t_L g496 ( .A(n_339), .Y(n_496) );
AND2x2_ASAP7_75t_L g358 ( .A(n_340), .B(n_349), .Y(n_358) );
AND2x2_ASAP7_75t_L g411 ( .A(n_340), .B(n_349), .Y(n_411) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_SL g400 ( .A(n_343), .Y(n_400) );
INVx1_ASAP7_75t_L g527 ( .A(n_343), .Y(n_527) );
INVx2_ASAP7_75t_L g605 ( .A(n_343), .Y(n_605) );
INVx2_ASAP7_75t_L g648 ( .A(n_343), .Y(n_648) );
INVx2_ASAP7_75t_L g692 ( .A(n_343), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_343), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_343), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_814) );
INVx6_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g811 ( .A(n_347), .Y(n_811) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
INVx3_ASAP7_75t_L g492 ( .A(n_348), .Y(n_492) );
AND2x4_ASAP7_75t_L g380 ( .A(n_349), .B(n_366), .Y(n_380) );
AND2x6_ASAP7_75t_L g447 ( .A(n_349), .B(n_366), .Y(n_447) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_350), .Y(n_355) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_SL g393 ( .A(n_353), .Y(n_393) );
INVx2_ASAP7_75t_L g494 ( .A(n_353), .Y(n_494) );
BUFx3_ASAP7_75t_L g626 ( .A(n_353), .Y(n_626) );
BUFx4f_ASAP7_75t_L g773 ( .A(n_353), .Y(n_773) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_361), .C(n_367), .D(n_374), .Y(n_356) );
BUFx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx6_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_SL g510 ( .A(n_365), .Y(n_510) );
BUFx2_ASAP7_75t_SL g590 ( .A(n_365), .Y(n_590) );
BUFx3_ASAP7_75t_L g668 ( .A(n_365), .Y(n_668) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
INVx2_ASAP7_75t_SL g512 ( .A(n_369), .Y(n_512) );
INVx2_ASAP7_75t_L g534 ( .A(n_369), .Y(n_534) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g635 ( .A(n_370), .Y(n_635) );
BUFx2_ASAP7_75t_L g663 ( .A(n_370), .Y(n_663) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g503 ( .A(n_372), .Y(n_503) );
INVx2_ASAP7_75t_L g641 ( .A(n_372), .Y(n_641) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_373), .Y(n_595) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx4_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
INVx2_ASAP7_75t_SL g538 ( .A(n_376), .Y(n_538) );
INVx3_ASAP7_75t_SL g640 ( .A(n_376), .Y(n_640) );
INVx2_ASAP7_75t_L g698 ( .A(n_376), .Y(n_698) );
INVx2_ASAP7_75t_SL g746 ( .A(n_376), .Y(n_746) );
INVx8_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g513 ( .A(n_379), .Y(n_513) );
INVx2_ASAP7_75t_L g597 ( .A(n_379), .Y(n_597) );
INVx2_ASAP7_75t_L g636 ( .A(n_379), .Y(n_636) );
INVx2_ASAP7_75t_SL g664 ( .A(n_379), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_379), .A2(n_781), .B1(n_782), .B2(n_783), .Y(n_780) );
INVx2_ASAP7_75t_L g821 ( .A(n_379), .Y(n_821) );
INVx8_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g450 ( .A(n_381), .Y(n_450) );
XNOR2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_421), .Y(n_381) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_401), .Y(n_384) );
NAND4xp25_ASAP7_75t_SL g385 ( .A(n_386), .B(n_389), .C(n_394), .D(n_398), .Y(n_385) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g813 ( .A(n_393), .Y(n_813) );
BUFx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx4f_ASAP7_75t_SL g604 ( .A(n_399), .Y(n_604) );
BUFx2_ASAP7_75t_L g647 ( .A(n_399), .Y(n_647) );
INVx1_ASAP7_75t_L g816 ( .A(n_399), .Y(n_816) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .C(n_407), .D(n_415), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g502 ( .A(n_404), .Y(n_502) );
INVx2_ASAP7_75t_L g589 ( .A(n_404), .Y(n_589) );
INVx3_ASAP7_75t_L g638 ( .A(n_404), .Y(n_638) );
INVx1_ASAP7_75t_SL g666 ( .A(n_404), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_404), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_406), .Y(n_509) );
INVx2_ASAP7_75t_L g593 ( .A(n_406), .Y(n_593) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g630 ( .A(n_410), .Y(n_630) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_411), .Y(n_505) );
BUFx3_ASAP7_75t_L g671 ( .A(n_411), .Y(n_671) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_413), .A2(n_786), .B1(n_787), .B2(n_789), .Y(n_785) );
INVx5_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g631 ( .A(n_414), .Y(n_631) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g749 ( .A(n_419), .Y(n_749) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_426), .B(n_438), .Y(n_425) );
NAND4xp25_ASAP7_75t_SL g426 ( .A(n_427), .B(n_429), .C(n_432), .D(n_435), .Y(n_426) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .C(n_445), .D(n_448), .Y(n_438) );
AO22x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_465), .B1(n_482), .B2(n_483), .Y(n_451) );
INVx1_ASAP7_75t_L g482 ( .A(n_452), .Y(n_482) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_459), .Y(n_453) );
NAND4xp25_ASAP7_75t_SL g454 ( .A(n_455), .B(n_456), .C(n_457), .D(n_458), .Y(n_454) );
NAND4xp25_ASAP7_75t_SL g459 ( .A(n_460), .B(n_461), .C(n_463), .D(n_464), .Y(n_459) );
INVx1_ASAP7_75t_L g483 ( .A(n_465), .Y(n_483) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .C(n_475), .Y(n_469) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .C(n_480), .D(n_481), .Y(n_477) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_516), .B1(n_573), .B2(n_574), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g573 ( .A(n_487), .Y(n_573) );
INVx1_ASAP7_75t_SL g514 ( .A(n_488), .Y(n_514) );
NOR4xp75_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .C(n_500), .D(n_507), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
INVx2_ASAP7_75t_SL g612 ( .A(n_491), .Y(n_612) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g531 ( .A(n_492), .Y(n_531) );
INVx1_ASAP7_75t_L g733 ( .A(n_492), .Y(n_733) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g614 ( .A(n_494), .Y(n_614) );
INVx1_ASAP7_75t_L g682 ( .A(n_496), .Y(n_682) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g677 ( .A(n_499), .Y(n_677) );
INVx1_ASAP7_75t_L g769 ( .A(n_499), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OA22x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_557), .B2(n_572), .Y(n_517) );
OA22x2_ASAP7_75t_L g575 ( .A1(n_518), .A2(n_519), .B1(n_557), .B2(n_572), .Y(n_575) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OA22x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_539), .B2(n_540), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
XNOR2x2_ASAP7_75t_SL g521 ( .A(n_522), .B(n_523), .Y(n_521) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_532), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .C(n_528), .D(n_530), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .C(n_536), .D(n_537), .Y(n_532) );
INVx3_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
XOR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_556), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVxp67_ASAP7_75t_L g572 ( .A(n_557), .Y(n_572) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g571 ( .A(n_559), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g559 ( .A(n_560), .B(n_565), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .D(n_564), .Y(n_560) );
NAND4xp25_ASAP7_75t_SL g565 ( .A(n_566), .B(n_567), .C(n_568), .D(n_569), .Y(n_565) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g761 ( .A(n_577), .Y(n_761) );
XOR2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_654), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_582), .B1(n_615), .B2(n_653), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_586), .B(n_598), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .C(n_591), .D(n_596), .Y(n_586) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g794 ( .A(n_595), .Y(n_794) );
NAND4xp25_ASAP7_75t_SL g598 ( .A(n_599), .B(n_603), .C(n_606), .D(n_610), .Y(n_598) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_601), .A2(n_725), .B1(n_726), .B2(n_727), .C(n_728), .Y(n_724) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g737 ( .A(n_604), .Y(n_737) );
BUFx6f_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g727 ( .A(n_608), .Y(n_727) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_614), .A2(n_730), .B1(n_731), .B2(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g653 ( .A(n_615), .Y(n_653) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND4xp75_ASAP7_75t_L g616 ( .A(n_617), .B(n_649), .C(n_651), .D(n_652), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_632), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_623), .C(n_628), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g679 ( .A(n_622), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g650 ( .A(n_624), .Y(n_650) );
BUFx6f_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx6f_ASAP7_75t_L g743 ( .A(n_630), .Y(n_743) );
INVx1_ASAP7_75t_L g788 ( .A(n_630), .Y(n_788) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_633), .B(n_642), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_637), .C(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
XNOR2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_718), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_684), .B2(n_685), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
XOR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_683), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_673), .Y(n_659) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_665), .C(n_669), .D(n_672), .Y(n_660) );
INVx1_ASAP7_75t_L g782 ( .A(n_662), .Y(n_782) );
BUFx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g779 ( .A(n_667), .Y(n_779) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .C(n_676), .D(n_680), .Y(n_673) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OA22x2_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_704), .B2(n_705), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g703 ( .A(n_688), .Y(n_703) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_696), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .C(n_693), .D(n_694), .Y(n_689) );
NAND4xp25_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .C(n_700), .D(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g792 ( .A(n_698), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_704), .A2(n_705), .B1(n_721), .B2(n_750), .Y(n_720) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_712), .C(n_715), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .C(n_710), .D(n_711), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g750 ( .A(n_721), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_739), .Y(n_722) );
NOR3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_729), .C(n_735), .Y(n_723) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_744), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_753), .B(n_756), .Y(n_828) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
OAI222xp33_ASAP7_75t_R g763 ( .A1(n_764), .A2(n_797), .B1(n_799), .B2(n_801), .C1(n_826), .C2(n_829), .Y(n_763) );
INVx1_ASAP7_75t_SL g796 ( .A(n_765), .Y(n_796) );
AND3x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_775), .C(n_784), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_771), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_768), .B(n_770), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_774), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_780), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_790), .Y(n_784) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_790) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_818), .Y(n_803) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_809), .C(n_814), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_808), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_823), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx1_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
CKINVDCx6p67_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
endmodule