module fake_jpeg_20018_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_28),
.B(n_17),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_36),
.C(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_26),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_19),
.B1(n_23),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_43),
.B1(n_38),
.B2(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_65),
.Y(n_92)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_24),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_25),
.B(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_94),
.B1(n_87),
.B2(n_75),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_43),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_26),
.B(n_47),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_23),
.B1(n_33),
.B2(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_88),
.B1(n_56),
.B2(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_94),
.Y(n_111)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_103),
.B1(n_109),
.B2(n_122),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_107),
.B(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_38),
.B1(n_47),
.B2(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_118),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_37),
.B(n_45),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_78),
.A2(n_38),
.B1(n_66),
.B2(n_55),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_88),
.B1(n_68),
.B2(n_93),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_36),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_24),
.C(n_27),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_32),
.A3(n_37),
.B1(n_60),
.B2(n_16),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_37),
.A3(n_31),
.B1(n_20),
.B2(n_16),
.Y(n_133)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_39),
.B1(n_35),
.B2(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_125),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_81),
.B(n_73),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_124),
.A2(n_130),
.B(n_133),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_37),
.CI(n_91),
.CON(n_125),
.SN(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_31),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_135),
.C(n_141),
.Y(n_161)
);

OAI21x1_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_90),
.B(n_84),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_68),
.B1(n_76),
.B2(n_74),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_115),
.B1(n_121),
.B2(n_119),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_145),
.Y(n_165)
);

NOR2x1p5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_35),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_144),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_27),
.B(n_24),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_143),
.B(n_146),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_52),
.C(n_60),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_102),
.B(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_35),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_83),
.B1(n_76),
.B2(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_39),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_148),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_29),
.A3(n_39),
.B1(n_34),
.B2(n_27),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_34),
.B(n_1),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_0),
.B(n_1),
.Y(n_159)
);

NOR2x1p5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_60),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_98),
.A3(n_121),
.B1(n_119),
.B2(n_96),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_155),
.A2(n_175),
.B1(n_178),
.B2(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_146),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_21),
.B1(n_95),
.B2(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_166),
.B(n_124),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_110),
.B1(n_96),
.B2(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_160),
.A2(n_171),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_167),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_129),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_137),
.B1(n_151),
.B2(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_122),
.B1(n_110),
.B2(n_104),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_180),
.B1(n_145),
.B2(n_148),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_118),
.B1(n_104),
.B2(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_120),
.B1(n_97),
.B2(n_95),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_123),
.C(n_135),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_211),
.C(n_180),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_195),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_138),
.B(n_129),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_140),
.B(n_131),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_194),
.B1(n_198),
.B2(n_203),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_125),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_199),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_183),
.B(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_201),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_29),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_15),
.B(n_14),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_159),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_12),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_155),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_11),
.C(n_3),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_173),
.B1(n_176),
.B2(n_172),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_220),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_191),
.B1(n_196),
.B2(n_212),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_219),
.A2(n_2),
.B(n_4),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_164),
.C(n_163),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_188),
.C(n_197),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_176),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_227),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_157),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_231),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_152),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_152),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_160),
.Y(n_236)
);

AOI211xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_170),
.B(n_167),
.C(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_11),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_194),
.B1(n_203),
.B2(n_198),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_247),
.B1(n_226),
.B2(n_232),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_246),
.C(n_251),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_188),
.C(n_190),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_196),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_260),
.B(n_216),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_211),
.B1(n_208),
.B2(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_213),
.C(n_204),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_219),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_204),
.B1(n_189),
.B2(n_206),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_6),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_205),
.C(n_3),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_215),
.C(n_220),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_223),
.B(n_217),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_227),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_7),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_225),
.C(n_230),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_276),
.C(n_246),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_272),
.Y(n_282)
);

MAJx2_ASAP7_75t_R g271 ( 
.A(n_260),
.B(n_228),
.C(n_231),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_236),
.B(n_226),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_274),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_4),
.B(n_5),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_277),
.B1(n_257),
.B2(n_253),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_6),
.C(n_7),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_265),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_264),
.A2(n_244),
.B1(n_255),
.B2(n_249),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_290),
.Y(n_301)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_243),
.B1(n_245),
.B2(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_288),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_241),
.C(n_243),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_256),
.B1(n_241),
.B2(n_9),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_292),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_304),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_269),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_299),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_273),
.B(n_262),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_272),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_263),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_288),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_276),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_279),
.B(n_267),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_268),
.C(n_274),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_301),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_312),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_310),
.B(n_314),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_282),
.B(n_280),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_284),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_302),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_292),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_298),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_318),
.Y(n_323)
);

AOI21x1_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_314),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_301),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_320),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_316),
.Y(n_326)
);

AOI321xp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_323),
.A3(n_322),
.B1(n_324),
.B2(n_318),
.C(n_321),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_313),
.B(n_9),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_8),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_10),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_10),
.Y(n_331)
);


endmodule