module fake_jpeg_23233_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_40),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_21),
.B2(n_23),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_15),
.B1(n_21),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_54),
.B1(n_16),
.B2(n_25),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_15),
.B1(n_18),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_30),
.B1(n_18),
.B2(n_27),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_32),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g101 ( 
.A(n_58),
.Y(n_101)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_72),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_53),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_77),
.B1(n_80),
.B2(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_18),
.B1(n_27),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_74),
.Y(n_103)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_69),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_75),
.Y(n_115)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_79),
.Y(n_95)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_42),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_47),
.B1(n_46),
.B2(n_24),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_16),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_89),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_88),
.B(n_94),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_53),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_0),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_93),
.B(n_99),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_1),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_113),
.B1(n_65),
.B2(n_76),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_79),
.B1(n_24),
.B2(n_25),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_67),
.A2(n_33),
.B(n_32),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_76),
.B1(n_112),
.B2(n_95),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_56),
.B(n_33),
.C(n_32),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_110),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_60),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_48),
.B1(n_25),
.B2(n_24),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_125),
.B(n_126),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_119),
.B1(n_127),
.B2(n_128),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_78),
.B1(n_62),
.B2(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_123),
.Y(n_152)
);

AO21x2_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_65),
.B(n_71),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_130),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_86),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_100),
.B(n_97),
.C(n_110),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_82),
.B1(n_76),
.B2(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_59),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_59),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_48),
.B1(n_64),
.B2(n_75),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_108),
.B1(n_114),
.B2(n_87),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_80),
.B1(n_44),
.B2(n_69),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_3),
.Y(n_176)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_79),
.B1(n_69),
.B2(n_80),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_87),
.B(n_105),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_144),
.A2(n_158),
.B(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_96),
.B(n_93),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_166),
.B(n_122),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_160),
.B1(n_165),
.B2(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_93),
.B1(n_108),
.B2(n_114),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_176),
.B1(n_120),
.B2(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_164),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_91),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_168),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_91),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_106),
.C(n_102),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_161),
.C(n_171),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_95),
.B1(n_94),
.B2(n_106),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_102),
.C(n_88),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_40),
.B(n_39),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_95),
.B1(n_39),
.B2(n_35),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_125),
.A2(n_39),
.B(n_35),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_35),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_33),
.B1(n_25),
.B2(n_16),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_1),
.C(n_2),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

NAND2xp67_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_3),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_178),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_181),
.B(n_182),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_129),
.B(n_134),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_141),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_187),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_119),
.B1(n_123),
.B2(n_142),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_171),
.B1(n_149),
.B2(n_151),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_128),
.B1(n_124),
.B2(n_131),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_191),
.B1(n_208),
.B2(n_175),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_135),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_150),
.B(n_161),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_159),
.B(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_193),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_174),
.B1(n_160),
.B2(n_163),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_136),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_175),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_152),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_198),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_155),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_204),
.B(n_207),
.Y(n_210)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_139),
.B1(n_137),
.B2(n_5),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_220),
.B1(n_228),
.B2(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_168),
.C(n_156),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_226),
.C(n_232),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_158),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_224),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_175),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_180),
.A2(n_3),
.B(n_4),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_181),
.B1(n_178),
.B2(n_184),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_10),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_191),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_6),
.C(n_8),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_229),
.B1(n_197),
.B2(n_216),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_252),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_182),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_225),
.B(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_192),
.C(n_195),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_224),
.C(n_222),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_195),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_242),
.Y(n_255)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_204),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_199),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_189),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_249),
.Y(n_257)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_208),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_215),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_210),
.B(n_185),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_188),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_179),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_243),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_264),
.C(n_235),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_228),
.B1(n_206),
.B2(n_201),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_242),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_210),
.C(n_232),
.Y(n_264)
);

FAx1_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_211),
.CI(n_220),
.CON(n_265),
.SN(n_265)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_262),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_217),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_245),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_273),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_247),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_238),
.C(n_235),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_283),
.C(n_245),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_270),
.B1(n_283),
.B2(n_273),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_257),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_231),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_6),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_274),
.B(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_263),
.C(n_260),
.Y(n_283)
);

FAx1_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_265),
.CI(n_240),
.CON(n_284),
.SN(n_284)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_289),
.B(n_10),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_294),
.C(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_9),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_255),
.C(n_8),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_297),
.B(n_303),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_287),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_9),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_10),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_308),
.C(n_291),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_14),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_285),
.B(n_284),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AO21x2_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_298),
.B(n_13),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_311),
.B(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_304),
.C(n_13),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_12),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_12),
.B(n_14),
.Y(n_318)
);


endmodule