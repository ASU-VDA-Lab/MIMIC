module fake_jpeg_1_n_467 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_48),
.Y(n_117)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_52),
.B(n_37),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_53),
.Y(n_143)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_23),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_95),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_86),
.B(n_14),
.Y(n_150)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_90),
.Y(n_142)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_91),
.B(n_92),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_93),
.Y(n_97)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_96),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_62),
.B1(n_70),
.B2(n_53),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_98),
.A2(n_120),
.B1(n_128),
.B2(n_132),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_47),
.B1(n_36),
.B2(n_34),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_110),
.A2(n_126),
.B1(n_29),
.B2(n_40),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_52),
.A2(n_36),
.B1(n_32),
.B2(n_34),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_19),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_79),
.A2(n_31),
.B1(n_33),
.B2(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_124),
.B(n_127),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_76),
.A2(n_33),
.B1(n_31),
.B2(n_37),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_44),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_82),
.A2(n_29),
.B1(n_42),
.B2(n_27),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_65),
.A2(n_77),
.B1(n_66),
.B2(n_92),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_54),
.A2(n_29),
.B1(n_27),
.B2(n_42),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_29),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_89),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_1),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_153),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_154),
.B(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_96),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_157),
.B(n_158),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_161),
.A2(n_146),
.B1(n_152),
.B2(n_108),
.Y(n_231)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_90),
.B(n_93),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_164),
.A2(n_140),
.B(n_133),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_119),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_63),
.C(n_29),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_135),
.C(n_114),
.Y(n_230)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_12),
.B(n_27),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_R g215 ( 
.A(n_169),
.B(n_110),
.Y(n_215)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_175),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_174),
.A2(n_200),
.B1(n_126),
.B2(n_119),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_177),
.Y(n_228)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_1),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_180),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_105),
.B(n_107),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_188),
.Y(n_214)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_134),
.B(n_2),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_192),
.Y(n_227)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_194),
.Y(n_220)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_197),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_2),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_202),
.Y(n_246)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_137),
.A2(n_40),
.B1(n_19),
.B2(n_5),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_141),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_98),
.Y(n_217)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_138),
.B1(n_97),
.B2(n_118),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_210),
.B1(n_164),
.B2(n_200),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_97),
.B1(n_118),
.B2(n_132),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_211),
.A2(n_153),
.B1(n_176),
.B2(n_159),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_225),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_240),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_231),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_144),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_249),
.A2(n_280),
.B1(n_215),
.B2(n_219),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_250),
.B(n_258),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_196),
.A3(n_167),
.B1(n_183),
.B2(n_160),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_182),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_192),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_266),
.Y(n_292)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_189),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_259),
.A2(n_282),
.B(n_242),
.Y(n_317)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_183),
.B1(n_174),
.B2(n_204),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_267),
.B1(n_273),
.B2(n_276),
.Y(n_305)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_187),
.B1(n_143),
.B2(n_194),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_213),
.B(n_184),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_269),
.Y(n_314)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_272),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_207),
.A2(n_191),
.B1(n_190),
.B2(n_185),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_277),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_165),
.B1(n_199),
.B2(n_202),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_210),
.A2(n_152),
.B1(n_168),
.B2(n_186),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_221),
.B1(n_219),
.B2(n_229),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_214),
.B(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_281),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_211),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_233),
.B(n_223),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_284),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_285),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_286),
.A2(n_309),
.B1(n_315),
.B2(n_4),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_253),
.A2(n_246),
.B(n_234),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_312),
.B(n_296),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_247),
.B(n_209),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_296),
.B(n_307),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_253),
.A2(n_222),
.B(n_232),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_206),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_297),
.B(n_282),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_206),
.C(n_226),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_285),
.C(n_283),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_265),
.A2(n_237),
.B1(n_226),
.B2(n_232),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_276),
.B(n_267),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_237),
.B1(n_222),
.B2(n_209),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_251),
.A2(n_229),
.B(n_234),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_275),
.A2(n_234),
.B(n_242),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_254),
.A2(n_242),
.B1(n_6),
.B2(n_7),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_317),
.A2(n_278),
.B1(n_266),
.B2(n_257),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_R g320 ( 
.A1(n_289),
.A2(n_263),
.B1(n_248),
.B2(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_322),
.B(n_348),
.Y(n_363)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_284),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_326),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_289),
.B(n_282),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_264),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_328),
.C(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_293),
.Y(n_331)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_281),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_336),
.C(n_342),
.Y(n_364)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_334),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_337),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_271),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_301),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_269),
.B1(n_6),
.B2(n_7),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_345),
.B1(n_346),
.B2(n_313),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_341),
.A2(n_343),
.B1(n_315),
.B2(n_287),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_310),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_286),
.B1(n_304),
.B2(n_290),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_312),
.B(n_299),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_4),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_9),
.Y(n_347)
);

XNOR2x2_ASAP7_75t_SL g351 ( 
.A(n_347),
.B(n_313),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_308),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_342),
.B(n_321),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_370),
.Y(n_381)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_354),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_319),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_360),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_287),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_307),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_367),
.C(n_328),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_369),
.B1(n_372),
.B2(n_341),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_336),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_330),
.B(n_294),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_368),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_343),
.A2(n_311),
.B1(n_305),
.B2(n_301),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_349),
.A2(n_317),
.B1(n_311),
.B2(n_318),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_318),
.B1(n_314),
.B2(n_295),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_325),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_370),
.A2(n_357),
.B1(n_325),
.B2(n_374),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_376),
.A2(n_384),
.B1(n_392),
.B2(n_395),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_366),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_385),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_364),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_321),
.C(n_344),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_367),
.C(n_368),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_374),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_389),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_371),
.A2(n_347),
.B(n_299),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_394),
.Y(n_401)
);

AOI21xp33_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_295),
.B(n_298),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_10),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_359),
.A2(n_340),
.B1(n_314),
.B2(n_298),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_375),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_306),
.B1(n_363),
.B2(n_10),
.Y(n_410)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_350),
.A2(n_334),
.B1(n_306),
.B2(n_300),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_355),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_360),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_352),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_404),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_364),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_394),
.A2(n_355),
.B1(n_361),
.B2(n_363),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_407),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_409),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_356),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_412),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_379),
.A2(n_10),
.B1(n_11),
.B2(n_387),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_413),
.A2(n_389),
.B1(n_393),
.B2(n_386),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_10),
.C(n_11),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_395),
.C(n_381),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_416),
.A2(n_418),
.B1(n_422),
.B2(n_423),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_400),
.A2(n_381),
.B1(n_386),
.B2(n_376),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g420 ( 
.A(n_415),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_420),
.B(n_409),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_393),
.Y(n_423)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_424),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_411),
.A2(n_381),
.B(n_392),
.Y(n_425)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_402),
.A2(n_11),
.B(n_401),
.Y(n_426)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_399),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_407),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_425),
.A2(n_402),
.B1(n_410),
.B2(n_398),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_436),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_429),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_408),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_434),
.B(n_439),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_414),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_440),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_421),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_419),
.B(n_427),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_441),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_446),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_426),
.Y(n_443)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_443),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_417),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_444),
.B(n_449),
.Y(n_453)
);

NAND2xp67_ASAP7_75t_SL g445 ( 
.A(n_431),
.B(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_445),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_435),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_448),
.A2(n_434),
.B(n_438),
.Y(n_451)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_451),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_447),
.A2(n_432),
.B(n_446),
.Y(n_452)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_452),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_456),
.B(n_451),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_454),
.Y(n_461)
);

OR2x6_ASAP7_75t_SL g460 ( 
.A(n_453),
.B(n_450),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_460),
.B(n_458),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_461),
.B(n_462),
.C(n_458),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_463),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_464),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_465),
.B(n_459),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_455),
.B(n_443),
.Y(n_467)
);


endmodule