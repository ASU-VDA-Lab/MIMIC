module fake_aes_11552_n_30 (n_3, n_1, n_2, n_0, n_30);
input n_3;
input n_1;
input n_2;
input n_0;
output n_30;
wire n_20;
wire n_5;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_4;
wire n_29;
wire n_7;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_2), .Y(n_4) );
NOR2xp33_ASAP7_75t_R g5 ( .A(n_3), .B(n_2), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_1), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_0), .Y(n_7) );
BUFx12f_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
NOR2xp33_ASAP7_75t_L g9 ( .A(n_6), .B(n_0), .Y(n_9) );
NOR3xp33_ASAP7_75t_SL g10 ( .A(n_6), .B(n_0), .C(n_1), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_7), .B(n_0), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx2_ASAP7_75t_SL g13 ( .A(n_8), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
NOR2xp67_ASAP7_75t_SL g15 ( .A(n_8), .B(n_7), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_9), .B(n_1), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_16), .B(n_11), .Y(n_18) );
INVxp67_ASAP7_75t_SL g19 ( .A(n_13), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_19), .B(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_15), .B1(n_5), .B2(n_10), .C(n_12), .Y(n_23) );
AOI322xp5_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_2), .A3(n_3), .B1(n_5), .B2(n_15), .C1(n_12), .C2(n_14), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_21), .B(n_3), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_25), .B(n_20), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_24), .B(n_12), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
INVx2_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_12), .B1(n_17), .B2(n_28), .Y(n_30) );
endmodule