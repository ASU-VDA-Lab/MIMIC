module real_jpeg_16329_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_0),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_71),
.B1(n_76),
.B2(n_80),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_2),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_3),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_4),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_35),
.B(n_215),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_243),
.A3(n_246),
.B1(n_250),
.B2(n_255),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_5),
.A2(n_243),
.A3(n_246),
.B1(n_250),
.B2(n_255),
.Y(n_281)
);

OAI32xp33_ASAP7_75t_L g283 ( 
.A1(n_5),
.A2(n_243),
.A3(n_246),
.B1(n_250),
.B2(n_255),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_5),
.A2(n_148),
.B1(n_296),
.B2(n_299),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_5),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_5),
.A2(n_50),
.B1(n_270),
.B2(n_388),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_177),
.B1(n_180),
.B2(n_186),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_6),
.A2(n_186),
.B1(n_259),
.B2(n_264),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_7),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_7),
.Y(n_185)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_7),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_7),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_8),
.A2(n_203),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_8),
.A2(n_138),
.B1(n_203),
.B2(n_319),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_84),
.B1(n_90),
.B2(n_95),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_95),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_9),
.A2(n_95),
.B1(n_311),
.B2(n_315),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_9),
.A2(n_95),
.B1(n_382),
.B2(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_11),
.A2(n_138),
.B1(n_143),
.B2(n_144),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_11),
.A2(n_143),
.B1(n_190),
.B2(n_194),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_13),
.Y(n_142)
);

BUFx4f_ASAP7_75t_L g263 ( 
.A(n_13),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_14),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_14),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_14),
.A2(n_126),
.B1(n_286),
.B2(n_289),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_14),
.A2(n_126),
.B1(n_370),
.B2(n_374),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_15),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_15),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_273),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_271),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_226),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_19),
.B(n_226),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_155),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_39),
.B2(n_44),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_38),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g208 ( 
.A1(n_39),
.A2(n_150),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_40),
.Y(n_213)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_42),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B1(n_66),
.B2(n_70),
.Y(n_49)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_50),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_50),
.A2(n_318),
.B1(n_322),
.B2(n_328),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_50),
.A2(n_369),
.B1(n_388),
.B2(n_392),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_51),
.Y(n_270)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_53),
.Y(n_146)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_55),
.Y(n_321)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_55),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_57),
.A2(n_136),
.B1(n_137),
.B2(n_146),
.Y(n_135)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_65),
.Y(n_373)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_76),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_134),
.C(n_147),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_82),
.B(n_229),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_96),
.B1(n_123),
.B2(n_133),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_83),
.A2(n_96),
.B1(n_133),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_89),
.Y(n_304)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_96),
.A2(n_123),
.B1(n_133),
.B2(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_105),
.B(n_111),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_117),
.B2(n_120),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_116),
.Y(n_236)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_119),
.Y(n_249)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_131),
.Y(n_298)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_133),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_134),
.A2(n_135),
.B1(n_147),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_136),
.A2(n_137),
.B1(n_258),
.B2(n_268),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_136),
.A2(n_268),
.B1(n_368),
.B2(n_376),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_141),
.Y(n_267)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_147),
.Y(n_230)
);

NOR2x1_ASAP7_75t_R g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_148),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_148),
.B(n_190),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_SL g359 ( 
.A1(n_148),
.A2(n_348),
.B(n_360),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_148),
.B(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_148),
.B(n_187),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_208),
.B1(n_214),
.B2(n_221),
.Y(n_207)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_207),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_199),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_176),
.B1(n_187),
.B2(n_188),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_158),
.A2(n_176),
.B1(n_187),
.B2(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_159),
.A2(n_233),
.B1(n_285),
.B2(n_292),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_159),
.A2(n_285),
.B1(n_292),
.B2(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_159),
.A2(n_292),
.B1(n_310),
.B2(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_167),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_170),
.Y(n_347)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_185),
.Y(n_362)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_187),
.Y(n_292)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.C(n_240),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_227),
.A2(n_228),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_231),
.A2(n_240),
.B1(n_241),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_256),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_249),
.Y(n_341)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_257),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_263),
.Y(n_375)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_267),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_305),
.B(n_400),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_275),
.B(n_279),
.Y(n_400)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.C(n_293),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_284),
.A2(n_293),
.B1(n_294),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

AOI21x1_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_335),
.B(n_399),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_332),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_332),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.C(n_329),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_308),
.A2(n_309),
.B1(n_329),
.B2(n_330),
.Y(n_364)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_364),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_318),
.Y(n_376)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_SL g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_325),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_365),
.B(n_398),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_363),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_363),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_357),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_338),
.A2(n_357),
.B1(n_358),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_342),
.A3(n_346),
.B1(n_348),
.B2(n_349),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_379),
.B(n_397),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_377),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_377),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_390),
.B(n_396),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_387),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_395),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_395),
.Y(n_396)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);


endmodule