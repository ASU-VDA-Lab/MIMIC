module fake_netlist_1_12180_n_21 (n_3, n_1, n_2, n_0, n_21);
input n_3;
input n_1;
input n_2;
input n_0;
output n_21;
wire n_20;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_4;
wire n_7;
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
OR2x6_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_SL g6 ( .A(n_2), .B(n_0), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_7), .B(n_0), .Y(n_8) );
AOI211x1_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_0), .B(n_1), .C(n_2), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_4), .B(n_1), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_8), .B(n_5), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_5), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_11), .B(n_5), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_11), .B(n_6), .Y(n_14) );
OAI21xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_12), .B(n_9), .Y(n_15) );
NOR2x1p5_ASAP7_75t_SL g16 ( .A(n_13), .B(n_2), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_15), .B(n_13), .Y(n_17) );
CKINVDCx16_ASAP7_75t_R g18 ( .A(n_16), .Y(n_18) );
NAND3xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_3), .C(n_2), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
AOI22xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_3), .B1(n_17), .B2(n_20), .Y(n_21) );
endmodule