module real_jpeg_23074_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_0),
.A2(n_28),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_0),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_0),
.A2(n_30),
.B1(n_32),
.B2(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_0),
.A2(n_57),
.B1(n_58),
.B2(n_130),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_0),
.A2(n_73),
.B1(n_74),
.B2(n_130),
.Y(n_251)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_4),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_7),
.A2(n_28),
.B1(n_52),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_7),
.A2(n_52),
.B1(n_73),
.B2(n_74),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_9),
.A2(n_35),
.B1(n_73),
.B2(n_74),
.Y(n_120)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_40),
.B1(n_73),
.B2(n_74),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_30),
.B1(n_32),
.B2(n_40),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_26),
.B(n_27),
.C(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_29),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_32),
.B(n_55),
.C(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_72),
.C(n_73),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_11),
.B(n_53),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_11),
.B(n_257),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_11),
.B(n_70),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_323),
.Y(n_16)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_41),
.B1(n_45),
.B2(n_320),
.C(n_322),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_18),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_18),
.B(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_18),
.B(n_41),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_19),
.A2(n_29),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_20),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_24),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_25),
.A2(n_32),
.B(n_40),
.Y(n_199)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_29),
.B(n_129),
.Y(n_169)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_30),
.A2(n_32),
.B1(n_55),
.B2(n_60),
.Y(n_63)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_34),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_38),
.B(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_40),
.A2(n_57),
.B(n_60),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_41),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_41),
.A2(n_96),
.B1(n_105),
.B2(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_42),
.A2(n_84),
.B(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_309),
.B(n_319),
.Y(n_45)
);

OAI211xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_133),
.B(n_148),
.C(n_308),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_106),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_48),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_48),
.B(n_106),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_48),
.B(n_135),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_81),
.CI(n_95),
.CON(n_48),
.SN(n_48)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_49),
.A2(n_50),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_65),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_61),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_53),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_54),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_54),
.B(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_54),
.A2(n_62),
.B(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_54)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_79)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_58),
.B(n_239),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_61),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_62),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_76),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_66),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_69),
.B(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_68),
.B(n_78),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_77),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_70),
.B(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_73),
.B(n_263),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_77),
.B(n_236),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_78),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_93),
.B1(n_137),
.B2(n_146),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_87),
.C(n_90),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_82),
.B(n_137),
.C(n_147),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_83),
.B(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_84),
.B(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_192),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_91),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_90),
.B(n_181),
.C(n_183),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_90),
.A2(n_91),
.B1(n_183),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_91),
.B(n_140),
.C(n_143),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_101),
.B(n_105),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_96),
.A2(n_102),
.B1(n_110),
.B2(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_96),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_96),
.A2(n_110),
.B1(n_221),
.B2(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_97),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_97),
.B(n_100),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_97),
.B(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_120),
.Y(n_164)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_104),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_104),
.B(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_111),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_126),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_114),
.B(n_121),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_115),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_117),
.A2(n_119),
.B(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_119),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_124),
.B(n_185),
.Y(n_276)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_149),
.C(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_147),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_144),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_173),
.B(n_307),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_170),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_152),
.B(n_170),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_153),
.B(n_156),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_158),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.C(n_168),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_159),
.A2(n_160),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_165),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_164),
.B(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_167),
.A2(n_168),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_167),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_167),
.A2(n_296),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_167),
.B(n_311),
.C(n_316),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_168),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_302),
.B(n_306),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_214),
.B(n_288),
.C(n_301),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_202),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_176),
.B(n_202),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_189),
.B2(n_201),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_179),
.B(n_188),
.C(n_201),
.Y(n_289)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_182),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_197),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_191),
.B(n_196),
.C(n_197),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_194),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_204),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_212),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_287),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_230),
.B(n_286),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_217),
.B(n_227),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_223),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_218),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_220),
.B(n_223),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_221),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_281),
.B(n_285),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_272),
.B(n_280),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_253),
.B(n_271),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_234),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_252),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_246),
.C(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_260),
.B(n_270),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_258),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_266),
.B(n_269),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_298),
.B2(n_299),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_299),
.C(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_318),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_318),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_317),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_313),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);


endmodule