module fake_aes_5488_n_31 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx6_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_12), .B(n_10), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_17), .B(n_0), .Y(n_19) );
AOI21x1_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_16), .B(n_15), .Y(n_20) );
A2O1A1Ixp33_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_13), .B(n_14), .C(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_13), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_14), .Y(n_23) );
AND2x4_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
AOI221x1_ASAP7_75t_SL g26 ( .A1(n_25), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_4), .Y(n_26) );
NOR3x1_ASAP7_75t_L g27 ( .A(n_25), .B(n_1), .C(n_3), .Y(n_27) );
AND4x1_ASAP7_75t_L g28 ( .A(n_27), .B(n_4), .C(n_5), .D(n_15), .Y(n_28) );
XNOR2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
AO221x1_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_14), .B1(n_8), .B2(n_11), .C(n_6), .Y(n_30) );
OA22x2_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_29), .B1(n_24), .B2(n_14), .Y(n_31) );
endmodule