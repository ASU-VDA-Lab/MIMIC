module real_aes_6927_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g175 ( .A1(n_0), .A2(n_176), .B(n_179), .C(n_183), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_1), .B(n_167), .Y(n_186) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_2), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g450 ( .A(n_2), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_3), .B(n_177), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_4), .A2(n_140), .B(n_143), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_5), .A2(n_135), .B(n_547), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_6), .A2(n_135), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_7), .B(n_167), .Y(n_553) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_8), .A2(n_169), .B(n_241), .Y(n_240) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_9), .A2(n_457), .B1(n_744), .B2(n_745), .C1(n_748), .C2(n_751), .Y(n_456) );
AND2x6_ASAP7_75t_L g140 ( .A(n_10), .B(n_141), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_11), .A2(n_140), .B(n_143), .C(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g513 ( .A(n_12), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_13), .B(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_13), .B(n_40), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_14), .B(n_182), .Y(n_524) );
INVx1_ASAP7_75t_L g161 ( .A(n_15), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_16), .B(n_177), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_17), .B(n_453), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_18), .A2(n_178), .B(n_533), .C(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_19), .B(n_167), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_20), .B(n_155), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_21), .A2(n_143), .B(n_146), .C(n_154), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_22), .A2(n_181), .B(n_249), .C(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_23), .B(n_182), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_24), .B(n_182), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_25), .Y(n_494) );
INVx1_ASAP7_75t_L g474 ( .A(n_26), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_27), .A2(n_143), .B(n_154), .C(n_244), .Y(n_243) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_29), .Y(n_520) );
INVx1_ASAP7_75t_L g488 ( .A(n_30), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_31), .A2(n_135), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_33), .A2(n_193), .B(n_194), .C(n_198), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_34), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_35), .A2(n_181), .B(n_550), .C(n_552), .Y(n_549) );
INVxp67_ASAP7_75t_L g489 ( .A(n_36), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_37), .B(n_246), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_38), .A2(n_143), .B(n_154), .C(n_473), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g548 ( .A(n_39), .Y(n_548) );
INVx1_ASAP7_75t_L g105 ( .A(n_40), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_41), .A2(n_183), .B(n_511), .C(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_42), .B(n_134), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_43), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_44), .B(n_177), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_45), .B(n_135), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_46), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_48), .A2(n_193), .B(n_198), .C(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g180 ( .A(n_49), .Y(n_180) );
INVx1_ASAP7_75t_L g224 ( .A(n_50), .Y(n_224) );
INVx1_ASAP7_75t_L g561 ( .A(n_51), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_52), .B(n_135), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_53), .Y(n_163) );
CKINVDCx14_ASAP7_75t_R g509 ( .A(n_54), .Y(n_509) );
INVx1_ASAP7_75t_L g141 ( .A(n_55), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_56), .B(n_135), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_57), .B(n_167), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_58), .A2(n_153), .B(n_209), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g160 ( .A(n_59), .Y(n_160) );
INVx1_ASAP7_75t_SL g551 ( .A(n_60), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_61), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_62), .B(n_177), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_63), .B(n_167), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_64), .B(n_178), .Y(n_259) );
INVx1_ASAP7_75t_L g497 ( .A(n_65), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_66), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_67), .B(n_148), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_68), .A2(n_143), .B(n_198), .C(n_207), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_69), .Y(n_233) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_71), .A2(n_135), .B(n_508), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_72), .A2(n_92), .B1(n_120), .B2(n_121), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_72), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_73), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_74), .A2(n_135), .B(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_75), .A2(n_100), .B1(n_746), .B2(n_747), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_75), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_76), .A2(n_134), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_77), .Y(n_471) );
INVx1_ASAP7_75t_L g531 ( .A(n_78), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_79), .B(n_151), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_80), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_81), .A2(n_135), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g534 ( .A(n_82), .Y(n_534) );
INVx2_ASAP7_75t_L g158 ( .A(n_83), .Y(n_158) );
INVx1_ASAP7_75t_L g523 ( .A(n_84), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_85), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_86), .B(n_182), .Y(n_260) );
INVx2_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
OR2x2_ASAP7_75t_L g447 ( .A(n_87), .B(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g460 ( .A(n_87), .B(n_449), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_88), .A2(n_143), .B(n_198), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_89), .B(n_135), .Y(n_191) );
INVx1_ASAP7_75t_L g195 ( .A(n_90), .Y(n_195) );
INVxp67_ASAP7_75t_L g236 ( .A(n_91), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_92), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_93), .B(n_169), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_94), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g208 ( .A(n_95), .Y(n_208) );
INVx1_ASAP7_75t_L g255 ( .A(n_96), .Y(n_255) );
INVx2_ASAP7_75t_L g564 ( .A(n_97), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_98), .A2(n_102), .B1(n_111), .B2(n_755), .Y(n_101) );
AND2x2_ASAP7_75t_L g226 ( .A(n_99), .B(n_157), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_100), .Y(n_746) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g756 ( .A(n_103), .Y(n_756) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
OR2x2_ASAP7_75t_L g463 ( .A(n_107), .B(n_449), .Y(n_463) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_107), .B(n_448), .Y(n_750) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_455), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g754 ( .A(n_113), .Y(n_754) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_445), .B(n_452), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_119), .B1(n_122), .B2(n_123), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_122), .A2(n_458), .B1(n_461), .B2(n_464), .Y(n_457) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_123), .A2(n_458), .B1(n_752), .B2(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_400), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_335), .Y(n_124) );
NAND4xp25_ASAP7_75t_SL g125 ( .A(n_126), .B(n_280), .C(n_304), .D(n_327), .Y(n_125) );
AOI221xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_217), .B1(n_251), .B2(n_264), .C(n_267), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_187), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_129), .A2(n_165), .B1(n_218), .B2(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_129), .B(n_188), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_129), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_129), .B(n_341), .Y(n_427) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
AND2x2_ASAP7_75t_L g295 ( .A(n_130), .B(n_188), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_130), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g318 ( .A(n_130), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g323 ( .A(n_130), .B(n_166), .Y(n_323) );
INVx2_ASAP7_75t_L g355 ( .A(n_130), .Y(n_355) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_130), .Y(n_399) );
AND2x2_ASAP7_75t_L g416 ( .A(n_130), .B(n_293), .Y(n_416) );
INVx5_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g334 ( .A(n_131), .B(n_293), .Y(n_334) );
AND2x4_ASAP7_75t_L g348 ( .A(n_131), .B(n_165), .Y(n_348) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_131), .Y(n_352) );
AND2x2_ASAP7_75t_L g372 ( .A(n_131), .B(n_287), .Y(n_372) );
AND2x2_ASAP7_75t_L g422 ( .A(n_131), .B(n_189), .Y(n_422) );
AND2x2_ASAP7_75t_L g432 ( .A(n_131), .B(n_166), .Y(n_432) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_162), .Y(n_131) );
AOI21xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_142), .B(n_155), .Y(n_132) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_136), .B(n_140), .Y(n_256) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g250 ( .A(n_138), .Y(n_250) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx3_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
INVx1_ASAP7_75t_L g246 ( .A(n_139), .Y(n_246) );
BUFx3_ASAP7_75t_L g154 ( .A(n_140), .Y(n_154) );
INVx4_ASAP7_75t_SL g185 ( .A(n_140), .Y(n_185) );
INVx5_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_144), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B(n_152), .Y(n_146) );
INVx2_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_151), .A2(n_195), .B(n_196), .C(n_197), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_151), .A2(n_197), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_151), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp5_ASAP7_75t_L g522 ( .A1(n_151), .A2(n_499), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_152), .A2(n_177), .B(n_474), .C(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_153), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_156), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g164 ( .A(n_157), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_157), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_157), .A2(n_221), .B(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_157), .A2(n_256), .B(n_471), .C(n_472), .Y(n_470) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_157), .A2(n_507), .B(n_514), .Y(n_506) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g170 ( .A(n_158), .B(n_159), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_164), .A2(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g288 ( .A(n_165), .B(n_188), .Y(n_288) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_165), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_165), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g378 ( .A(n_165), .Y(n_378) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g266 ( .A(n_166), .B(n_203), .Y(n_266) );
AND2x2_ASAP7_75t_L g293 ( .A(n_166), .B(n_204), .Y(n_293) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_171), .B(n_186), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_168), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_168), .A2(n_205), .B(n_215), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_168), .B(n_216), .Y(n_215) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_168), .A2(n_254), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_168), .B(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_168), .A2(n_493), .B(n_500), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_168), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_169), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_169), .A2(n_242), .B(n_243), .Y(n_241) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g263 ( .A(n_170), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_185), .Y(n_172) );
INVx2_ASAP7_75t_L g193 ( .A(n_174), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_174), .A2(n_185), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_174), .A2(n_185), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_174), .A2(n_185), .B(n_509), .C(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_174), .A2(n_185), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_174), .A2(n_185), .B(n_548), .C(n_549), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_SL g560 ( .A1(n_174), .A2(n_185), .B(n_561), .C(n_562), .Y(n_560) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_177), .B(n_236), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_177), .A2(n_210), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_178), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_181), .B(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g511 ( .A(n_182), .Y(n_511) );
INVx2_ASAP7_75t_L g499 ( .A(n_183), .Y(n_499) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_184), .Y(n_197) );
INVx1_ASAP7_75t_L g535 ( .A(n_184), .Y(n_535) );
INVx1_ASAP7_75t_L g198 ( .A(n_185), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_187), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_201), .Y(n_187) );
OR2x2_ASAP7_75t_L g319 ( .A(n_188), .B(n_202), .Y(n_319) );
AND2x2_ASAP7_75t_L g356 ( .A(n_188), .B(n_266), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_188), .B(n_287), .Y(n_367) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_188), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_188), .B(n_323), .Y(n_440) );
INVx5_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g265 ( .A(n_189), .Y(n_265) );
AND2x2_ASAP7_75t_L g274 ( .A(n_189), .B(n_202), .Y(n_274) );
AND2x2_ASAP7_75t_L g390 ( .A(n_189), .B(n_285), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_189), .B(n_323), .Y(n_412) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_199), .Y(n_189) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_202), .Y(n_358) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_203), .Y(n_310) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g287 ( .A(n_204), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_214), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_211), .C(n_212), .Y(n_207) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_210), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_210), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g552 ( .A(n_213), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_227), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_218), .B(n_300), .Y(n_419) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_219), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g271 ( .A(n_219), .B(n_272), .Y(n_271) );
INVx5_ASAP7_75t_SL g279 ( .A(n_219), .Y(n_279) );
OR2x2_ASAP7_75t_L g302 ( .A(n_219), .B(n_272), .Y(n_302) );
OR2x2_ASAP7_75t_L g312 ( .A(n_219), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g375 ( .A(n_219), .B(n_229), .Y(n_375) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_219), .B(n_228), .Y(n_413) );
NOR4xp25_ASAP7_75t_L g434 ( .A(n_219), .B(n_355), .C(n_435), .D(n_436), .Y(n_434) );
AND2x2_ASAP7_75t_L g444 ( .A(n_219), .B(n_276), .Y(n_444) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g269 ( .A(n_228), .B(n_265), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_228), .B(n_271), .Y(n_438) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_238), .Y(n_228) );
OR2x2_ASAP7_75t_L g278 ( .A(n_229), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g285 ( .A(n_229), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_229), .B(n_253), .Y(n_297) );
INVxp67_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_229), .B(n_272), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_229), .B(n_239), .Y(n_366) );
AND2x2_ASAP7_75t_L g381 ( .A(n_229), .B(n_276), .Y(n_381) );
OR2x2_ASAP7_75t_L g410 ( .A(n_229), .B(n_239), .Y(n_410) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_237), .Y(n_229) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_230), .A2(n_529), .B(n_536), .Y(n_528) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_230), .A2(n_546), .B(n_553), .Y(n_545) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_230), .A2(n_559), .B(n_565), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_238), .B(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_238), .B(n_279), .Y(n_418) );
OR2x2_ASAP7_75t_L g439 ( .A(n_238), .B(n_316), .Y(n_439) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g252 ( .A(n_239), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g276 ( .A(n_239), .B(n_272), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_239), .B(n_253), .Y(n_291) );
AND2x2_ASAP7_75t_L g361 ( .A(n_239), .B(n_285), .Y(n_361) );
AND2x2_ASAP7_75t_L g395 ( .A(n_239), .B(n_279), .Y(n_395) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_240), .B(n_279), .Y(n_298) );
AND2x2_ASAP7_75t_L g326 ( .A(n_240), .B(n_253), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B(n_248), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_248), .A2(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_251), .B(n_334), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_252), .A2(n_341), .B1(n_377), .B2(n_394), .C(n_396), .Y(n_393) );
INVx5_ASAP7_75t_SL g272 ( .A(n_253), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_257), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_256), .A2(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_256), .A2(n_520), .B(n_521), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g482 ( .A(n_263), .Y(n_482) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OAI33xp33_ASAP7_75t_L g292 ( .A1(n_265), .A2(n_293), .A3(n_294), .B1(n_296), .B2(n_299), .B3(n_303), .Y(n_292) );
OR2x2_ASAP7_75t_L g308 ( .A(n_265), .B(n_309), .Y(n_308) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_265), .A2(n_334), .A3(n_341), .B1(n_418), .B2(n_419), .C1(n_420), .C2(n_423), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_265), .B(n_293), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_SL g441 ( .A1(n_265), .A2(n_293), .B(n_442), .C(n_444), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_266), .A2(n_281), .B1(n_286), .B2(n_289), .C(n_292), .Y(n_280) );
INVx1_ASAP7_75t_L g373 ( .A(n_266), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_266), .B(n_422), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_270), .B1(n_273), .B2(n_275), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g350 ( .A(n_271), .B(n_285), .Y(n_350) );
AND2x2_ASAP7_75t_L g408 ( .A(n_271), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g316 ( .A(n_272), .B(n_279), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_272), .B(n_285), .Y(n_344) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_274), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_274), .B(n_352), .Y(n_406) );
OAI321xp33_ASAP7_75t_L g425 ( .A1(n_274), .A2(n_347), .A3(n_426), .B1(n_427), .B2(n_428), .C(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g392 ( .A(n_275), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_276), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g331 ( .A(n_276), .B(n_279), .Y(n_331) );
AOI321xp33_ASAP7_75t_L g389 ( .A1(n_276), .A2(n_293), .A3(n_390), .B1(n_391), .B2(n_392), .C(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g306 ( .A(n_278), .B(n_291), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_279), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_279), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_279), .B(n_365), .Y(n_402) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g325 ( .A(n_283), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g290 ( .A(n_284), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g398 ( .A(n_285), .Y(n_398) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_288), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g321 ( .A(n_293), .Y(n_321) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_295), .B(n_330), .Y(n_379) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OR2x2_ASAP7_75t_L g343 ( .A(n_298), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g388 ( .A(n_298), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_299), .A2(n_346), .B1(n_349), .B2(n_351), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g443 ( .A(n_302), .B(n_366), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B1(n_311), .B2(n_317), .C(n_320), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx2_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx1_ASAP7_75t_SL g387 ( .A(n_313), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_315), .B(n_365), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_315), .A2(n_383), .B(n_385), .Y(n_382) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g428 ( .A(n_316), .B(n_410), .Y(n_428) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g330 ( .A(n_319), .Y(n_330) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g374 ( .A(n_326), .B(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g436 ( .A(n_326), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B(n_332), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_330), .B(n_348), .Y(n_384) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g405 ( .A(n_334), .Y(n_405) );
NAND5xp2_ASAP7_75t_L g335 ( .A(n_336), .B(n_353), .C(n_362), .D(n_382), .E(n_389), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B(n_342), .C(n_345), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_349), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
OAI21xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_357), .B(n_359), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_354), .A2(n_408), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_407) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AOI321xp33_ASAP7_75t_L g362 ( .A1(n_355), .A2(n_363), .A3(n_367), .B1(n_368), .B2(n_374), .C(n_376), .Y(n_362) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g433 ( .A(n_367), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g385 ( .A(n_370), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NOR2xp67_ASAP7_75t_SL g397 ( .A(n_371), .B(n_378), .Y(n_397) );
AOI321xp33_ASAP7_75t_SL g429 ( .A1(n_374), .A2(n_430), .A3(n_431), .B1(n_432), .B2(n_433), .C(n_434), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_379), .C(n_380), .Y(n_376) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_387), .B(n_395), .Y(n_424) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .C(n_399), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_425), .C(n_437), .Y(n_400) );
OAI211xp5_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_403), .B(n_407), .C(n_417), .Y(n_401) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_405), .B(n_406), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_406), .A2(n_438), .B1(n_439), .B2(n_440), .C(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g426 ( .A(n_408), .Y(n_426) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g430 ( .A(n_428), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g455 ( .A1(n_452), .A2(n_456), .B(n_754), .Y(n_455) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g753 ( .A(n_462), .Y(n_753) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g752 ( .A(n_464), .Y(n_752) );
OR4x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_634), .C(n_681), .D(n_721), .Y(n_464) );
NAND3xp33_ASAP7_75t_SL g465 ( .A(n_466), .B(n_580), .C(n_609), .Y(n_465) );
AOI211xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_502), .B(n_537), .C(n_573), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_467), .A2(n_593), .B(n_610), .C(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_469), .B(n_572), .Y(n_571) );
INVx3_ASAP7_75t_SL g576 ( .A(n_469), .Y(n_576) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_469), .Y(n_588) );
AND2x4_ASAP7_75t_L g592 ( .A(n_469), .B(n_544), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_469), .B(n_492), .Y(n_603) );
OR2x2_ASAP7_75t_L g627 ( .A(n_469), .B(n_540), .Y(n_627) );
AND2x2_ASAP7_75t_L g640 ( .A(n_469), .B(n_545), .Y(n_640) );
AND2x2_ASAP7_75t_L g680 ( .A(n_469), .B(n_666), .Y(n_680) );
AND2x2_ASAP7_75t_L g687 ( .A(n_469), .B(n_650), .Y(n_687) );
AND2x2_ASAP7_75t_L g717 ( .A(n_469), .B(n_479), .Y(n_717) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_478), .B(n_644), .Y(n_656) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_479), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g594 ( .A(n_479), .B(n_491), .Y(n_594) );
BUFx3_ASAP7_75t_L g602 ( .A(n_479), .Y(n_602) );
OR2x2_ASAP7_75t_L g623 ( .A(n_479), .B(n_505), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_479), .B(n_644), .Y(n_734) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_481), .A2(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g541 ( .A(n_483), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_490), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_491), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g587 ( .A(n_491), .Y(n_587) );
AND2x2_ASAP7_75t_L g650 ( .A(n_491), .B(n_545), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_491), .A2(n_653), .B1(n_655), .B2(n_657), .C(n_658), .Y(n_652) );
AND2x2_ASAP7_75t_L g666 ( .A(n_491), .B(n_540), .Y(n_666) );
AND2x2_ASAP7_75t_L g692 ( .A(n_491), .B(n_576), .Y(n_692) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g572 ( .A(n_492), .B(n_545), .Y(n_572) );
BUFx2_ASAP7_75t_L g706 ( .A(n_492), .Y(n_706) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI32xp33_ASAP7_75t_L g672 ( .A1(n_503), .A2(n_633), .A3(n_647), .B1(n_673), .B2(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
AND2x2_ASAP7_75t_L g613 ( .A(n_504), .B(n_557), .Y(n_613) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_505), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g667 ( .A(n_505), .B(n_557), .Y(n_667) );
AND2x2_ASAP7_75t_L g678 ( .A(n_505), .B(n_570), .Y(n_678) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g579 ( .A(n_506), .B(n_558), .Y(n_579) );
AND2x2_ASAP7_75t_L g583 ( .A(n_506), .B(n_558), .Y(n_583) );
AND2x2_ASAP7_75t_L g618 ( .A(n_506), .B(n_569), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_506), .B(n_527), .Y(n_625) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_506), .A2(n_576), .B(n_587), .C(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g684 ( .A(n_506), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_506), .B(n_517), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_515), .B(n_567), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_515), .B(n_583), .Y(n_673) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g578 ( .A(n_516), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
AND2x2_ASAP7_75t_L g570 ( .A(n_517), .B(n_528), .Y(n_570) );
OR2x2_ASAP7_75t_L g585 ( .A(n_517), .B(n_528), .Y(n_585) );
AND2x2_ASAP7_75t_L g608 ( .A(n_517), .B(n_569), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_517), .Y(n_612) );
AND2x2_ASAP7_75t_L g631 ( .A(n_517), .B(n_568), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_517), .A2(n_596), .B1(n_642), .B2(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_517), .B(n_684), .Y(n_708) );
AND2x2_ASAP7_75t_L g723 ( .A(n_517), .B(n_583), .Y(n_723) );
INVx4_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx3_ASAP7_75t_L g555 ( .A(n_518), .Y(n_555) );
AND2x2_ASAP7_75t_L g597 ( .A(n_518), .B(n_528), .Y(n_597) );
AND2x2_ASAP7_75t_L g599 ( .A(n_518), .B(n_557), .Y(n_599) );
AND3x2_ASAP7_75t_L g661 ( .A(n_518), .B(n_625), .C(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g696 ( .A(n_527), .B(n_568), .Y(n_696) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_528), .B(n_567), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_528), .B(n_608), .C(n_684), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_554), .B1(n_566), .B2(n_571), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_540), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g648 ( .A(n_540), .Y(n_648) );
OAI31xp33_ASAP7_75t_L g664 ( .A1(n_543), .A2(n_665), .A3(n_666), .B(n_667), .Y(n_664) );
AND2x2_ASAP7_75t_L g689 ( .A(n_543), .B(n_576), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_543), .B(n_602), .Y(n_735) );
AND2x2_ASAP7_75t_L g644 ( .A(n_544), .B(n_576), .Y(n_644) );
AND2x2_ASAP7_75t_L g705 ( .A(n_544), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g575 ( .A(n_545), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g633 ( .A(n_545), .Y(n_633) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g654 ( .A(n_555), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_556), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AOI221x1_ASAP7_75t_SL g621 ( .A1(n_557), .A2(n_622), .B1(n_624), .B2(n_626), .C(n_628), .Y(n_621) );
INVx2_ASAP7_75t_L g569 ( .A(n_558), .Y(n_569) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_558), .Y(n_663) );
INVx1_ASAP7_75t_L g651 ( .A(n_566), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_567), .B(n_584), .Y(n_676) );
INVx1_ASAP7_75t_SL g739 ( .A(n_567), .Y(n_739) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g657 ( .A(n_570), .B(n_583), .Y(n_657) );
INVx1_ASAP7_75t_L g725 ( .A(n_571), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_571), .B(n_654), .Y(n_738) );
INVx2_ASAP7_75t_SL g577 ( .A(n_572), .Y(n_577) );
AND2x2_ASAP7_75t_L g620 ( .A(n_572), .B(n_576), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_572), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_572), .B(n_647), .Y(n_674) );
AOI21xp33_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_577), .B(n_578), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_575), .B(n_647), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_575), .B(n_602), .Y(n_743) );
OR2x2_ASAP7_75t_L g615 ( .A(n_576), .B(n_594), .Y(n_615) );
AND2x2_ASAP7_75t_L g714 ( .A(n_576), .B(n_705), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_577), .A2(n_590), .B1(n_595), .B2(n_598), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_577), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g637 ( .A(n_579), .B(n_585), .Y(n_637) );
INVx1_ASAP7_75t_L g701 ( .A(n_579), .Y(n_701) );
AOI311xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_586), .A3(n_588), .B(n_589), .C(n_600), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_584), .A2(n_716), .B1(n_728), .B2(n_731), .C(n_733), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_584), .B(n_739), .Y(n_741) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g638 ( .A(n_586), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_587), .A2(n_629), .B(n_630), .C(n_632), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_SL g697 ( .A1(n_591), .A2(n_593), .B(n_698), .C(n_699), .Y(n_697) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_592), .B(n_666), .Y(n_732) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_595), .A2(n_615), .B1(n_616), .B2(n_619), .C(n_621), .Y(n_614) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g617 ( .A(n_597), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g700 ( .A(n_597), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g658 ( .A1(n_601), .A2(n_659), .B(n_660), .C(n_664), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_602), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_602), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g624 ( .A(n_608), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_612), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g726 ( .A(n_615), .Y(n_726) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_618), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g653 ( .A(n_618), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g730 ( .A(n_618), .Y(n_730) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g671 ( .A(n_620), .B(n_647), .Y(n_671) );
INVx1_ASAP7_75t_SL g665 ( .A(n_627), .Y(n_665) );
INVx1_ASAP7_75t_L g642 ( .A(n_633), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_652), .C(n_668), .Y(n_634) );
AOI322xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .A3(n_639), .B1(n_641), .B2(n_645), .C1(n_649), .C2(n_651), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_636), .A2(n_689), .B(n_690), .C(n_697), .Y(n_688) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_639), .A2(n_660), .B1(n_691), .B2(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g649 ( .A(n_647), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g686 ( .A(n_647), .B(n_687), .Y(n_686) );
AOI32xp33_ASAP7_75t_L g737 ( .A1(n_647), .A2(n_738), .A3(n_739), .B1(n_740), .B2(n_742), .Y(n_737) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g659 ( .A(n_650), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_650), .A2(n_703), .B1(n_707), .B2(n_709), .C(n_712), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_650), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g719 ( .A(n_654), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g729 ( .A(n_654), .B(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g720 ( .A(n_663), .B(n_684), .Y(n_720) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_675), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_685), .B(n_688), .C(n_702), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_696), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g711 ( .A(n_708), .Y(n_711) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_718), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI211xp5_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_724), .B(n_727), .C(n_737), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
endmodule