module fake_jpeg_9445_n_241 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_20),
.Y(n_61)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_44),
.Y(n_58)
);

NOR2xp67_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_1),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_24),
.CON(n_64),
.SN(n_64)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_52),
.Y(n_76)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_59),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_17),
.B1(n_21),
.B2(n_28),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_20),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_68),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_17),
.B1(n_21),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_72),
.B(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_75),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_40),
.C(n_39),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_90),
.C(n_91),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_18),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_96),
.A3(n_57),
.B1(n_25),
.B2(n_34),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_33),
.B(n_18),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_27),
.B(n_34),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_38),
.C(n_36),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_32),
.B(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_33),
.A3(n_25),
.B1(n_22),
.B2(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_103),
.B1(n_114),
.B2(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_112),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_25),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_90),
.C(n_78),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_19),
.B(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_20),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_25),
.A3(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_57),
.B1(n_65),
.B2(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_22),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_119),
.Y(n_132)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_22),
.Y(n_119)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_27),
.B(n_26),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_83),
.B(n_31),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_25),
.C(n_120),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_92),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_85),
.B1(n_96),
.B2(n_81),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_149),
.B1(n_150),
.B2(n_114),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_134),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_23),
.B(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_140),
.Y(n_165)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_30),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_79),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_73),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_106),
.B(n_117),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_105),
.B(n_25),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_148),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_120),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_93),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_93),
.B1(n_49),
.B2(n_87),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_87),
.B1(n_75),
.B2(n_71),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_123),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_124),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_161),
.C(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_174),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_118),
.B1(n_71),
.B2(n_102),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_149),
.B1(n_134),
.B2(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_163),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_173),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_128),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_80),
.B(n_105),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_171),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_29),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_129),
.C(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_16),
.C(n_14),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_99),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_134),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_167),
.B1(n_155),
.B2(n_152),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_144),
.B1(n_133),
.B2(n_138),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_147),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_194),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_129),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_192),
.C(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_168),
.C(n_165),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_132),
.C(n_136),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_142),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_205),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.C(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_206),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_159),
.B1(n_157),
.B2(n_160),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_188),
.B1(n_177),
.B2(n_193),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_169),
.C(n_154),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_169),
.C(n_172),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_166),
.C(n_173),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_144),
.C(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_181),
.B1(n_183),
.B2(n_131),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_196),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_2),
.B(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_2),
.B(n_3),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_219),
.B(n_212),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_204),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_226),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_198),
.Y(n_226)
);

XOR2x1_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_210),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_228),
.B(n_12),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_222),
.A2(n_214),
.B1(n_218),
.B2(n_137),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_4),
.B(n_5),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_4),
.B(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_235),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_4),
.C(n_5),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_231),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_231),
.B(n_9),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_239),
.A2(n_236),
.B(n_237),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_10),
.Y(n_241)
);


endmodule