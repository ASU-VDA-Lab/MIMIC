module fake_jpeg_1212_n_687 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_687);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_687;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_544;
wire n_455;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_13),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_61),
.Y(n_233)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_73),
.Y(n_193)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_78),
.Y(n_203)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_79),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_10),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_80),
.B(n_92),
.Y(n_160)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_11),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_93),
.Y(n_161)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_89),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_90),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_9),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_12),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_45),
.B(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_124),
.Y(n_166)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_20),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_119),
.Y(n_230)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_120),
.Y(n_232)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_123),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_28),
.A2(n_8),
.B(n_18),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_27),
.Y(n_125)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_128),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

BUFx4f_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_13),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_19),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_19),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_34),
.Y(n_132)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_56),
.B1(n_34),
.B2(n_37),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g260 ( 
.A1(n_142),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_40),
.B1(n_34),
.B2(n_37),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_147),
.A2(n_200),
.B1(n_221),
.B2(n_31),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_151),
.B(n_183),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_92),
.A2(n_40),
.B1(n_37),
.B2(n_57),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_93),
.A2(n_40),
.B1(n_37),
.B2(n_57),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_40),
.B1(n_57),
.B2(n_28),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_80),
.B1(n_112),
.B2(n_96),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_156),
.A2(n_165),
.B1(n_188),
.B2(n_191),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_62),
.A2(n_41),
.B1(n_51),
.B2(n_50),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_72),
.A2(n_25),
.B1(n_36),
.B2(n_54),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_167),
.A2(n_187),
.B1(n_224),
.B2(n_32),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_169),
.B(n_182),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_85),
.B(n_25),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_77),
.B(n_54),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_132),
.A2(n_24),
.B1(n_36),
.B2(n_52),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_81),
.A2(n_52),
.B1(n_46),
.B2(n_30),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_110),
.A2(n_41),
.B1(n_51),
.B2(n_50),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_60),
.Y(n_194)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_66),
.A2(n_51),
.B1(n_50),
.B2(n_41),
.Y(n_200)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_71),
.Y(n_205)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_78),
.B(n_24),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_206),
.B(n_207),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_89),
.B(n_33),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_90),
.B(n_46),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_211),
.B(n_213),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_91),
.B(n_28),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_95),
.B(n_35),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_218),
.B(n_3),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_98),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_115),
.B(n_35),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_100),
.A2(n_35),
.B1(n_30),
.B2(n_32),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_101),
.B(n_30),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_222),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_107),
.B(n_14),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_111),
.A2(n_31),
.B1(n_14),
.B2(n_18),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_130),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_114),
.Y(n_226)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_114),
.Y(n_227)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_32),
.B1(n_31),
.B2(n_14),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_234),
.A2(n_248),
.B1(n_281),
.B2(n_287),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_145),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_235),
.B(n_280),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_150),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_236),
.Y(n_343)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_0),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_239),
.B(n_252),
.Y(n_360)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_240),
.Y(n_368)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_241),
.Y(n_373)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_242),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_145),
.A2(n_32),
.B1(n_31),
.B2(n_18),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_243),
.A2(n_250),
.B1(n_265),
.B2(n_269),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_140),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_244),
.Y(n_324)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_245),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_249),
.Y(n_330)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_168),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_251),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_156),
.B(n_0),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_17),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_152),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_256),
.A2(n_229),
.B1(n_135),
.B2(n_195),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_163),
.B(n_161),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_133),
.Y(n_259)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_259),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_179),
.B(n_17),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_261),
.Y(n_354)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_153),
.A2(n_16),
.B1(n_15),
.B2(n_2),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_148),
.Y(n_266)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_266),
.Y(n_380)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_267),
.Y(n_345)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_268),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_155),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_137),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_270),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_185),
.B(n_0),
.C(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_271),
.B(n_244),
.C(n_237),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_173),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_273),
.A2(n_276),
.B1(n_295),
.B2(n_298),
.Y(n_338)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_275),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_147),
.A2(n_223),
.B1(n_142),
.B2(n_200),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_279),
.Y(n_371)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_221),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_282),
.B(n_291),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_286),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_159),
.B(n_3),
.Y(n_285)
);

AND2x2_ASAP7_75t_SL g340 ( 
.A(n_285),
.B(n_290),
.Y(n_340)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_196),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_186),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_288),
.B(n_292),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_289),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_149),
.B(n_5),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_202),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_184),
.B(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_293),
.B(n_302),
.Y(n_335)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_202),
.Y(n_294)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_294),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_165),
.A2(n_5),
.B1(n_6),
.B2(n_191),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_171),
.Y(n_296)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_217),
.A2(n_6),
.B1(n_215),
.B2(n_209),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_141),
.Y(n_299)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_201),
.Y(n_300)
);

INVx11_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_170),
.B(n_180),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_146),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_303),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_217),
.A2(n_198),
.B1(n_209),
.B2(n_189),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_304),
.A2(n_319),
.B1(n_248),
.B2(n_238),
.Y(n_356)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_305),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_138),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_307),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_136),
.A2(n_6),
.B1(n_198),
.B2(n_189),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_309),
.B1(n_313),
.B2(n_317),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_199),
.A2(n_181),
.B1(n_210),
.B2(n_230),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_164),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_212),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_162),
.B(n_232),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_311),
.B(n_315),
.Y(n_369)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_195),
.Y(n_313)
);

AO22x1_ASAP7_75t_SL g314 ( 
.A1(n_176),
.A2(n_208),
.B1(n_228),
.B2(n_203),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_134),
.B(n_168),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_164),
.A2(n_201),
.B(n_228),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_290),
.B(n_310),
.C(n_260),
.Y(n_359)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_136),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_318),
.A2(n_321),
.B1(n_197),
.B2(n_134),
.Y(n_348)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_205),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_323),
.B(n_327),
.Y(n_404)
);

AOI32xp33_ASAP7_75t_L g327 ( 
.A1(n_252),
.A2(n_239),
.A3(n_264),
.B1(n_267),
.B2(n_247),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_154),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_332),
.B(n_355),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_278),
.A2(n_197),
.B1(n_154),
.B2(n_157),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_336),
.A2(n_322),
.B1(n_343),
.B2(n_324),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_260),
.A2(n_164),
.B1(n_157),
.B2(n_212),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_L g406 ( 
.A1(n_350),
.A2(n_352),
.B(n_359),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_320),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_362),
.C(n_370),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_215),
.Y(n_355)
);

AO21x2_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_314),
.B(n_304),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_285),
.B(n_246),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_365),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_272),
.B(n_244),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_290),
.B(n_306),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_271),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_260),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_399),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_382),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_389),
.Y(n_447)
);

OAI22x1_ASAP7_75t_SL g387 ( 
.A1(n_378),
.A2(n_260),
.B1(n_306),
.B2(n_281),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_387),
.A2(n_403),
.B1(n_410),
.B2(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_382),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_390),
.A2(n_402),
.B1(n_409),
.B2(n_417),
.Y(n_441)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_347),
.B(n_262),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_392),
.B(n_413),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_368),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_412),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_242),
.B(n_277),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_395),
.A2(n_426),
.B(n_379),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_332),
.B(n_314),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_396),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_375),
.A2(n_359),
.B(n_344),
.C(n_345),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_398),
.A2(n_380),
.B(n_358),
.C(n_367),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_324),
.B(n_316),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_344),
.A2(n_275),
.B(n_274),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_400),
.A2(n_401),
.B(n_414),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_345),
.A2(n_299),
.B(n_303),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_322),
.B1(n_356),
.B2(n_363),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_338),
.A2(n_305),
.B1(n_301),
.B2(n_294),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_353),
.B(n_263),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_405),
.B(n_416),
.Y(n_457)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_363),
.A2(n_369),
.B1(n_335),
.B2(n_334),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_326),
.A2(n_259),
.B1(n_317),
.B2(n_321),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_368),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_255),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_369),
.A2(n_289),
.B(n_257),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_360),
.B(n_266),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_421),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_327),
.B(n_236),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_335),
.A2(n_251),
.B1(n_245),
.B2(n_313),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_341),
.B(n_241),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_340),
.A2(n_268),
.B1(n_318),
.B2(n_249),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_340),
.B(n_240),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_340),
.A2(n_279),
.B1(n_296),
.B2(n_300),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_422),
.A2(n_424),
.B1(n_430),
.B2(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_423),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_340),
.A2(n_357),
.B1(n_355),
.B2(n_341),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_362),
.A2(n_254),
.B1(n_236),
.B2(n_297),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_352),
.B1(n_349),
.B2(n_377),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_328),
.A2(n_333),
.B(n_370),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_384),
.Y(n_427)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_360),
.B(n_254),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_432),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_328),
.B(n_351),
.C(n_342),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_342),
.C(n_364),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_346),
.A2(n_352),
.B1(n_361),
.B2(n_383),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_351),
.B(n_379),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_434),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_432),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_435),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_413),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_477),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_464),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_442),
.A2(n_453),
.B1(n_461),
.B2(n_465),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_444),
.C(n_459),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_372),
.C(n_349),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_401),
.Y(n_445)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_399),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_449),
.B(n_469),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_404),
.A2(n_361),
.B1(n_339),
.B2(n_367),
.Y(n_450)
);

OAI22x1_ASAP7_75t_L g487 ( 
.A1(n_450),
.A2(n_425),
.B1(n_396),
.B2(n_417),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_416),
.A2(n_377),
.B1(n_383),
.B2(n_371),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_418),
.B(n_374),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_395),
.Y(n_460)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_460),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_416),
.A2(n_371),
.B1(n_339),
.B2(n_337),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_380),
.C(n_358),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_418),
.A2(n_337),
.B1(n_330),
.B2(n_374),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_402),
.A2(n_337),
.B1(n_330),
.B2(n_373),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_468),
.A2(n_470),
.B1(n_422),
.B2(n_420),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_399),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_404),
.A2(n_387),
.B1(n_390),
.B2(n_397),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_373),
.C(n_368),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_400),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_476),
.A2(n_414),
.B1(n_419),
.B2(n_408),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_386),
.B(n_325),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_463),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_481),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_476),
.A2(n_387),
.B1(n_390),
.B2(n_397),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_479),
.A2(n_515),
.B1(n_512),
.B2(n_505),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_463),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_398),
.B(n_406),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_484),
.A2(n_517),
.B(n_439),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_447),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_485),
.B(n_493),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_389),
.Y(n_486)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_486),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_487),
.A2(n_439),
.B1(n_467),
.B2(n_445),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_435),
.B(n_393),
.Y(n_489)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_393),
.Y(n_491)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_437),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_495),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_436),
.B(n_438),
.Y(n_496)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_496),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_437),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_498),
.B(n_503),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_467),
.Y(n_500)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_501),
.B(n_510),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_440),
.B(n_405),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_502),
.B(n_486),
.Y(n_545)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_454),
.A2(n_390),
.B1(n_430),
.B2(n_396),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_505),
.A2(n_508),
.B1(n_511),
.B2(n_512),
.Y(n_550)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_446),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_506),
.B(n_507),
.Y(n_546)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_452),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_509),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_459),
.B(n_424),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_470),
.A2(n_398),
.B1(n_385),
.B2(n_390),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_454),
.A2(n_390),
.B1(n_410),
.B2(n_421),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_441),
.A2(n_403),
.B1(n_426),
.B2(n_415),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_513),
.A2(n_516),
.B1(n_439),
.B2(n_467),
.Y(n_528)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_514),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_441),
.A2(n_453),
.B1(n_456),
.B2(n_460),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_452),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_518),
.A2(n_526),
.B1(n_544),
.B2(n_484),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_444),
.C(n_464),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_520),
.B(n_535),
.C(n_536),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_459),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_523),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_457),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_510),
.B(n_457),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g582 ( 
.A(n_524),
.B(n_532),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_525),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_528),
.A2(n_529),
.B1(n_540),
.B2(n_549),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_511),
.A2(n_473),
.B1(n_450),
.B2(n_467),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_482),
.B(n_443),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_530),
.B(n_533),
.Y(n_583)
);

MAJx2_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_473),
.C(n_462),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_462),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_504),
.B(n_429),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_475),
.C(n_472),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_489),
.B(n_414),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_480),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_492),
.B(n_442),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_542),
.C(n_547),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_516),
.A2(n_431),
.B1(n_471),
.B2(n_466),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_480),
.B(n_472),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_479),
.A2(n_503),
.B1(n_490),
.B2(n_497),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_545),
.B(n_514),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_501),
.B(n_471),
.C(n_451),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_513),
.A2(n_431),
.B1(n_448),
.B2(n_466),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_490),
.A2(n_431),
.B1(n_451),
.B2(n_474),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_551),
.A2(n_478),
.B1(n_481),
.B2(n_487),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_498),
.B(n_474),
.C(n_427),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_554),
.B(n_521),
.C(n_547),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_543),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_564),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_SL g590 ( 
.A(n_558),
.B(n_584),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_559),
.A2(n_560),
.B1(n_570),
.B2(n_572),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_526),
.A2(n_544),
.B1(n_552),
.B2(n_534),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_527),
.Y(n_561)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_543),
.Y(n_562)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_562),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_520),
.B(n_392),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_546),
.Y(n_565)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_565),
.Y(n_599)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_554),
.Y(n_567)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_567),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_555),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_569),
.B(n_571),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_553),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_550),
.A2(n_485),
.B1(n_508),
.B2(n_491),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_528),
.A2(n_517),
.B1(n_509),
.B2(n_494),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_573),
.A2(n_578),
.B1(n_581),
.B2(n_585),
.Y(n_593)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_542),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_575),
.B(n_576),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_483),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_525),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_577),
.Y(n_598)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_579),
.B(n_586),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_530),
.B(n_494),
.C(n_507),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_580),
.B(n_536),
.C(n_535),
.Y(n_587)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g584 ( 
.A(n_523),
.B(n_483),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_548),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_587),
.B(n_595),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_563),
.A2(n_518),
.B(n_539),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_588),
.A2(n_563),
.B(n_559),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_579),
.B(n_522),
.Y(n_591)
);

MAJx2_ASAP7_75t_L g618 ( 
.A(n_591),
.B(n_594),
.C(n_609),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_566),
.B(n_522),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_568),
.B(n_524),
.C(n_533),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_568),
.B(n_549),
.C(n_540),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_597),
.B(n_600),
.C(n_602),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_566),
.B(n_529),
.C(n_537),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_583),
.B(n_538),
.C(n_532),
.Y(n_602)
);

AOI21x1_ASAP7_75t_L g605 ( 
.A1(n_575),
.A2(n_506),
.B(n_499),
.Y(n_605)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_605),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_583),
.B(n_551),
.C(n_499),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_607),
.C(n_608),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_574),
.B(n_458),
.C(n_455),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_455),
.C(n_423),
.Y(n_608)
);

XOR2x2_ASAP7_75t_L g609 ( 
.A(n_558),
.B(n_468),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_580),
.B(n_434),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_569),
.Y(n_619)
);

MAJx2_ASAP7_75t_L g638 ( 
.A(n_613),
.B(n_590),
.C(n_610),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_576),
.Y(n_615)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_615),
.Y(n_640)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_604),
.Y(n_616)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_616),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_592),
.A2(n_560),
.B1(n_557),
.B2(n_567),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_617),
.A2(n_595),
.B1(n_366),
.B2(n_329),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_621),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_584),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_593),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_622),
.B(n_628),
.Y(n_635)
);

OAI221xp5_ASAP7_75t_L g623 ( 
.A1(n_611),
.A2(n_573),
.B1(n_582),
.B2(n_578),
.C(n_581),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_623),
.A2(n_602),
.B(n_609),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_600),
.B(n_606),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_625),
.B(n_632),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_598),
.A2(n_557),
.B1(n_585),
.B2(n_586),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_627),
.A2(n_629),
.B1(n_589),
.B2(n_597),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_598),
.B(n_565),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_596),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_588),
.A2(n_582),
.B(n_391),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_630),
.A2(n_631),
.B(n_590),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_601),
.A2(n_388),
.B(n_412),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_612),
.B(n_433),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_603),
.A2(n_394),
.B1(n_330),
.B2(n_325),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_633),
.A2(n_325),
.B1(n_608),
.B2(n_607),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_638),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_636),
.A2(n_641),
.B(n_646),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_620),
.B(n_610),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_637),
.B(n_649),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_615),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_639),
.B(n_643),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_642),
.B(n_645),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_626),
.B(n_587),
.C(n_591),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_623),
.A2(n_366),
.B(n_329),
.Y(n_646)
);

AOI21x1_ASAP7_75t_L g647 ( 
.A1(n_614),
.A2(n_366),
.B(n_613),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_647),
.B(n_631),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_616),
.B(n_628),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_626),
.B(n_625),
.C(n_624),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_650),
.B(n_618),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_651),
.B(n_617),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_654),
.B(n_656),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_650),
.B(n_624),
.C(n_622),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_636),
.A2(n_614),
.B(n_627),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_657),
.A2(n_661),
.B(n_655),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_658),
.B(n_662),
.Y(n_670)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_659),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_629),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_635),
.B(n_633),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_663),
.B(n_664),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_643),
.B(n_632),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_653),
.A2(n_640),
.B(n_641),
.Y(n_666)
);

AOI21x1_ASAP7_75t_SL g674 ( 
.A1(n_666),
.A2(n_668),
.B(n_669),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_660),
.A2(n_644),
.B(n_651),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_656),
.B(n_635),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_672),
.Y(n_677)
);

CKINVDCx14_ASAP7_75t_R g672 ( 
.A(n_655),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_670),
.A2(n_661),
.B(n_647),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_675),
.A2(n_676),
.B(n_667),
.Y(n_679)
);

NAND2x1_ASAP7_75t_L g676 ( 
.A(n_673),
.B(n_654),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_671),
.B(n_645),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_678),
.B(n_659),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_679),
.B(n_681),
.C(n_676),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_677),
.A2(n_665),
.B(n_646),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_680),
.A2(n_674),
.B(n_642),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_682),
.A2(n_683),
.B(n_630),
.Y(n_684)
);

BUFx24_ASAP7_75t_SL g685 ( 
.A(n_684),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_685),
.A2(n_652),
.B(n_644),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_686),
.B(n_652),
.Y(n_687)
);


endmodule