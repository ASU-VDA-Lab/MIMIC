module fake_netlist_1_5212_n_417 (n_45, n_20, n_2, n_38, n_44, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_12, n_9, n_17, n_14, n_10, n_15, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_417);
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_417;
wire n_117;
wire n_361;
wire n_185;
wire n_57;
wire n_407;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_53;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_54;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_70;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_396;
wire n_168;
wire n_398;
wire n_134;
wire n_233;
wire n_82;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_52;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_56;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_58;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_55;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_414;
wire n_350;
wire n_164;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g52 ( .A(n_16), .Y(n_52) );
INVx1_ASAP7_75t_L g53 ( .A(n_25), .Y(n_53) );
INVxp67_ASAP7_75t_SL g54 ( .A(n_26), .Y(n_54) );
INVx1_ASAP7_75t_L g55 ( .A(n_14), .Y(n_55) );
INVx1_ASAP7_75t_L g56 ( .A(n_19), .Y(n_56) );
CKINVDCx16_ASAP7_75t_R g57 ( .A(n_33), .Y(n_57) );
BUFx3_ASAP7_75t_L g58 ( .A(n_0), .Y(n_58) );
INVx1_ASAP7_75t_L g59 ( .A(n_40), .Y(n_59) );
NOR2xp67_ASAP7_75t_L g60 ( .A(n_5), .B(n_46), .Y(n_60) );
INVxp33_ASAP7_75t_L g61 ( .A(n_22), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_41), .Y(n_62) );
INVx1_ASAP7_75t_L g63 ( .A(n_38), .Y(n_63) );
INVx2_ASAP7_75t_L g64 ( .A(n_8), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_49), .Y(n_65) );
CKINVDCx16_ASAP7_75t_R g66 ( .A(n_50), .Y(n_66) );
CKINVDCx5p33_ASAP7_75t_R g67 ( .A(n_29), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_35), .Y(n_68) );
INVxp33_ASAP7_75t_L g69 ( .A(n_47), .Y(n_69) );
BUFx2_ASAP7_75t_SL g70 ( .A(n_42), .Y(n_70) );
INVxp33_ASAP7_75t_L g71 ( .A(n_3), .Y(n_71) );
INVx2_ASAP7_75t_L g72 ( .A(n_21), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_8), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_15), .Y(n_74) );
INVxp67_ASAP7_75t_SL g75 ( .A(n_39), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_6), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_4), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_43), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_3), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_30), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_36), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_18), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_28), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_31), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_72), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_72), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_79), .Y(n_89) );
AND2x2_ASAP7_75t_L g90 ( .A(n_71), .B(n_0), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_57), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_58), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_72), .Y(n_93) );
OAI21x1_ASAP7_75t_L g94 ( .A1(n_52), .A2(n_27), .B(n_48), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_58), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_58), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_64), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_52), .Y(n_98) );
NOR2xp67_ASAP7_75t_L g99 ( .A(n_84), .B(n_1), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_57), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_66), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_66), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_61), .B(n_1), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_67), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_64), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_69), .B(n_2), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_64), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_81), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_53), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_53), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_102), .B(n_78), .Y(n_111) );
NAND3xp33_ASAP7_75t_L g112 ( .A(n_103), .B(n_73), .C(n_76), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_102), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_87), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_87), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_91), .B(n_63), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_92), .B(n_73), .Y(n_118) );
AND2x4_ASAP7_75t_L g119 ( .A(n_92), .B(n_76), .Y(n_119) );
INVx4_ASAP7_75t_L g120 ( .A(n_109), .Y(n_120) );
OAI21xp33_ASAP7_75t_L g121 ( .A1(n_110), .A2(n_77), .B(n_85), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_88), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_88), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_110), .B(n_68), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_95), .B(n_86), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_98), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_109), .B(n_85), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_104), .B(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_97), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_95), .B(n_83), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_129), .B(n_103), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_120), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
OR2x6_ASAP7_75t_L g143 ( .A(n_118), .B(n_90), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_118), .B(n_106), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_118), .B(n_90), .Y(n_146) );
INVxp67_ASAP7_75t_SL g147 ( .A(n_133), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_135), .A2(n_109), .B(n_96), .C(n_98), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
OR2x2_ASAP7_75t_L g152 ( .A(n_113), .B(n_105), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_114), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_115), .B(n_106), .Y(n_154) );
INVxp67_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
NOR2x1p5_ASAP7_75t_L g156 ( .A(n_111), .B(n_100), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_118), .B(n_108), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_119), .B(n_99), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_124), .Y(n_161) );
NOR3xp33_ASAP7_75t_SL g162 ( .A(n_134), .B(n_77), .C(n_75), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_120), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_119), .B(n_99), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_119), .B(n_105), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_116), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_111), .B(n_96), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_112), .B(n_94), .Y(n_170) );
NAND2x1p5_ASAP7_75t_L g171 ( .A(n_120), .B(n_94), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_143), .A2(n_126), .B1(n_89), .B2(n_127), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_155), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx6_ASAP7_75t_L g179 ( .A(n_140), .Y(n_179) );
INVx6_ASAP7_75t_SL g180 ( .A(n_143), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_172), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_146), .B(n_137), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_152), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_146), .B(n_127), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_143), .B(n_116), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
BUFx12f_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_143), .B(n_122), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_172), .A2(n_117), .B1(n_121), .B2(n_122), .Y(n_195) );
CKINVDCx8_ASAP7_75t_R g196 ( .A(n_146), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_146), .B(n_131), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_139), .A2(n_94), .B(n_131), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_145), .A2(n_128), .B(n_125), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx3_ASAP7_75t_R g206 ( .A(n_165), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_193), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_198), .B(n_160), .Y(n_208) );
AND2x4_ASAP7_75t_SL g209 ( .A(n_200), .B(n_199), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_185), .A2(n_156), .B1(n_152), .B2(n_165), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_193), .B(n_144), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_198), .B(n_149), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_201), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_173), .A2(n_165), .B1(n_154), .B2(n_157), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_201), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_197), .B(n_149), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_174), .A2(n_153), .B1(n_168), .B2(n_163), .Y(n_218) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_202), .A2(n_170), .B(n_148), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_188), .A2(n_165), .B1(n_154), .B2(n_166), .Y(n_220) );
BUFx2_ASAP7_75t_L g221 ( .A(n_180), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_195), .B(n_170), .C(n_162), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_181), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_205), .Y(n_225) );
OR2x6_ASAP7_75t_L g226 ( .A(n_181), .B(n_149), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_205), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_184), .A2(n_169), .B1(n_158), .B2(n_170), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_188), .B(n_153), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_193), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_178), .B(n_163), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_208), .B(n_193), .Y(n_232) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_218), .A2(n_170), .B(n_204), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_215), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_226), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_214), .A2(n_191), .B1(n_180), .B2(n_175), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_210), .A2(n_196), .B1(n_187), .B2(n_192), .C(n_178), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_222), .A2(n_191), .B1(n_180), .B2(n_199), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_222), .A2(n_199), .B1(n_192), .B2(n_203), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_213), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_231), .Y(n_243) );
BUFx4f_ASAP7_75t_SL g244 ( .A(n_207), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_226), .A2(n_203), .B1(n_182), .B2(n_197), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_231), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_226), .A2(n_182), .B1(n_197), .B2(n_200), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_223), .B(n_196), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_218), .A2(n_177), .B(n_189), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_226), .A2(n_197), .B1(n_200), .B2(n_176), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_244), .Y(n_252) );
OAI221xp5_ASAP7_75t_L g253 ( .A1(n_237), .A2(n_220), .B1(n_228), .B2(n_226), .C(n_221), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_238), .A2(n_212), .B1(n_229), .B2(n_208), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_240), .A2(n_212), .B1(n_229), .B2(n_208), .Y(n_255) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_228), .B1(n_221), .B2(n_212), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_232), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_242), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_232), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_243), .A2(n_246), .B1(n_241), .B2(n_234), .C(n_239), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_242), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_241), .B(n_213), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_248), .B(n_212), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
OR2x6_ASAP7_75t_L g267 ( .A(n_236), .B(n_211), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_250), .B(n_216), .Y(n_268) );
OAI321xp33_ASAP7_75t_L g269 ( .A1(n_233), .A2(n_59), .A3(n_55), .B1(n_56), .B2(n_62), .C(n_82), .Y(n_269) );
INVx8_ASAP7_75t_L g270 ( .A(n_232), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_233), .Y(n_271) );
OAI31xp33_ASAP7_75t_L g272 ( .A1(n_253), .A2(n_209), .A3(n_232), .B(n_211), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_264), .B(n_216), .Y(n_273) );
NAND4xp25_ASAP7_75t_SL g274 ( .A(n_252), .B(n_245), .C(n_251), .D(n_247), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g275 ( .A1(n_270), .A2(n_235), .B1(n_207), .B2(n_230), .Y(n_275) );
AND2x2_ASAP7_75t_SL g276 ( .A(n_254), .B(n_235), .Y(n_276) );
INVx5_ASAP7_75t_L g277 ( .A(n_267), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_255), .A2(n_262), .B1(n_260), .B2(n_252), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_258), .B(n_235), .Y(n_279) );
AOI211xp5_ASAP7_75t_SL g280 ( .A1(n_269), .A2(n_230), .B(n_224), .C(n_60), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
OAI31xp33_ASAP7_75t_L g282 ( .A1(n_256), .A2(n_209), .A3(n_211), .B(n_217), .Y(n_282) );
AOI33xp33_ASAP7_75t_L g283 ( .A1(n_261), .A2(n_56), .A3(n_59), .B1(n_62), .B2(n_63), .B3(n_65), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_259), .B(n_225), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_263), .B(n_225), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_260), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_257), .B(n_235), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_268), .A2(n_249), .B(n_227), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_271), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
OAI221xp5_ASAP7_75t_L g294 ( .A1(n_265), .A2(n_70), .B1(n_107), .B2(n_97), .C(n_55), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_267), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_267), .B(n_227), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_270), .B(n_235), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_270), .B(n_209), .Y(n_298) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_276), .B(n_270), .Y(n_299) );
NAND3xp33_ASAP7_75t_SL g300 ( .A(n_280), .B(n_74), .C(n_68), .Y(n_300) );
NAND2xp33_ASAP7_75t_SL g301 ( .A(n_295), .B(n_206), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_281), .B(n_219), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_273), .B(n_217), .Y(n_303) );
AOI22x1_ASAP7_75t_L g304 ( .A1(n_289), .A2(n_65), .B1(n_74), .B2(n_54), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_295), .B(n_224), .Y(n_305) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_276), .B(n_224), .Y(n_306) );
AOI31xp33_ASAP7_75t_L g307 ( .A1(n_278), .A2(n_171), .A3(n_80), .B(n_107), .Y(n_307) );
NAND2xp33_ASAP7_75t_R g308 ( .A(n_295), .B(n_230), .Y(n_308) );
OAI31xp33_ASAP7_75t_L g309 ( .A1(n_274), .A2(n_217), .A3(n_230), .B(n_171), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_295), .B(n_219), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_287), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_279), .B(n_2), .Y(n_313) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_297), .B(n_219), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_292), .B(n_219), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
AND3x1_ASAP7_75t_L g317 ( .A(n_272), .B(n_5), .C(n_6), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_284), .B(n_7), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_294), .A2(n_171), .B(n_125), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
XOR2xp5_ASAP7_75t_L g321 ( .A(n_297), .B(n_9), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_276), .B(n_296), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_282), .A2(n_189), .B(n_177), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_277), .B(n_194), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_285), .B(n_9), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
NAND3xp33_ASAP7_75t_SL g328 ( .A(n_283), .B(n_10), .C(n_11), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_293), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_321), .B(n_10), .Y(n_331) );
OA21x2_ASAP7_75t_SL g332 ( .A1(n_301), .A2(n_272), .B(n_298), .Y(n_332) );
NAND3xp33_ASAP7_75t_SL g333 ( .A(n_309), .B(n_275), .C(n_282), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g334 ( .A1(n_307), .A2(n_290), .B(n_291), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_330), .B(n_277), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_320), .B(n_277), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_299), .B(n_277), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_317), .A2(n_200), .B1(n_197), .B2(n_128), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_301), .A2(n_176), .B(n_186), .C(n_190), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_316), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_324), .A2(n_177), .B(n_194), .Y(n_342) );
AOI31xp33_ASAP7_75t_L g343 ( .A1(n_308), .A2(n_12), .A3(n_13), .B(n_168), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_322), .B(n_12), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_306), .A2(n_200), .B1(n_179), .B2(n_177), .Y(n_346) );
NOR2x1_ASAP7_75t_L g347 ( .A(n_300), .B(n_190), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_328), .A2(n_183), .B1(n_189), .B2(n_194), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_179), .B1(n_176), .B2(n_186), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_302), .B(n_130), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_325), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_327), .B(n_130), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_322), .B(n_17), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_324), .A2(n_194), .B(n_189), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_308), .A2(n_179), .B1(n_186), .B2(n_189), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_303), .B(n_20), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_318), .B(n_141), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_304), .A2(n_138), .B1(n_141), .B2(n_161), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_359), .B(n_311), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_356), .B(n_314), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_333), .A2(n_323), .B(n_326), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_SL g365 ( .A1(n_337), .A2(n_319), .B(n_305), .C(n_311), .Y(n_365) );
OAI21xp33_ASAP7_75t_SL g366 ( .A1(n_343), .A2(n_305), .B(n_311), .Y(n_366) );
NOR2xp33_ASAP7_75t_R g367 ( .A(n_332), .B(n_23), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
HAxp5_ASAP7_75t_SL g369 ( .A(n_338), .B(n_24), .CON(n_369), .SN(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_341), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g371 ( .A(n_344), .B(n_141), .C(n_138), .D(n_159), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_336), .B(n_34), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_345), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_351), .B(n_37), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_346), .B(n_167), .Y(n_375) );
AND2x2_ASAP7_75t_SL g376 ( .A(n_353), .B(n_164), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_355), .B(n_335), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
NAND2xp33_ASAP7_75t_L g379 ( .A(n_334), .B(n_161), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_350), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_366), .B(n_357), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_363), .A2(n_331), .B1(n_348), .B2(n_360), .C(n_349), .Y(n_382) );
XOR2x1_ASAP7_75t_L g383 ( .A(n_367), .B(n_361), .Y(n_383) );
AOI321xp33_ASAP7_75t_L g384 ( .A1(n_364), .A2(n_347), .A3(n_358), .B1(n_349), .B2(n_340), .C(n_342), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_377), .Y(n_385) );
NOR3xp33_ASAP7_75t_L g386 ( .A(n_379), .B(n_354), .C(n_138), .Y(n_386) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_379), .B(n_164), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_373), .Y(n_388) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_371), .A2(n_150), .B(n_44), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_362), .B(n_51), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_376), .A2(n_380), .B1(n_378), .B2(n_375), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_368), .B(n_370), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_376), .B(n_372), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_374), .B(n_365), .Y(n_394) );
NOR2x1p5_ASAP7_75t_L g395 ( .A(n_383), .B(n_369), .Y(n_395) );
NOR2xp33_ASAP7_75t_SL g396 ( .A(n_391), .B(n_393), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_392), .B(n_385), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_384), .B(n_382), .C(n_389), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_390), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g400 ( .A1(n_387), .A2(n_366), .B(n_367), .C(n_381), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_388), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_386), .A2(n_366), .B1(n_381), .B2(n_391), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_381), .A2(n_391), .B1(n_385), .B2(n_388), .C(n_366), .Y(n_403) );
OAI22xp33_ASAP7_75t_SL g404 ( .A1(n_381), .A2(n_394), .B1(n_391), .B2(n_385), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_399), .Y(n_405) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_403), .B(n_400), .C(n_402), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_397), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_397), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_401), .Y(n_409) );
XNOR2xp5_ASAP7_75t_L g410 ( .A(n_405), .B(n_395), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_408), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_409), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_410), .B(n_404), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_411), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_414), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_415), .A2(n_413), .B1(n_406), .B2(n_412), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_416), .A2(n_410), .B1(n_407), .B2(n_398), .C(n_396), .Y(n_417) );
endmodule