module fake_jpeg_8675_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_14),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_35),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_26),
.B1(n_35),
.B2(n_25),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_27),
.B1(n_30),
.B2(n_23),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_29),
.B(n_22),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_58),
.Y(n_80)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_76),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_84),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_55),
.B(n_49),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_26),
.B1(n_41),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_23),
.B1(n_33),
.B2(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_40),
.B1(n_45),
.B2(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_45),
.B1(n_22),
.B2(n_29),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_98),
.B1(n_101),
.B2(n_49),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_46),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_40),
.B1(n_19),
.B2(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_33),
.B1(n_20),
.B2(n_28),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_102),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_131),
.B1(n_93),
.B2(n_79),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_69),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_75),
.C(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_20),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_114),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_124),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_96),
.B(n_39),
.Y(n_149)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_31),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_70),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_101),
.B1(n_81),
.B2(n_76),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_137),
.B1(n_151),
.B2(n_158),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_141),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_93),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_121),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_93),
.B1(n_77),
.B2(n_83),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_130),
.B1(n_117),
.B2(n_24),
.Y(n_192)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_122),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_93),
.B1(n_75),
.B2(n_79),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_147),
.B1(n_143),
.B2(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_95),
.B(n_84),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_149),
.B(n_157),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_107),
.C(n_18),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_98),
.B1(n_89),
.B2(n_86),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_150),
.B(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_86),
.B1(n_87),
.B2(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_104),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_32),
.B(n_87),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_74),
.B1(n_91),
.B2(n_92),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_104),
.A2(n_92),
.B1(n_19),
.B2(n_21),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_120),
.B1(n_119),
.B2(n_106),
.Y(n_172)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_121),
.B(n_123),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_129),
.B(n_115),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_164),
.A2(n_170),
.B(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_175),
.C(n_187),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_185),
.B1(n_192),
.B2(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_173),
.B(n_174),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_106),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_188),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_137),
.B1(n_158),
.B2(n_133),
.Y(n_199)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_183),
.Y(n_214)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_141),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_117),
.B1(n_130),
.B2(n_112),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_51),
.C(n_39),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_39),
.B(n_31),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_144),
.B(n_18),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_191),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_18),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_127),
.B1(n_113),
.B2(n_21),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_28),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_196),
.C(n_0),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_133),
.B(n_28),
.C(n_19),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_139),
.B(n_14),
.C(n_12),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_197),
.A2(n_152),
.B(n_134),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_208),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_207),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_135),
.B1(n_132),
.B2(n_19),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_213),
.B1(n_216),
.B2(n_222),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_132),
.B1(n_24),
.B2(n_32),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_167),
.C(n_191),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_176),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_170),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_3),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_171),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_188),
.B(n_164),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_243),
.B(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_166),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_239),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_190),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_232),
.C(n_236),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_180),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_195),
.C(n_167),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_175),
.C(n_187),
.Y(n_239)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_193),
.B(n_168),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_246),
.B1(n_213),
.B2(n_250),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_189),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_215),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_196),
.C(n_168),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_198),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_235),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_194),
.B(n_184),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_199),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_274),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_221),
.B1(n_205),
.B2(n_211),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_265),
.B1(n_266),
.B2(n_255),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_241),
.B1(n_222),
.B2(n_205),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_266),
.B1(n_228),
.B2(n_246),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_224),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_267),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_226),
.B(n_217),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_265),
.A2(n_268),
.B(n_225),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_212),
.B1(n_218),
.B2(n_216),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_206),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_228),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_220),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_274),
.C(n_273),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_280),
.C(n_282),
.Y(n_298)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_236),
.C(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_248),
.C(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_284),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_229),
.B1(n_245),
.B2(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_234),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_259),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_237),
.B(n_215),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_261),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_263),
.CI(n_262),
.CON(n_292),
.SN(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_285),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_290),
.B1(n_283),
.B2(n_278),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_272),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_276),
.B(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_303),
.C(n_280),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_209),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_257),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_304),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_237),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_289),
.B(n_254),
.Y(n_304)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_294),
.B(n_306),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_287),
.C(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_310),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.C(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_299),
.C(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_317),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_301),
.A2(n_281),
.B1(n_11),
.B2(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_292),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_3),
.C(n_4),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_5),
.C(n_6),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_322),
.B(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_309),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_307),
.B(n_317),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_328),
.A2(n_330),
.B(n_331),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_321),
.B(n_6),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_6),
.B(n_7),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_326),
.B(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_336),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_332),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_329),
.B(n_334),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_325),
.B(n_7),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.B(n_8),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_8),
.B(n_334),
.Y(n_342)
);


endmodule