module fake_jpeg_25221_n_74 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_2),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_40),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_34),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_48)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_1),
.CON(n_39),
.SN(n_39)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_4),
.Y(n_47)
);

CKINVDCx12_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_5),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_34),
.B(n_15),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_52),
.B(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_54),
.B1(n_56),
.B2(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_7),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_18),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_7),
.B(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_9),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_27),
.B1(n_14),
.B2(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_11),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_44),
.B1(n_47),
.B2(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_64),
.B1(n_43),
.B2(n_22),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_63),
.B(n_21),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_59),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_62),
.C(n_60),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_57),
.C(n_61),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_63),
.Y(n_74)
);


endmodule