module real_jpeg_26981_n_7 (n_5, n_4, n_0, n_1, n_2, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_38;
wire n_35;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_58;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_48;
wire n_27;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_0),
.B(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_1),
.A2(n_14),
.B1(n_16),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_3),
.A2(n_14),
.B1(n_16),
.B2(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_3),
.A2(n_22),
.B1(n_49),
.B2(n_55),
.Y(n_59)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_5),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_14),
.B(n_17),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_18),
.B1(n_49),
.B2(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_38),
.Y(n_7)
);

OAI21xp5_ASAP7_75t_SL g8 ( 
.A1(n_9),
.A2(n_29),
.B(n_37),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_19),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_10),
.B(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_18),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_12)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_13),
.A2(n_18),
.B(n_48),
.C(n_49),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_13),
.A2(n_17),
.B1(n_49),
.B2(n_55),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_60),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);


endmodule