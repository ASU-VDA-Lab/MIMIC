module fake_jpeg_9965_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_33),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_16),
.B1(n_31),
.B2(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_15),
.B1(n_24),
.B2(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_19),
.B2(n_27),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_48),
.B1(n_39),
.B2(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_16),
.B1(n_31),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_52),
.B1(n_18),
.B2(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_23),
.B1(n_18),
.B2(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_57),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_76),
.B1(n_43),
.B2(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_61),
.Y(n_85)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_32),
.B1(n_40),
.B2(n_35),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_75),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_32),
.B1(n_20),
.B2(n_21),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_71),
.Y(n_106)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_0),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_30),
.C(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_0),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_0),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_33),
.B1(n_30),
.B2(n_4),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_104),
.B1(n_33),
.B2(n_3),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_1),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_5),
.C(n_6),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_43),
.B1(n_45),
.B2(n_36),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_80),
.B1(n_74),
.B2(n_71),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_25),
.B1(n_33),
.B2(n_30),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_107),
.B(n_109),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_62),
.C(n_79),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_114),
.C(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_110),
.A2(n_118),
.B1(n_98),
.B2(n_6),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_57),
.B1(n_89),
.B2(n_97),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_124),
.B1(n_91),
.B2(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_115),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_77),
.C(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_126),
.B1(n_131),
.B2(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_121),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_81),
.B(n_73),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_81),
.B1(n_73),
.B2(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_116),
.B1(n_109),
.B2(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_69),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_84),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_2),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_2),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_83),
.B(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_104),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_33),
.C(n_3),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_2),
.B(n_5),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_105),
.B(n_103),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_105),
.B(n_99),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_93),
.A3(n_83),
.B1(n_92),
.B2(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_143),
.B1(n_145),
.B2(n_147),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_96),
.B(n_92),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_142),
.C(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_91),
.C(n_96),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_104),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_98),
.B(n_95),
.Y(n_147)
);

OAI21x1_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_130),
.B(n_124),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_7),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_127),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_173),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_145),
.B1(n_163),
.B2(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_167),
.C(n_168),
.Y(n_176)
);

NAND5xp2_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_123),
.C(n_129),
.D(n_12),
.E(n_13),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_153),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_135),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_7),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_155),
.Y(n_185)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_135),
.C(n_142),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_188),
.B1(n_175),
.B2(n_163),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_143),
.B1(n_149),
.B2(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_165),
.B(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_183),
.B(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_146),
.C(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_171),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_164),
.CI(n_160),
.CON(n_199),
.SN(n_199)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_134),
.B1(n_136),
.B2(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_179),
.B(n_144),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_186),
.B(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_10),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_159),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_199),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_161),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_201),
.B(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_161),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_188),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_208),
.C(n_176),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_181),
.B1(n_178),
.B2(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_184),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_12),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_204),
.C(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_176),
.C(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_13),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_227),
.C(n_222),
.Y(n_231)
);

OAI321xp33_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_205),
.A3(n_190),
.B1(n_211),
.B2(n_214),
.C(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_168),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_223),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_231),
.A2(n_199),
.B(n_172),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_229),
.B(n_166),
.Y(n_234)
);

OAI221xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_232),
.B1(n_110),
.B2(n_14),
.C(n_13),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_14),
.Y(n_236)
);


endmodule