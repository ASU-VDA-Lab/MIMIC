module fake_jpeg_10982_n_135 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_4),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_29),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_21),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_3),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_23),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_36),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_22),
.B1(n_20),
.B2(n_14),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_33),
.B1(n_43),
.B2(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_15),
.C(n_12),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_66),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_12),
.C(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_5),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_35),
.B(n_12),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_98)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_71),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_90),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_75),
.B1(n_74),
.B2(n_91),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_62),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_87),
.B(n_90),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_104),
.B(n_89),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_82),
.B(n_86),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_88),
.B1(n_79),
.B2(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_88),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_106),
.B(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_85),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_104),
.C(n_94),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_97),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_113),
.B(n_92),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_104),
.B(n_102),
.Y(n_123)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_107),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_123),
.B(n_117),
.C(n_119),
.D(n_110),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_127),
.B(n_123),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_95),
.B(n_96),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_96),
.Y(n_135)
);


endmodule