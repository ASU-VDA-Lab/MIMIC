module fake_netlist_1_59_n_548 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_548);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_548;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_476;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_163;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_56), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_38), .Y(n_76) );
INVxp33_ASAP7_75t_L g77 ( .A(n_62), .Y(n_77) );
INVxp67_ASAP7_75t_L g78 ( .A(n_12), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_13), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_57), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_49), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_71), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_69), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_52), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_41), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_66), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_30), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_2), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_8), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_18), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_12), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_47), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_22), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_26), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_28), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_32), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_11), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_13), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_31), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_67), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_51), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_61), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_39), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_20), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_53), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_45), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_35), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_21), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_27), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_112), .B(n_0), .Y(n_125) );
OAI21x1_ASAP7_75t_L g126 ( .A1(n_113), .A2(n_34), .B(n_73), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_94), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_98), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_117), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_82), .B(n_1), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_117), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_77), .B(n_1), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_96), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_75), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_107), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_110), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_111), .B(n_2), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_90), .B(n_3), .Y(n_148) );
OR2x2_ASAP7_75t_L g149 ( .A(n_81), .B(n_3), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_78), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_76), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_119), .B(n_4), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_76), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_105), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_95), .B(n_4), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_102), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_128), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_148), .B(n_86), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_157), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_134), .B(n_97), .Y(n_169) );
INVx4_ASAP7_75t_SL g170 ( .A(n_143), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_134), .B(n_97), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_125), .B(n_120), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_128), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_125), .B(n_86), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVxp67_ASAP7_75t_SL g183 ( .A(n_135), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_158), .B(n_91), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_142), .B(n_99), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_149), .A2(n_93), .B1(n_104), .B2(n_99), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_135), .B(n_101), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_128), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g193 ( .A1(n_162), .A2(n_106), .B1(n_89), .B2(n_115), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_156), .B(n_106), .Y(n_194) );
INVx1_ASAP7_75t_SL g195 ( .A(n_147), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_152), .B(n_108), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_156), .B(n_108), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_160), .B(n_88), .Y(n_198) );
BUFx2_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
INVx6_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_132), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_160), .B(n_109), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_152), .B(n_109), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_139), .B(n_88), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_144), .B(n_118), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_132), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_141), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_141), .B(n_115), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_146), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_128), .Y(n_214) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_150), .B(n_114), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_128), .Y(n_218) );
BUFx4f_ASAP7_75t_L g219 ( .A(n_166), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_175), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_211), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_211), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g226 ( .A1(n_193), .A2(n_140), .B1(n_131), .B2(n_130), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_194), .B(n_147), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_211), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_194), .B(n_137), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_194), .B(n_137), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_197), .B(n_155), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_168), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_177), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_166), .Y(n_236) );
INVxp67_ASAP7_75t_SL g237 ( .A(n_166), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_215), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_179), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_164), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_164), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_169), .B(n_145), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_197), .B(n_155), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_197), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_191), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_198), .B(n_149), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_191), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_172), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_198), .B(n_126), .Y(n_253) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_198), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_205), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_186), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_205), .B(n_126), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_195), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_189), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_207), .B(n_161), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_201), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_181), .B(n_126), .Y(n_267) );
NAND2xp33_ASAP7_75t_SL g268 ( .A(n_199), .B(n_89), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_200), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_165), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_217), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_165), .B(n_123), .Y(n_272) );
BUFx4f_ASAP7_75t_L g273 ( .A(n_181), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_207), .B(n_127), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_181), .B(n_123), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_169), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_202), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_173), .Y(n_279) );
BUFx4f_ASAP7_75t_L g280 ( .A(n_223), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_260), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_237), .A2(n_173), .B1(n_187), .B2(n_190), .Y(n_282) );
NAND2xp33_ASAP7_75t_L g283 ( .A(n_224), .B(n_203), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_228), .B(n_196), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_238), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_230), .B(n_176), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_261), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_274), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_261), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_276), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_228), .A2(n_176), .B1(n_196), .B2(n_206), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_228), .A2(n_176), .B1(n_206), .B2(n_213), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_219), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_236), .Y(n_298) );
OAI21x1_ASAP7_75t_SL g299 ( .A1(n_229), .A2(n_209), .B(n_216), .Y(n_299) );
AOI22xp33_ASAP7_75t_SL g300 ( .A1(n_270), .A2(n_208), .B1(n_184), .B2(n_210), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_219), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_227), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_248), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_253), .A2(n_212), .B(n_174), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_275), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_234), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_264), .B(n_151), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_234), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_236), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_219), .A2(n_138), .B1(n_136), .B2(n_133), .Y(n_310) );
OAI21xp33_ASAP7_75t_L g311 ( .A1(n_231), .A2(n_136), .B(n_138), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_275), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_248), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_233), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_264), .B(n_151), .Y(n_315) );
BUFx12f_ASAP7_75t_L g316 ( .A(n_248), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_255), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_255), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_270), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_233), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_251), .A2(n_136), .B1(n_138), .B2(n_159), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_245), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_234), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_240), .A2(n_92), .B1(n_114), .B2(n_123), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_232), .B(n_151), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_245), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_253), .A2(n_182), .B(n_167), .Y(n_327) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_300), .A2(n_279), .B1(n_249), .B2(n_277), .C(n_268), .Y(n_328) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_286), .A2(n_226), .B1(n_280), .B2(n_277), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_327), .A2(n_253), .B(n_259), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_325), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_325), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_286), .A2(n_241), .B1(n_246), .B2(n_273), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_319), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_284), .A2(n_268), .B1(n_250), .B2(n_262), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_297), .B(n_301), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_265), .B1(n_244), .B2(n_225), .C(n_272), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_298), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_281), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_287), .B(n_273), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_280), .A2(n_273), .B1(n_312), .B2(n_305), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_284), .A2(n_252), .B1(n_247), .B2(n_267), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_290), .A2(n_267), .B1(n_259), .B2(n_243), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_295), .B(n_272), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_304), .A2(n_259), .B(n_283), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_316), .B(n_267), .Y(n_349) );
AO221x1_ASAP7_75t_L g350 ( .A1(n_298), .A2(n_258), .B1(n_92), .B2(n_159), .C(n_269), .Y(n_350) );
INVx4_ASAP7_75t_SL g351 ( .A(n_297), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_315), .B(n_263), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_291), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g354 ( .A1(n_282), .A2(n_242), .B1(n_258), .B2(n_235), .C(n_271), .Y(n_354) );
CKINVDCx11_ASAP7_75t_R g355 ( .A(n_316), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_280), .B(n_220), .Y(n_356) );
OAI211xp5_ASAP7_75t_SL g357 ( .A1(n_328), .A2(n_321), .B(n_123), .C(n_127), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_346), .B(n_305), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_329), .A2(n_283), .B1(n_318), .B2(n_293), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_350), .A2(n_311), .B(n_314), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_329), .A2(n_318), .B1(n_314), .B2(n_320), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_339), .A2(n_320), .B1(n_312), .B2(n_324), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_349), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_348), .A2(n_299), .B(n_310), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g365 ( .A1(n_337), .A2(n_301), .B(n_303), .C(n_285), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_344), .B(n_296), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_330), .A2(n_296), .B(n_302), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_334), .A2(n_298), .B1(n_309), .B2(n_302), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_341), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_344), .B(n_288), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_355), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_331), .B(n_288), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_352), .B(n_298), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_343), .A2(n_289), .B(n_292), .Y(n_374) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_353), .A2(n_127), .B1(n_151), .B2(n_235), .C1(n_317), .C2(n_306), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
BUFx4f_ASAP7_75t_SL g377 ( .A(n_336), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_343), .A2(n_185), .B(n_167), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_349), .B(n_309), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_347), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_358), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_366), .B(n_345), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_371), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_376), .B(n_337), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_366), .B(n_345), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_380), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_355), .B(n_127), .C(n_342), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_376), .A2(n_354), .B1(n_338), .B2(n_308), .C(n_323), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_378), .B(n_349), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_370), .B(n_335), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_377), .A2(n_309), .B1(n_288), .B2(n_289), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_370), .B(n_335), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_363), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_380), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_378), .A2(n_338), .B1(n_356), .B2(n_100), .C(n_116), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
NOR2xp33_ASAP7_75t_R g399 ( .A(n_363), .B(n_309), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_380), .B(n_335), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_309), .B1(n_313), .B2(n_351), .Y(n_401) );
NOR2xp33_ASAP7_75t_R g402 ( .A(n_363), .B(n_340), .Y(n_402) );
AOI222xp33_ASAP7_75t_L g403 ( .A1(n_369), .A2(n_351), .B1(n_239), .B2(n_257), .C1(n_242), .C2(n_222), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_373), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_357), .A2(n_313), .B1(n_351), .B2(n_340), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_357), .A2(n_326), .B1(n_322), .B2(n_335), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_381), .B(n_326), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_374), .A2(n_180), .B(n_185), .Y(n_408) );
OAI332xp33_ASAP7_75t_L g409 ( .A1(n_362), .A2(n_121), .A3(n_122), .B1(n_124), .B2(n_9), .B3(n_10), .C1(n_11), .C2(n_14), .Y(n_409) );
OAI21x1_ASAP7_75t_L g410 ( .A1(n_367), .A2(n_182), .B(n_204), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_385), .B(n_391), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_404), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_398), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_384), .B(n_379), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g419 ( .A(n_397), .B(n_375), .C(n_365), .D(n_372), .Y(n_419) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_390), .B(n_360), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_387), .B(n_379), .Y(n_422) );
AOI33xp33_ASAP7_75t_L g423 ( .A1(n_391), .A2(n_368), .A3(n_121), .B1(n_122), .B2(n_124), .B3(n_380), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_387), .B(n_379), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_402), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_383), .B(n_364), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_400), .B(n_364), .Y(n_427) );
AOI31xp33_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_365), .A3(n_374), .B(n_375), .Y(n_428) );
NAND3xp33_ASAP7_75t_SL g429 ( .A(n_403), .B(n_121), .C(n_122), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_392), .B(n_360), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_399), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_408), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_411), .B(n_360), .Y(n_434) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_386), .A2(n_360), .B(n_124), .C(n_159), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_407), .Y(n_436) );
AND2x4_ASAP7_75t_SL g437 ( .A(n_400), .B(n_322), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_409), .B(n_5), .Y(n_438) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_406), .A2(n_257), .B(n_239), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_392), .B(n_5), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_401), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_407), .B(n_6), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_408), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_388), .A2(n_128), .B1(n_129), .B2(n_220), .C(n_221), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_392), .B(n_14), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_393), .B(n_180), .C(n_174), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_394), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_388), .B(n_15), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_438), .A2(n_396), .B1(n_405), .B2(n_394), .C(n_129), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_422), .B(n_400), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_413), .B(n_396), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g455 ( .A1(n_420), .A2(n_129), .B(n_204), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_448), .B(n_410), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_424), .B(n_129), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_418), .B(n_15), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_424), .B(n_129), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_447), .B(n_16), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_431), .Y(n_462) );
AOI21xp33_ASAP7_75t_L g463 ( .A1(n_428), .A2(n_129), .B(n_326), .Y(n_463) );
NAND2xp33_ASAP7_75t_R g464 ( .A(n_431), .B(n_17), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_436), .B(n_322), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_419), .B(n_202), .C(n_24), .D(n_25), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_426), .B(n_445), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_426), .B(n_202), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_427), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_445), .B(n_202), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_415), .B(n_19), .Y(n_474) );
NAND5xp2_ASAP7_75t_SL g475 ( .A(n_420), .B(n_33), .C(n_36), .D(n_37), .E(n_40), .Y(n_475) );
INVx3_ASAP7_75t_SL g476 ( .A(n_416), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_435), .A2(n_266), .B(n_256), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
AOI221x1_ASAP7_75t_L g479 ( .A1(n_441), .A2(n_218), .B1(n_214), .B2(n_192), .C(n_178), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_448), .B(n_42), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_440), .B(n_43), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_414), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_450), .B(n_44), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_417), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_451), .B(n_46), .C(n_48), .D(n_50), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_417), .Y(n_486) );
OAI21x1_ASAP7_75t_L g487 ( .A1(n_479), .A2(n_433), .B(n_444), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_476), .A2(n_442), .B1(n_412), .B2(n_415), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g489 ( .A1(n_461), .A2(n_434), .B1(n_430), .B2(n_429), .C1(n_443), .C2(n_433), .Y(n_489) );
OAI322xp33_ASAP7_75t_L g490 ( .A1(n_457), .A2(n_427), .A3(n_432), .B1(n_423), .B2(n_218), .C1(n_163), .C2(n_214), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_478), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_476), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_468), .A2(n_439), .B(n_446), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_464), .A2(n_449), .B1(n_266), .B2(n_256), .C(n_245), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_453), .B(n_437), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_463), .B(n_486), .C(n_484), .Y(n_496) );
OAI311xp33_ASAP7_75t_L g497 ( .A1(n_452), .A2(n_437), .A3(n_60), .B1(n_63), .C1(n_65), .Y(n_497) );
OAI32xp33_ASAP7_75t_L g498 ( .A1(n_462), .A2(n_54), .A3(n_68), .B1(n_72), .B2(n_74), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_485), .A2(n_266), .B(n_256), .C(n_245), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_466), .B(n_170), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_454), .B(n_170), .C(n_163), .D(n_178), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_467), .A2(n_278), .B1(n_178), .B2(n_192), .Y(n_502) );
NAND2x1_ASAP7_75t_SL g503 ( .A(n_467), .B(n_170), .Y(n_503) );
INVxp67_ASAP7_75t_L g504 ( .A(n_458), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_471), .A2(n_278), .B1(n_192), .B2(n_214), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_459), .B(n_163), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_460), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_471), .B(n_192), .Y(n_509) );
INVxp33_ASAP7_75t_L g510 ( .A(n_494), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_489), .B(n_481), .C(n_455), .D(n_474), .Y(n_511) );
AND2x6_ASAP7_75t_SL g512 ( .A(n_492), .B(n_483), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_499), .A2(n_475), .B(n_472), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_506), .B(n_456), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_491), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_487), .Y(n_516) );
NAND2x1_ASAP7_75t_L g517 ( .A(n_495), .B(n_472), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_488), .B(n_467), .C(n_473), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_508), .B(n_482), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_504), .B(n_469), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_503), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_515), .B(n_509), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_510), .A2(n_499), .B1(n_493), .B2(n_496), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_517), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_510), .A2(n_490), .B(n_501), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g526 ( .A1(n_518), .A2(n_502), .B(n_498), .C(n_507), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_521), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_511), .A2(n_507), .B1(n_502), .B2(n_480), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_SL g529 ( .A1(n_516), .A2(n_505), .B(n_473), .C(n_500), .Y(n_529) );
AOI211xp5_ASAP7_75t_L g530 ( .A1(n_513), .A2(n_497), .B(n_465), .C(n_477), .Y(n_530) );
XOR2x2_ASAP7_75t_L g531 ( .A(n_512), .B(n_278), .Y(n_531) );
NOR2x1p5_ASAP7_75t_L g532 ( .A(n_527), .B(n_516), .Y(n_532) );
AOI22x1_ASAP7_75t_L g533 ( .A1(n_524), .A2(n_521), .B1(n_520), .B2(n_514), .Y(n_533) );
NOR2xp33_ASAP7_75t_R g534 ( .A(n_522), .B(n_519), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_530), .A2(n_529), .B(n_525), .C(n_510), .Y(n_535) );
NAND3xp33_ASAP7_75t_SL g536 ( .A(n_528), .B(n_523), .C(n_525), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_531), .B(n_523), .C(n_526), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_537), .B(n_535), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_536), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_534), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_540), .Y(n_541) );
AND3x4_ASAP7_75t_L g542 ( .A(n_539), .B(n_532), .C(n_533), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_541), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_542), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_543), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_544), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_545), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_547), .A2(n_538), .B(n_546), .Y(n_548) );
endmodule