module fake_aes_5854_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx5_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
OA21x2_ASAP7_75t_L g15 ( .A1(n_8), .A2(n_10), .B(n_12), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
NAND2x1_ASAP7_75t_L g19 ( .A(n_16), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_15), .B(n_14), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_18), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_16), .Y(n_23) );
AOI32xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_17), .A3(n_2), .B1(n_3), .B2(n_4), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
NAND4xp25_ASAP7_75t_L g26 ( .A(n_25), .B(n_21), .C(n_3), .D(n_1), .Y(n_26) );
NOR2xp67_ASAP7_75t_L g27 ( .A(n_26), .B(n_1), .Y(n_27) );
OAI22xp5_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_15), .B1(n_14), .B2(n_9), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_14), .B1(n_7), .B2(n_11), .C(n_6), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
endmodule