module fake_jpeg_22360_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_1),
.B(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_26),
.B1(n_17),
.B2(n_28),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_26),
.B1(n_17),
.B2(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_26),
.B1(n_17),
.B2(n_20),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_26),
.B1(n_36),
.B2(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_21),
.B1(n_25),
.B2(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_89),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_88),
.B1(n_106),
.B2(n_20),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_77),
.B1(n_105),
.B2(n_64),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_91),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_28),
.B1(n_45),
.B2(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_92),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_24),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_34),
.B1(n_45),
.B2(n_38),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_64),
.B1(n_67),
.B2(n_63),
.Y(n_115)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_60),
.B(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_23),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_20),
.B1(n_27),
.B2(n_36),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_24),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_29),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_94),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_50),
.B1(n_29),
.B2(n_19),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_52),
.B(n_53),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_104),
.B(n_82),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_126),
.B1(n_85),
.B2(n_77),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_62),
.B1(n_23),
.B2(n_25),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_62),
.B1(n_23),
.B2(n_29),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_29),
.B(n_30),
.C(n_19),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_121),
.C(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_99),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_105),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_19),
.B1(n_22),
.B2(n_30),
.Y(n_126)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_84),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_21),
.B1(n_33),
.B2(n_19),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_135),
.A2(n_98),
.B1(n_86),
.B2(n_37),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_33),
.B1(n_22),
.B2(n_30),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_78),
.B1(n_75),
.B2(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_138),
.B(n_153),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_139),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_149),
.B1(n_131),
.B2(n_110),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_89),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_150),
.B(n_113),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_87),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_146),
.A2(n_37),
.B(n_34),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_88),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_157),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_108),
.A2(n_97),
.B(n_86),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_34),
.B(n_37),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_93),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_159),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_117),
.B(n_34),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_131),
.B1(n_126),
.B2(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_97),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_22),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_124),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_97),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_122),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_169),
.A2(n_181),
.B(n_191),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_190),
.B1(n_151),
.B2(n_155),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_127),
.C(n_136),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_163),
.C(n_159),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_177),
.B1(n_188),
.B2(n_192),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_110),
.B1(n_115),
.B2(n_119),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_112),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_31),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_115),
.B(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_183),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_115),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_187),
.Y(n_227)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_119),
.B1(n_135),
.B2(n_78),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_119),
.B1(n_59),
.B2(n_56),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_141),
.A2(n_122),
.B1(n_133),
.B2(n_101),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_122),
.B1(n_67),
.B2(n_63),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_155),
.B1(n_160),
.B2(n_137),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_200),
.B(n_34),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_210),
.B1(n_221),
.B2(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_215),
.C(n_172),
.Y(n_237)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_137),
.B1(n_157),
.B2(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_230),
.B1(n_193),
.B2(n_192),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_150),
.B1(n_151),
.B2(n_146),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_224),
.B1(n_225),
.B2(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_216),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_150),
.C(n_146),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_219),
.B(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_169),
.A2(n_139),
.B1(n_59),
.B2(n_56),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_179),
.A2(n_139),
.B1(n_30),
.B2(n_22),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_34),
.B1(n_31),
.B2(n_2),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_176),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_9),
.B(n_15),
.C(n_14),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_235),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_242),
.C(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_239),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_245),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_184),
.C(n_200),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_178),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_184),
.C(n_181),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_177),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_202),
.B1(n_208),
.B2(n_222),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_253),
.A2(n_231),
.B1(n_219),
.B2(n_220),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_211),
.B(n_205),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_267),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_171),
.B1(n_180),
.B2(n_214),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_264),
.A2(n_241),
.B1(n_277),
.B2(n_187),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_171),
.B(n_183),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_168),
.C(n_182),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_168),
.C(n_216),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_275),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_243),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_234),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_229),
.C(n_191),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_257),
.B1(n_242),
.B2(n_241),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_283),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_260),
.B1(n_269),
.B2(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_294),
.B1(n_295),
.B2(n_244),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_265),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_245),
.B(n_253),
.C(n_256),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_288),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_278),
.Y(n_298)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_297),
.B1(n_185),
.B2(n_230),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_264),
.A2(n_266),
.B(n_259),
.C(n_258),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_244),
.B1(n_271),
.B2(n_270),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_254),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_296),
.B(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_299),
.B(n_305),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_273),
.B1(n_279),
.B2(n_209),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_284),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_297),
.B1(n_284),
.B2(n_294),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_268),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_186),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_233),
.B(n_279),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_206),
.C(n_167),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_312),
.C(n_285),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_16),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_185),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_288),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_2),
.C(n_3),
.Y(n_312)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_321),
.B1(n_300),
.B2(n_12),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_282),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_280),
.C(n_294),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_312),
.C(n_303),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_280),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_306),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_294),
.B1(n_284),
.B2(n_12),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_324),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_307),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_327),
.B(n_11),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_313),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_332),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_333),
.C(n_316),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_302),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_336),
.B1(n_340),
.B2(n_4),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_339),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_328),
.A2(n_313),
.B1(n_11),
.B2(n_13),
.Y(n_336)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_327),
.B(n_325),
.Y(n_338)
);

AOI21x1_ASAP7_75t_SL g342 ( 
.A1(n_338),
.A2(n_13),
.B(n_14),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_4),
.Y(n_339)
);

OAI321xp33_ASAP7_75t_L g345 ( 
.A1(n_342),
.A2(n_343),
.A3(n_344),
.B1(n_339),
.B2(n_6),
.C(n_7),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_337),
.A2(n_16),
.B1(n_5),
.B2(n_6),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_341),
.C(n_342),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_4),
.B(n_6),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_347),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_7),
.Y(n_349)
);


endmodule