module fake_jpeg_18005_n_167 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_4),
.B(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_55),
.B1(n_43),
.B2(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_43),
.B1(n_59),
.B2(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_89),
.Y(n_94)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_50),
.B1(n_44),
.B2(n_47),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_57),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_60),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_88),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

BUFx16f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_46),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_0),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_53),
.B1(n_45),
.B2(n_3),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_16),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_114),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_111),
.Y(n_122)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_1),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_2),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_4),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_105),
.B(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_110),
.B1(n_103),
.B2(n_7),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_139),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_116),
.C(n_131),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_145),
.B(n_146),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_124),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_122),
.B1(n_117),
.B2(n_6),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_145),
.C(n_96),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_149),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_151),
.B1(n_23),
.B2(n_9),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_22),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_27),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_21),
.Y(n_158)
);

OAI21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_29),
.B(n_40),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_19),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_17),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_33),
.C(n_38),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_15),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_13),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_34),
.B(n_41),
.Y(n_167)
);


endmodule