module real_jpeg_26434_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_29),
.B1(n_33),
.B2(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_4),
.B(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_4),
.B(n_39),
.C(n_61),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_36),
.B1(n_133),
.B2(n_137),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx8_ASAP7_75t_SL g81 ( 
.A(n_6),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_29),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_53),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_53),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_11),
.A2(n_22),
.B1(n_23),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_66),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_13),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_13),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_100),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_67),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_18),
.B(n_67),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.C(n_54),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_19),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_34),
.B2(n_35),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B(n_27),
.C(n_32),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_22),
.A2(n_23),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_26),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_23),
.B(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

HAxp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.CON(n_28),
.SN(n_28)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_29),
.A2(n_33),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_31),
.B(n_63),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_31),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_42),
.B(n_44),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_36),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_36),
.A2(n_126),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_37),
.B(n_45),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_37),
.A2(n_86),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_39),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_38),
.B(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_40),
.Y(n_134)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_42),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_47),
.B(n_54),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_64),
.B2(n_65),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_59),
.B1(n_63),
.B2(n_109),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_64),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_90),
.B2(n_91),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_89),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_144),
.B(n_148),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_122),
.B(n_143),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_110),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_106),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_118),
.C(n_121),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_129),
.B(n_142),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_128),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_135),
.B(n_141),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);


endmodule