module fake_jpeg_31019_n_261 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_29),
.Y(n_64)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_45),
.Y(n_75)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_16),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_12),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_32),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_23),
.B1(n_14),
.B2(n_31),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_55),
.A2(n_66),
.B1(n_92),
.B2(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_61),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_22),
.B1(n_17),
.B2(n_31),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_73),
.B1(n_81),
.B2(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_64),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_24),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_36),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_32),
.B(n_26),
.C(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_34),
.B1(n_24),
.B2(n_16),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_85),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_25),
.B1(n_23),
.B2(n_17),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_83),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_24),
.B1(n_30),
.B2(n_27),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_38),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_26),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_89),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_44),
.A2(n_33),
.B1(n_29),
.B2(n_17),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_38),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_8),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_30),
.B1(n_27),
.B2(n_5),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_3),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_45),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_39),
.B(n_4),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OR2x2_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_5),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_109),
.B1(n_54),
.B2(n_62),
.Y(n_138)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_67),
.B(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_9),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_69),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_10),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_10),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_95),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_84),
.B1(n_88),
.B2(n_73),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_89),
.B1(n_76),
.B2(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_152),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_133),
.B(n_149),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_90),
.B1(n_55),
.B2(n_58),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_58),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_55),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_147),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_120),
.B(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_66),
.B1(n_90),
.B2(n_82),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_92),
.B1(n_65),
.B2(n_56),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_92),
.B1(n_65),
.B2(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_71),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_86),
.B1(n_77),
.B2(n_71),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_69),
.B1(n_91),
.B2(n_62),
.Y(n_148)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_54),
.B1(n_116),
.B2(n_112),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_101),
.B(n_117),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_123),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_102),
.B(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_176),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_167),
.C(n_126),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_120),
.C(n_119),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_113),
.C(n_105),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_113),
.C(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_134),
.Y(n_186)
);

CKINVDCx10_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_122),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_199),
.B1(n_143),
.B2(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_133),
.B(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_195),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_165),
.B1(n_171),
.B2(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_126),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_197),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_153),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_168),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_203),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_169),
.C(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_205),
.C(n_206),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_159),
.C(n_164),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_186),
.A2(n_174),
.B1(n_175),
.B2(n_145),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_179),
.B1(n_188),
.B2(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_207),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_174),
.C(n_156),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_189),
.C(n_183),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_158),
.B1(n_142),
.B2(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_217),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_222),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_200),
.A2(n_190),
.B(n_158),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_223),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_178),
.C(n_181),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_202),
.C(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_185),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_209),
.B(n_211),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_235),
.C(n_236),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_212),
.C(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_233),
.B1(n_234),
.B2(n_232),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_221),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_218),
.B(n_216),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_243),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_217),
.B(n_216),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_241),
.A2(n_221),
.B(n_235),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_185),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_249),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_215),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_181),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_247),
.A2(n_242),
.B1(n_240),
.B2(n_244),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_154),
.C(n_139),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_173),
.B(n_178),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_248),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_257),
.B1(n_139),
.B2(n_141),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_177),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_256),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_180),
.B(n_254),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_258),
.Y(n_261)
);


endmodule