module fake_jpeg_4763_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_51),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_29),
.B1(n_38),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_59),
.B1(n_33),
.B2(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_58),
.Y(n_72)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_73),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_25),
.B1(n_30),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_80),
.B1(n_26),
.B2(n_50),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_57),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_77),
.B1(n_17),
.B2(n_19),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_25),
.B1(n_27),
.B2(n_20),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_91),
.B1(n_17),
.B2(n_16),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_28),
.C(n_16),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_70),
.C(n_77),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_58),
.B1(n_45),
.B2(n_57),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_32),
.B1(n_1),
.B2(n_3),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_86),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_21),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_46),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_102),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_115),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_108),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_73),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_48),
.B1(n_55),
.B2(n_54),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_106),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_63),
.A2(n_55),
.B1(n_54),
.B2(n_48),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_52),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_70),
.Y(n_123)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_83),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_43),
.B1(n_56),
.B2(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_85),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_81),
.B(n_68),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_132),
.B(n_134),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_89),
.B1(n_92),
.B2(n_81),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_145),
.B1(n_114),
.B2(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_71),
.B(n_68),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_71),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_141),
.C(n_120),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_79),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_65),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_150),
.B(n_1),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_32),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_32),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_94),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_144),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_43),
.B1(n_67),
.B2(n_32),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_142),
.B1(n_122),
.B2(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_0),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_0),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_104),
.B1(n_116),
.B2(n_113),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_154),
.A2(n_172),
.B1(n_178),
.B2(n_180),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_117),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_179),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_182),
.C(n_141),
.Y(n_205)
);

OR2x6_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_96),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_146),
.B(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_138),
.B(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_83),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_136),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_87),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_43),
.B1(n_109),
.B2(n_111),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_122),
.A2(n_111),
.B1(n_1),
.B2(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_126),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_10),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_196),
.B1(n_198),
.B2(n_203),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_182),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_161),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_121),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_205),
.C(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_164),
.A2(n_132),
.B1(n_135),
.B2(n_123),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_168),
.B1(n_156),
.B2(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_132),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_156),
.B1(n_170),
.B2(n_163),
.Y(n_203)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_209),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_175),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_137),
.C(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_212),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_151),
.A2(n_147),
.B1(n_148),
.B2(n_4),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_231),
.Y(n_244)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_151),
.B1(n_152),
.B2(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_166),
.C(n_161),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_188),
.C(n_205),
.Y(n_239)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_236),
.Y(n_238)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_232),
.B(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_173),
.B1(n_159),
.B2(n_176),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_176),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_237),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_169),
.B1(n_148),
.B2(n_6),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_185),
.B(n_4),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_241),
.C(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_203),
.C(n_190),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_197),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_198),
.C(n_186),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_196),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_232),
.B(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_199),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_194),
.C(n_213),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_193),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_228),
.Y(n_279)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_248),
.B1(n_219),
.B2(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_222),
.C(n_214),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_245),
.C(n_241),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_225),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_267),
.B(n_269),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_218),
.B(n_235),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_236),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_268),
.B(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_229),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_224),
.B1(n_233),
.B2(n_217),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_237),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_265),
.B(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_277),
.A2(n_280),
.B(n_283),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_244),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_244),
.C(n_246),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_228),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_238),
.C(n_11),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_261),
.C(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_263),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_292),
.C(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_269),
.B1(n_266),
.B2(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_262),
.B1(n_267),
.B2(n_4),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_9),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_297),
.B(n_298),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_12),
.B1(n_14),
.B2(n_6),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_6),
.C(n_7),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_4),
.B(n_5),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_277),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_302),
.C(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_286),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_278),
.B(n_12),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_292),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_310),
.B(n_15),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_13),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_13),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_303),
.B(n_15),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_313),
.C(n_314),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_308),
.B(n_309),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_15),
.C(n_5),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_5),
.Y(n_318)
);


endmodule