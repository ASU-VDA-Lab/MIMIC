module fake_jpeg_329_n_110 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_23),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_13),
.C(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_38),
.B1(n_35),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_39),
.B1(n_30),
.B2(n_34),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_50),
.B1(n_32),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_41),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_45),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_41),
.B1(n_45),
.B2(n_40),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_44),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_52),
.B(n_40),
.C(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_31),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_41),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_65),
.C(n_14),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_6),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_86),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_2),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_65),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_65),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_92),
.Y(n_97)
);

OAI322xp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_93),
.A3(n_94),
.B1(n_96),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_28),
.C(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_3),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_94)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_79),
.B(n_85),
.C(n_76),
.D(n_84),
.Y(n_99)
);

OA21x2_ASAP7_75t_SL g102 ( 
.A1(n_99),
.A2(n_101),
.B(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);

OAI221xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_98),
.B1(n_79),
.B2(n_95),
.C(n_20),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_98),
.Y(n_110)
);


endmodule