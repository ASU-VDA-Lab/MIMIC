module fake_aes_6920_n_755 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_755);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_755;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g83 ( .A(n_22), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_81), .Y(n_84) );
INVx1_ASAP7_75t_SL g85 ( .A(n_5), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_69), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_29), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_54), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_73), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_52), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_57), .Y(n_92) );
NOR2xp33_ASAP7_75t_L g93 ( .A(n_12), .B(n_19), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_49), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_72), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_50), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_51), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_37), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_40), .Y(n_101) );
INVx1_ASAP7_75t_SL g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_63), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_3), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_1), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_82), .Y(n_107) );
BUFx10_ASAP7_75t_L g108 ( .A(n_32), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_67), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_46), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_58), .Y(n_112) );
BUFx5_ASAP7_75t_L g113 ( .A(n_65), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_79), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_39), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_70), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_24), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_60), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_35), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_17), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_59), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_34), .Y(n_125) );
BUFx10_ASAP7_75t_L g126 ( .A(n_31), .Y(n_126) );
INVxp33_ASAP7_75t_L g127 ( .A(n_61), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_18), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_38), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_53), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_75), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_12), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_28), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_122), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_132), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_135) );
INVx4_ASAP7_75t_L g136 ( .A(n_112), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_127), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_122), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_127), .B(n_3), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_114), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_95), .B(n_4), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_132), .B(n_4), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_95), .Y(n_143) );
INVxp67_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_114), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_118), .A2(n_42), .B(n_77), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_87), .Y(n_152) );
AND2x4_ASAP7_75t_SL g153 ( .A(n_108), .B(n_36), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g154 ( .A1(n_106), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_113), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_119), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_119), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_120), .B(n_6), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_113), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_113), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_87), .B(n_44), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_120), .B(n_43), .Y(n_164) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_128), .A2(n_45), .B(n_76), .Y(n_165) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_128), .A2(n_33), .B(n_74), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_105), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_96), .Y(n_172) );
NOR2x1_ASAP7_75t_L g173 ( .A(n_97), .B(n_30), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_108), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_98), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_88), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_108), .B(n_8), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_101), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_103), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_136), .B(n_126), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_176), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_176), .B(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_136), .B(n_126), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_174), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
XOR2xp5_ASAP7_75t_SL g188 ( .A(n_135), .B(n_130), .Y(n_188) );
INVxp67_ASAP7_75t_SL g189 ( .A(n_137), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_174), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_155), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
BUFx10_ASAP7_75t_L g198 ( .A(n_152), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_136), .B(n_88), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_174), .B(n_89), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_152), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_144), .B(n_89), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_159), .B(n_125), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_141), .B(n_121), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_141), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_175), .B(n_131), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_177), .A2(n_133), .B1(n_131), .B2(n_124), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_175), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_167), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_172), .Y(n_220) );
CKINVDCx6p67_ASAP7_75t_R g221 ( .A(n_177), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_151), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_151), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_172), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_146), .B(n_111), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_164), .Y(n_228) );
INVx5_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
XNOR2xp5_ASAP7_75t_L g230 ( .A(n_154), .B(n_85), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_142), .B(n_104), .Y(n_231) );
NAND3xp33_ASAP7_75t_L g232 ( .A(n_171), .B(n_133), .C(n_124), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_146), .A2(n_93), .B1(n_102), .B2(n_109), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_151), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_153), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_156), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_148), .B(n_117), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_156), .Y(n_238) );
NAND2xp33_ASAP7_75t_SL g239 ( .A(n_139), .B(n_107), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_156), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_153), .Y(n_241) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_150), .A2(n_113), .B(n_115), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_140), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_172), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_161), .B(n_113), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_148), .A2(n_116), .B1(n_110), .B2(n_100), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_156), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_164), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_149), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_189), .B(n_179), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_243), .B(n_179), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_241), .B(n_178), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_249), .B(n_163), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_243), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_198), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_196), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_249), .B(n_178), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_182), .A2(n_157), .B1(n_149), .B2(n_169), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_200), .B(n_157), .Y(n_260) );
NOR2xp33_ASAP7_75t_SL g261 ( .A(n_203), .B(n_198), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_213), .B(n_140), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_242), .A2(n_166), .B(n_165), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_180), .B(n_143), .Y(n_264) );
NOR2xp67_ASAP7_75t_L g265 ( .A(n_232), .B(n_138), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_196), .A2(n_172), .B1(n_164), .B2(n_170), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_182), .A2(n_173), .B1(n_172), .B2(n_164), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_237), .B(n_134), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_185), .Y(n_269) );
BUFx8_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
AND2x6_ASAP7_75t_SL g271 ( .A(n_231), .B(n_138), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g272 ( .A1(n_210), .A2(n_134), .B(n_165), .C(n_166), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_196), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_218), .B(n_92), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_184), .B(n_99), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_181), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_208), .A2(n_170), .B1(n_168), .B2(n_158), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_245), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_218), .B(n_166), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_202), .B(n_166), .Y(n_280) );
OAI221xp5_ASAP7_75t_L g281 ( .A1(n_217), .A2(n_170), .B1(n_168), .B2(n_158), .C(n_156), .Y(n_281) );
OAI22xp33_ASAP7_75t_L g282 ( .A1(n_221), .A2(n_170), .B1(n_168), .B2(n_158), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_221), .A2(n_168), .B1(n_158), .B2(n_170), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_231), .A2(n_165), .B1(n_168), .B2(n_158), .Y(n_285) );
INVxp33_ASAP7_75t_L g286 ( .A(n_230), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_231), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_185), .B(n_165), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_208), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_289) );
INVxp33_ASAP7_75t_L g290 ( .A(n_230), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_206), .B(n_10), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_206), .B(n_11), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_206), .B(n_14), .Y(n_293) );
NAND2xp33_ASAP7_75t_L g294 ( .A(n_208), .B(n_55), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_241), .B(n_48), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_209), .B(n_56), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_209), .B(n_47), .Y(n_297) );
INVx5_ASAP7_75t_L g298 ( .A(n_208), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_208), .A2(n_14), .B1(n_16), .B2(n_21), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_211), .B(n_16), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_245), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_211), .B(n_23), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_228), .B(n_25), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_190), .A2(n_27), .B(n_62), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_190), .B(n_64), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_220), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_204), .B(n_66), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_231), .B(n_78), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_208), .A2(n_68), .B1(n_71), .B2(n_235), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_235), .A2(n_246), .B1(n_233), .B2(n_227), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_228), .B(n_198), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_228), .B(n_239), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_183), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_183), .B(n_216), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_192), .B(n_216), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_248), .B(n_197), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_197), .B(n_229), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_192), .B(n_219), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_193), .B(n_219), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_186), .A2(n_214), .B1(n_215), .B2(n_205), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_193), .B(n_214), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_195), .B(n_215), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_195), .B(n_205), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_201), .B(n_248), .Y(n_324) );
A2O1A1Ixp33_ASAP7_75t_L g325 ( .A1(n_260), .A2(n_201), .B(n_186), .C(n_229), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_280), .A2(n_186), .B(n_226), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_250), .B(n_186), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_303), .A2(n_238), .B(n_236), .C(n_223), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_298), .B(n_197), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_251), .B(n_186), .Y(n_331) );
OA22x2_ASAP7_75t_L g332 ( .A1(n_258), .A2(n_188), .B1(n_242), .B2(n_244), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_279), .A2(n_229), .B(n_226), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_278), .B(n_229), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_298), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_276), .B(n_188), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_301), .B(n_229), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_256), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_298), .B(n_226), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_310), .B(n_226), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_255), .B(n_244), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_288), .A2(n_226), .B(n_197), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_287), .B(n_197), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_SL g346 ( .A1(n_307), .A2(n_244), .B(n_225), .C(n_194), .Y(n_346) );
AOI22xp5_ASAP7_75t_SL g347 ( .A1(n_300), .A2(n_223), .B1(n_238), .B2(n_236), .Y(n_347) );
NOR2xp67_ASAP7_75t_SL g348 ( .A(n_298), .B(n_225), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_269), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_272), .A2(n_222), .B(n_191), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_270), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_263), .A2(n_324), .B(n_257), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_273), .Y(n_353) );
NAND2xp33_ASAP7_75t_SL g354 ( .A(n_276), .B(n_225), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_261), .B(n_222), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_254), .B(n_187), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_300), .A2(n_187), .B1(n_191), .B2(n_194), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_252), .B(n_199), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_252), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_312), .A2(n_199), .B(n_207), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_315), .A2(n_207), .B(n_212), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_289), .A2(n_212), .B1(n_224), .B2(n_234), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_318), .Y(n_364) );
OA22x2_ASAP7_75t_L g365 ( .A1(n_252), .A2(n_224), .B1(n_234), .B2(n_240), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_319), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_321), .A2(n_240), .B(n_247), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_291), .B(n_247), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_322), .A2(n_323), .B(n_262), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_268), .B(n_265), .Y(n_370) );
A2O1A1Ixp33_ASAP7_75t_L g371 ( .A1(n_267), .A2(n_307), .B(n_293), .C(n_292), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_264), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_275), .B(n_308), .C(n_274), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_281), .A2(n_253), .B(n_282), .C(n_289), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_299), .A2(n_309), .B1(n_294), .B2(n_282), .Y(n_375) );
AOI21x1_ASAP7_75t_L g376 ( .A1(n_296), .A2(n_297), .B(n_302), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_285), .A2(n_320), .B(n_275), .C(n_299), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_320), .A2(n_311), .B1(n_305), .B2(n_266), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_283), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_316), .A2(n_317), .B(n_259), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_271), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_284), .Y(n_382) );
NAND2xp33_ASAP7_75t_SL g383 ( .A(n_360), .B(n_286), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_SL g384 ( .A1(n_371), .A2(n_295), .B(n_304), .C(n_306), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_326), .A2(n_266), .B(n_277), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_377), .A2(n_277), .B(n_290), .C(n_370), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_333), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_355), .B(n_364), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_SL g390 ( .A1(n_346), .A2(n_325), .B(n_356), .C(n_331), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_350), .A2(n_352), .B(n_334), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g392 ( .A1(n_372), .A2(n_338), .B(n_373), .C(n_374), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_342), .A2(n_379), .B(n_381), .C(n_369), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
AO31x2_ASAP7_75t_L g395 ( .A1(n_378), .A2(n_358), .A3(n_363), .B(n_327), .Y(n_395) );
AO31x2_ASAP7_75t_L g396 ( .A1(n_358), .A2(n_363), .A3(n_362), .B(n_367), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_337), .B(n_351), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_375), .B(n_347), .C(n_354), .Y(n_398) );
BUFx2_ASAP7_75t_SL g399 ( .A(n_360), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_344), .A2(n_365), .B(n_376), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_360), .B(n_347), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_340), .B(n_332), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_L g403 ( .A1(n_357), .A2(n_335), .B(n_339), .C(n_368), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_336), .Y(n_404) );
BUFx10_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
CKINVDCx11_ASAP7_75t_R g406 ( .A(n_336), .Y(n_406) );
AO31x2_ASAP7_75t_L g407 ( .A1(n_361), .A2(n_380), .A3(n_359), .B(n_382), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_343), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_368), .B1(n_329), .B2(n_349), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_368), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_329), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_345), .A2(n_328), .B(n_330), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_349), .B(n_348), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_341), .B(n_360), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_326), .A2(n_280), .B(n_279), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_326), .A2(n_280), .B(n_279), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_337), .Y(n_417) );
AO31x2_ASAP7_75t_L g418 ( .A1(n_325), .A2(n_377), .A3(n_371), .B(n_352), .Y(n_418) );
OA21x2_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_416), .B(n_415), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
OA21x2_ASAP7_75t_L g421 ( .A1(n_400), .A2(n_398), .B(n_409), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_384), .A2(n_390), .B(n_393), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_392), .A2(n_387), .B(n_398), .Y(n_423) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_403), .A2(n_386), .B(n_389), .Y(n_424) );
OR2x6_ASAP7_75t_L g425 ( .A(n_399), .B(n_409), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_407), .Y(n_426) );
BUFx8_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_404), .B(n_401), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_417), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_412), .A2(n_413), .B(n_385), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_402), .A2(n_413), .B(n_395), .Y(n_432) );
OAI21x1_ASAP7_75t_L g433 ( .A1(n_385), .A2(n_414), .B(n_411), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_394), .B(n_410), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_410), .B(n_408), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_383), .B(n_406), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
OAI21x1_ASAP7_75t_L g439 ( .A1(n_418), .A2(n_396), .B(n_395), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_418), .B(n_395), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_396), .A2(n_392), .B(n_393), .C(n_387), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
OAI21x1_ASAP7_75t_L g444 ( .A1(n_405), .A2(n_391), .B(n_415), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_386), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_384), .A2(n_390), .B(n_415), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_386), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_386), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_386), .B(n_389), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_437), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_449), .B(n_448), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_426), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_427), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_437), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_438), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_429), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_429), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_420), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_420), .B(n_448), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_445), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_445), .Y(n_465) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_446), .A2(n_422), .B(n_431), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_447), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_434), .B(n_432), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_447), .B(n_427), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_426), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_432), .B(n_423), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_419), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_424), .B(n_443), .Y(n_474) );
AO31x2_ASAP7_75t_L g475 ( .A1(n_442), .A2(n_440), .A3(n_443), .B(n_441), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_441), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g477 ( .A1(n_430), .A2(n_436), .B1(n_425), .B2(n_428), .C(n_429), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_427), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_441), .Y(n_479) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_439), .A2(n_444), .B(n_433), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_419), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_439), .A2(n_444), .B(n_419), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_421), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_421), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_458), .B(n_421), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_468), .B(n_421), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_470), .B(n_425), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_469), .B(n_427), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
AND2x4_ASAP7_75t_SL g494 ( .A(n_460), .B(n_425), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_463), .B(n_425), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_455), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_470), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_458), .B(n_435), .Y(n_498) );
NAND2x1_ASAP7_75t_L g499 ( .A(n_461), .B(n_435), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_453), .B(n_435), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_473), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_463), .B(n_465), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_459), .B(n_435), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_461), .B(n_428), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_473), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_481), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_481), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_455), .B(n_428), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_456), .B(n_457), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_456), .B(n_457), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_468), .B(n_471), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_484), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_460), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_460), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_476), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_462), .B(n_467), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_464), .B(n_479), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_460), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_471), .B(n_474), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_462), .B(n_465), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_467), .B(n_474), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_459), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_479), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_482), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_472), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_475), .B(n_464), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_475), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_475), .B(n_486), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_501), .B(n_475), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_519), .B(n_451), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_523), .B(n_475), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_523), .B(n_475), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_526), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_492), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_519), .B(n_454), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_490), .B(n_484), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_504), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_515), .B(n_477), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_502), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_515), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_524), .B(n_478), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_511), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_524), .B(n_485), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_525), .B(n_511), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_501), .B(n_485), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_513), .B(n_485), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_511), .Y(n_554) );
OAI21xp33_ASAP7_75t_L g555 ( .A1(n_532), .A2(n_486), .B(n_483), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_512), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_502), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_502), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_501), .B(n_486), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_513), .B(n_483), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_526), .A2(n_480), .B(n_466), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_512), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_525), .B(n_466), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_497), .B(n_480), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_487), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_487), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_531), .B(n_480), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_491), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_531), .B(n_466), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_491), .B(n_496), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_498), .B(n_497), .Y(n_575) );
AND2x4_ASAP7_75t_SL g576 ( .A(n_515), .B(n_498), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_527), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_515), .B(n_526), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_517), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_517), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_507), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_507), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_518), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_527), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_500), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_533), .B(n_490), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_529), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_522), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_533), .B(n_490), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_499), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_510), .B(n_506), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_499), .B(n_516), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_588), .B(n_533), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_575), .B(n_500), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_549), .B(n_495), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_551), .B(n_493), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_568), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_571), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_574), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_579), .Y(n_604) );
OAI332xp33_ASAP7_75t_L g605 ( .A1(n_565), .A2(n_532), .A3(n_489), .B1(n_495), .B2(n_530), .B3(n_522), .C1(n_528), .C2(n_521), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_554), .B(n_510), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_541), .B(n_493), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_580), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_546), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_588), .B(n_488), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_536), .B(n_489), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_546), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_592), .B(n_510), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_540), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_582), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_556), .B(n_530), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_540), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_592), .B(n_488), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_550), .B(n_508), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_557), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_570), .B(n_520), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_577), .B(n_508), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_570), .B(n_520), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_585), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_576), .B(n_520), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_564), .B(n_506), .Y(n_626) );
NAND2x1_ASAP7_75t_SL g627 ( .A(n_545), .B(n_520), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_576), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_562), .B(n_534), .C(n_514), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_557), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_548), .B(n_494), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_567), .B(n_508), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_573), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_535), .B(n_522), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_572), .B(n_534), .Y(n_635) );
INVx2_ASAP7_75t_SL g636 ( .A(n_547), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_587), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_572), .B(n_534), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_539), .A2(n_494), .B1(n_505), .B2(n_516), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_543), .B(n_509), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_553), .B(n_528), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_535), .B(n_514), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_589), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_544), .B(n_509), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g645 ( .A(n_547), .B(n_516), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_539), .B(n_494), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_590), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_578), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_553), .B(n_528), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_586), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_558), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_611), .B(n_538), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_651), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_637), .A2(n_578), .B(n_534), .C(n_514), .Y(n_655) );
OA21x2_ASAP7_75t_L g656 ( .A1(n_629), .A2(n_555), .B(n_542), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_542), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_637), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_596), .B(n_542), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_633), .B(n_538), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_600), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_601), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_627), .Y(n_663) );
NAND2x1_ASAP7_75t_L g664 ( .A(n_636), .B(n_547), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_642), .A2(n_537), .B1(n_594), .B2(n_593), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_622), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_602), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_605), .B(n_537), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_610), .B(n_566), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_650), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_603), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_604), .Y(n_672) );
NAND5xp2_ASAP7_75t_L g673 ( .A(n_639), .B(n_595), .C(n_591), .D(n_559), .E(n_552), .Y(n_673) );
AOI33xp33_ASAP7_75t_L g674 ( .A1(n_614), .A2(n_559), .A3(n_552), .B1(n_583), .B2(n_563), .B3(n_581), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_610), .B(n_514), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_618), .B(n_560), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_618), .B(n_560), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_648), .A2(n_593), .B(n_595), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_628), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_635), .B(n_566), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_645), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_609), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_609), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_636), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_635), .B(n_561), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_638), .B(n_561), .Y(n_686) );
AOI21xp33_ASAP7_75t_SL g687 ( .A1(n_645), .A2(n_595), .B(n_593), .Y(n_687) );
INVx2_ASAP7_75t_SL g688 ( .A(n_625), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_617), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_608), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_599), .B(n_597), .Y(n_691) );
INVxp67_ASAP7_75t_L g692 ( .A(n_679), .Y(n_692) );
NAND2xp33_ASAP7_75t_SL g693 ( .A(n_674), .B(n_631), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_657), .B(n_642), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_658), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_682), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_668), .B(n_638), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_679), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_665), .A2(n_648), .B1(n_607), .B2(n_646), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_689), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_666), .B(n_613), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_689), .A2(n_634), .B1(n_621), .B2(n_623), .Y(n_702) );
OAI222xp33_ASAP7_75t_L g703 ( .A1(n_664), .A2(n_623), .B1(n_621), .B2(n_646), .C1(n_626), .C2(n_598), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_670), .B(n_615), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_687), .A2(n_640), .B(n_644), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_671), .A2(n_624), .B1(n_647), .B2(n_643), .C(n_616), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_660), .A2(n_606), .B1(n_632), .B2(n_619), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_682), .Y(n_708) );
OAI211xp5_ASAP7_75t_SL g709 ( .A1(n_655), .A2(n_649), .B(n_641), .C(n_630), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_656), .B(n_612), .C(n_620), .Y(n_710) );
INVxp67_ASAP7_75t_L g711 ( .A(n_684), .Y(n_711) );
OAI31xp33_ASAP7_75t_L g712 ( .A1(n_663), .A2(n_620), .A3(n_612), .B(n_558), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_657), .B(n_584), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_661), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g715 ( .A1(n_697), .A2(n_673), .B(n_675), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_710), .B(n_663), .C(n_681), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_695), .B(n_680), .Y(n_717) );
OA211x2_ASAP7_75t_L g718 ( .A1(n_712), .A2(n_664), .B(n_676), .C(n_677), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_714), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_702), .A2(n_688), .B1(n_669), .B2(n_681), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_706), .B(n_675), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_693), .A2(n_678), .B(n_684), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_707), .B(n_662), .Y(n_723) );
NAND2x1_ASAP7_75t_L g724 ( .A(n_700), .B(n_681), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_693), .A2(n_688), .B1(n_653), .B2(n_656), .C(n_691), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_704), .B(n_690), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_699), .A2(n_653), .B1(n_656), .B2(n_659), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_692), .A2(n_656), .B(n_654), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_704), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_698), .A2(n_659), .B(n_686), .C(n_685), .Y(n_730) );
OAI211xp5_ASAP7_75t_L g731 ( .A1(n_702), .A2(n_690), .B(n_661), .C(n_662), .Y(n_731) );
O2A1O1Ixp33_ASAP7_75t_SL g732 ( .A1(n_703), .A2(n_652), .B(n_654), .C(n_672), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_705), .A2(n_652), .B(n_672), .Y(n_733) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_709), .A2(n_667), .B(n_683), .C(n_686), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_711), .B(n_667), .C(n_683), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_701), .B(n_685), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_696), .B(n_708), .Y(n_737) );
AOI21xp33_ASAP7_75t_L g738 ( .A1(n_725), .A2(n_722), .B(n_734), .Y(n_738) );
OA211x2_ASAP7_75t_L g739 ( .A1(n_724), .A2(n_715), .B(n_727), .C(n_728), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_716), .B(n_720), .Y(n_740) );
NOR2xp67_ASAP7_75t_L g741 ( .A(n_731), .B(n_735), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_716), .B(n_732), .C(n_733), .Y(n_742) );
NAND3xp33_ASAP7_75t_SL g743 ( .A(n_740), .B(n_742), .C(n_739), .Y(n_743) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_741), .B(n_718), .Y(n_744) );
NOR2x1_ASAP7_75t_L g745 ( .A(n_738), .B(n_730), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_745), .B(n_729), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_744), .B(n_717), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_747), .B(n_743), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_746), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_749), .Y(n_750) );
OAI22x1_ASAP7_75t_L g751 ( .A1(n_750), .A2(n_748), .B1(n_721), .B2(n_723), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_751), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_752), .B(n_719), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_726), .B(n_736), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_754), .A2(n_737), .B1(n_694), .B2(n_713), .Y(n_755) );
endmodule