module fake_ariane_2483_n_172 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_172);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_172;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_121;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVxp33_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx2_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_0),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_32),
.B1(n_43),
.B2(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_56),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_49),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_55),
.B(n_63),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_63),
.B(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_84),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_69),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_60),
.Y(n_92)
);

AO32x2_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_44),
.A3(n_60),
.B1(n_69),
.B2(n_59),
.Y(n_93)
);

OAI21x1_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_60),
.B(n_58),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_87),
.B(n_72),
.C(n_74),
.Y(n_95)
);

AO31x2_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_68),
.A3(n_67),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_61),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_61),
.B(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_86),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_85),
.B1(n_86),
.B2(n_71),
.Y(n_105)
);

AOI221x1_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_68),
.B1(n_67),
.B2(n_64),
.C(n_62),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_116),
.Y(n_119)
);

NAND2x1_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_114),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NAND4xp25_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_106),
.C(n_110),
.D(n_104),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_112),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_46),
.B1(n_36),
.B2(n_31),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_111),
.B(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_124),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_123),
.B(n_120),
.Y(n_135)
);

AOI222xp33_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_127),
.B1(n_81),
.B2(n_87),
.C1(n_76),
.C2(n_72),
.Y(n_136)
);

OAI221xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_120),
.B1(n_91),
.B2(n_81),
.C(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_1),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_128),
.B(n_126),
.Y(n_139)
);

AOI211xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_89),
.B(n_77),
.C(n_82),
.Y(n_140)
);

AOI311xp33_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_1),
.A3(n_4),
.B(n_5),
.C(n_6),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_4),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_79),
.C(n_77),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_5),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_147),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_136),
.Y(n_151)
);

AOI222xp33_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_125),
.B1(n_121),
.B2(n_107),
.C1(n_88),
.C2(n_8),
.Y(n_152)
);

AND4x1_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_143),
.C(n_144),
.D(n_148),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_94),
.C(n_10),
.Y(n_156)
);

OAI221xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_11),
.B1(n_93),
.B2(n_102),
.C(n_96),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_93),
.C(n_96),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_93),
.C(n_96),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_93),
.C(n_15),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_12),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_154),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_155),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_164),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_163),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_172)
);


endmodule