module fake_aes_5489_n_252 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_252);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_252;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_214;
wire n_204;
wire n_221;
wire n_249;
wire n_185;
wire n_203;
wire n_88;
wire n_244;
wire n_102;
wire n_119;
wire n_141;
wire n_115;
wire n_97;
wire n_167;
wire n_107;
wire n_158;
wire n_114;
wire n_121;
wire n_171;
wire n_94;
wire n_196;
wire n_125;
wire n_192;
wire n_240;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_239;
wire n_137;
wire n_87;
wire n_180;
wire n_104;
wire n_160;
wire n_98;
wire n_154;
wire n_195;
wire n_165;
wire n_146;
wire n_85;
wire n_250;
wire n_237;
wire n_181;
wire n_101;
wire n_215;
wire n_91;
wire n_116;
wire n_108;
wire n_155;
wire n_217;
wire n_209;
wire n_139;
wire n_229;
wire n_230;
wire n_198;
wire n_169;
wire n_193;
wire n_152;
wire n_113;
wire n_241;
wire n_95;
wire n_124;
wire n_156;
wire n_238;
wire n_128;
wire n_129;
wire n_120;
wire n_90;
wire n_206;
wire n_135;
wire n_188;
wire n_247;
wire n_197;
wire n_201;
wire n_242;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_202;
wire n_210;
wire n_142;
wire n_184;
wire n_245;
wire n_191;
wire n_232;
wire n_208;
wire n_200;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_84;
wire n_131;
wire n_112;
wire n_205;
wire n_86;
wire n_143;
wire n_213;
wire n_235;
wire n_243;
wire n_182;
wire n_166;
wire n_162;
wire n_186;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_248;
wire n_231;
wire n_136;
wire n_89;
wire n_176;
wire n_144;
wire n_183;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_83;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_251;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_82;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_246;
wire n_153;
wire n_99;
wire n_132;
wire n_93;
wire n_109;
wire n_151;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_225;
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_50), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_38), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_71), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_36), .Y(n_85) );
BUFx5_ASAP7_75t_L g86 ( .A(n_77), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_51), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_18), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_56), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_57), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_76), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_31), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_37), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_66), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_25), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_28), .Y(n_97) );
BUFx10_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_2), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_22), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_5), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_79), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_80), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_43), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_74), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_69), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_30), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_44), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_21), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
INVx2_ASAP7_75t_SL g114 ( .A(n_29), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_33), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_54), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_40), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_78), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_42), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_55), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_72), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_61), .Y(n_123) );
INVx2_ASAP7_75t_SL g124 ( .A(n_70), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_98), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_91), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_114), .B(n_115), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_91), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_116), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_124), .B(n_1), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_111), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_127), .B(n_84), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_125), .B(n_89), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_133), .B(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_131), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_126), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_143), .B(n_142), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_136), .A2(n_117), .B(n_90), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_138), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_139), .B(n_93), .Y(n_149) );
OAI22xp33_ASAP7_75t_L g150 ( .A1(n_141), .A2(n_129), .B1(n_99), .B2(n_96), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
BUFx5_ASAP7_75t_L g153 ( .A(n_138), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_137), .B(n_97), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_147), .A2(n_152), .B(n_145), .Y(n_155) );
O2A1O1Ixp5_ASAP7_75t_L g156 ( .A1(n_149), .A2(n_88), .B(n_102), .C(n_92), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_148), .A2(n_95), .B(n_94), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_153), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_151), .A2(n_101), .B(n_100), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_153), .B(n_118), .Y(n_160) );
AOI21x1_ASAP7_75t_L g161 ( .A1(n_150), .A2(n_105), .B(n_104), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_154), .B(n_123), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_160), .B(n_119), .Y(n_164) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_156), .A2(n_121), .B(n_120), .Y(n_165) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_108), .B(n_103), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_157), .A2(n_113), .B(n_112), .Y(n_168) );
BUFx12f_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
OAI21x1_ASAP7_75t_SL g170 ( .A1(n_161), .A2(n_3), .B(n_4), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_155), .A2(n_107), .B(n_106), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_162), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_170), .Y(n_173) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_166), .A2(n_132), .B(n_128), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_168), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_171), .A2(n_110), .B(n_109), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_169), .Y(n_177) );
OAI21x1_ASAP7_75t_L g178 ( .A1(n_165), .A2(n_7), .B(n_6), .Y(n_178) );
INVxp67_ASAP7_75t_L g179 ( .A(n_172), .Y(n_179) );
INVx5_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_172), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_172), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_164), .A2(n_122), .B(n_11), .Y(n_183) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_166), .A2(n_12), .B(n_13), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_180), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_173), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_181), .Y(n_187) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_175), .A2(n_14), .B(n_15), .Y(n_188) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_174), .A2(n_16), .B(n_17), .Y(n_189) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_174), .A2(n_19), .B(n_20), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_178), .Y(n_191) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_184), .A2(n_183), .B(n_176), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_182), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_179), .B(n_23), .Y(n_194) );
OR2x6_ASAP7_75t_L g195 ( .A(n_177), .B(n_24), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_173), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_193), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_185), .B(n_26), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_187), .B(n_81), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_197), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_186), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_185), .B(n_27), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_196), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_195), .B(n_75), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_194), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_188), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_191), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_189), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_190), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_192), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_198), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_202), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_201), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_204), .B(n_34), .Y(n_215) );
INVx5_ASAP7_75t_L g216 ( .A(n_199), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_208), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_206), .B(n_39), .Y(n_218) );
INVxp67_ASAP7_75t_L g219 ( .A(n_205), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_203), .Y(n_220) );
OR2x2_ASAP7_75t_L g221 ( .A(n_200), .B(n_41), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_214), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_219), .B(n_211), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_213), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_220), .B(n_207), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_212), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_217), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_216), .B(n_209), .Y(n_228) );
INVxp67_ASAP7_75t_SL g229 ( .A(n_226), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_222), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_225), .B(n_223), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_224), .B(n_215), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_228), .B(n_210), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_229), .B(n_227), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_230), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_234), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_235), .B(n_231), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_237), .A2(n_233), .B(n_232), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_236), .A2(n_221), .B(n_218), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_238), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_239), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_240), .B(n_73), .Y(n_242) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_242), .B(n_241), .Y(n_243) );
XNOR2xp5_ASAP7_75t_L g244 ( .A(n_243), .B(n_46), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_244), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_245), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_246), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_247), .A2(n_52), .B(n_53), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_248), .A2(n_58), .B(n_59), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_249), .A2(n_62), .B(n_63), .Y(n_250) );
NAND2xp33_ASAP7_75t_L g251 ( .A(n_250), .B(n_64), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_251), .A2(n_65), .B1(n_67), .B2(n_68), .Y(n_252) );
endmodule