module fake_jpeg_12415_n_113 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.C(n_36),
.Y(n_37)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_19),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_30),
.B(n_14),
.C(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_13),
.B1(n_20),
.B2(n_25),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_44),
.B1(n_31),
.B2(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_13),
.B1(n_20),
.B2(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_21),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_28),
.B1(n_27),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_43),
.B1(n_42),
.B2(n_49),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_64),
.B(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_51),
.B1(n_43),
.B2(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_28),
.C(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_14),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_75),
.B1(n_52),
.B2(n_42),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_51),
.B1(n_50),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_51),
.B1(n_39),
.B2(n_41),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_77),
.B1(n_65),
.B2(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_56),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_82),
.C(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

AO221x1_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_85),
.B1(n_42),
.B2(n_65),
.C(n_68),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_74),
.B(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_70),
.C(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_95),
.C(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_84),
.B1(n_75),
.B2(n_79),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_70),
.C(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_73),
.Y(n_98)
);

OAI21x1_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_55),
.B(n_53),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_87),
.B1(n_85),
.B2(n_95),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_83),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

OAI22x1_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_97),
.B1(n_100),
.B2(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_8),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_109),
.B(n_10),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_103),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_106),
.B(n_102),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.C(n_2),
.Y(n_112)
);

AOI222xp33_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_96),
.C2(n_15),
.Y(n_113)
);


endmodule