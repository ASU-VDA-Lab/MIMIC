module fake_netlist_6_1971_n_1054 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1054);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1054;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_689;
wire n_354;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_882;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_81),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_12),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_36),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_44),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_61),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_182),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_217),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_48),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_153),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_76),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_189),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_74),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_26),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_67),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_7),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_146),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_88),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_60),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_64),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_187),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_161),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_163),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_120),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_190),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_78),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_4),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_124),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_209),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_107),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_223),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_174),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_3),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_3),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_99),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_105),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_91),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_136),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_183),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_72),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_122),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_89),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_129),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_79),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_137),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_114),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_104),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_113),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_147),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_25),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_97),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_80),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_138),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_109),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_235),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_18),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_215),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_51),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_144),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_166),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_90),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_43),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_127),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_156),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_148),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_59),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_131),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_165),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_24),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_117),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_234),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_195),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_20),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_126),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_13),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_211),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_121),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_13),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_52),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_83),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_37),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_198),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_92),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_95),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_27),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_119),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_204),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_25),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_239),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_238),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_282),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_243),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_250),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_252),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_276),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_245),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_288),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_242),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_309),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_260),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_265),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_326),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_327),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_247),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_248),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_265),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_240),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_241),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_249),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_293),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_281),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_244),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_246),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_253),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_257),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_254),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_251),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_315),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_275),
.B(n_0),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_340),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_255),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_306),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_258),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_256),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_330),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_259),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_261),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_263),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_319),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_268),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_270),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_271),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_262),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_0),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_324),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_264),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

OA21x2_ASAP7_75t_L g398 ( 
.A1(n_373),
.A2(n_292),
.B(n_290),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_343),
.B(n_267),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_347),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_307),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_314),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_367),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_294),
.Y(n_412)
);

BUFx8_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

BUFx8_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_386),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_361),
.B(n_296),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_369),
.B(n_266),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_362),
.B(n_298),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_359),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_394),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_299),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_374),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_273),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_346),
.B(n_273),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_396),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_365),
.B(n_301),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_269),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_395),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_350),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_351),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_352),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_354),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_428),
.B(n_334),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_401),
.B(n_356),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_429),
.Y(n_461)
);

INVx4_ASAP7_75t_SL g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_447),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_360),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_447),
.B(n_338),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_412),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_308),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_414),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_432),
.A2(n_273),
.B1(n_278),
.B2(n_283),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_409),
.A2(n_278),
.B1(n_280),
.B2(n_283),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_421),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_272),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_454),
.B(n_452),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_405),
.Y(n_481)
);

NAND2x1p5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_278),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_274),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_447),
.B(n_277),
.Y(n_487)
);

INVx4_ASAP7_75t_SL g488 ( 
.A(n_437),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_399),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_279),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_399),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_405),
.Y(n_495)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_278),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_411),
.B(n_311),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_454),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_402),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_450),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_321),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_411),
.B(n_284),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_444),
.B(n_438),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_431),
.B(n_328),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_280),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_437),
.B(n_285),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_438),
.B(n_286),
.Y(n_514)
);

NOR2x1p5_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_287),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_439),
.B(n_280),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_426),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_439),
.B(n_289),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_433),
.B(n_291),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_435),
.B(n_280),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_443),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_440),
.B(n_283),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_441),
.B(n_295),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_436),
.A2(n_318),
.B1(n_302),
.B2(n_303),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_404),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_468),
.B(n_430),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_500),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_476),
.A2(n_450),
.B1(n_409),
.B2(n_441),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_478),
.Y(n_535)
);

OAI221xp5_ASAP7_75t_L g536 ( 
.A1(n_504),
.A2(n_419),
.B1(n_424),
.B2(n_427),
.C(n_420),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_460),
.A2(n_409),
.B1(n_448),
.B2(n_446),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_486),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_L g539 ( 
.A(n_463),
.B(n_509),
.Y(n_539)
);

OAI221xp5_ASAP7_75t_L g540 ( 
.A1(n_507),
.A2(n_424),
.B1(n_427),
.B2(n_420),
.C(n_331),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_466),
.A2(n_448),
.B1(n_449),
.B2(n_452),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_520),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_464),
.A2(n_446),
.B1(n_297),
.B2(n_304),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_454),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_505),
.B(n_420),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_473),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_457),
.B(n_451),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_458),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_458),
.B(n_398),
.Y(n_551)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_494),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

BUFx8_ASAP7_75t_L g556 ( 
.A(n_503),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

AO22x2_ASAP7_75t_L g558 ( 
.A1(n_501),
.A2(n_449),
.B1(n_455),
.B2(n_453),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_527),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_493),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_477),
.A2(n_455),
.B1(n_453),
.B2(n_451),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_497),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_526),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_502),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_483),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_510),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_517),
.Y(n_569)
);

BUFx8_ASAP7_75t_L g570 ( 
.A(n_531),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_489),
.Y(n_571)
);

NAND2x1p5_ASAP7_75t_L g572 ( 
.A(n_456),
.B(n_454),
.Y(n_572)
);

BUFx6f_ASAP7_75t_SL g573 ( 
.A(n_469),
.Y(n_573)
);

AND3x1_ASAP7_75t_L g574 ( 
.A(n_490),
.B(n_451),
.C(n_336),
.Y(n_574)
);

AO22x2_ASAP7_75t_L g575 ( 
.A1(n_469),
.A2(n_341),
.B1(n_370),
.B2(n_4),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_454),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_530),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_499),
.A2(n_341),
.B1(n_370),
.B2(n_5),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_515),
.B(n_402),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_434),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_487),
.B(n_434),
.Y(n_583)
);

AO22x2_ASAP7_75t_L g584 ( 
.A1(n_514),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_584)
);

OAI221xp5_ASAP7_75t_L g585 ( 
.A1(n_475),
.A2(n_322),
.B1(n_305),
.B2(n_310),
.C(n_312),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_492),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_518),
.B(n_398),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_521),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_513),
.Y(n_589)
);

NAND2x1p5_ASAP7_75t_L g590 ( 
.A(n_456),
.B(n_398),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_522),
.A2(n_329),
.B1(n_313),
.B2(n_316),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_467),
.B(n_400),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_462),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_594)
);

NOR2xp67_ASAP7_75t_L g595 ( 
.A(n_528),
.B(n_397),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_472),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_525),
.Y(n_597)
);

AO22x2_ASAP7_75t_L g598 ( 
.A1(n_462),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_484),
.B(n_397),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_467),
.B(n_400),
.Y(n_600)
);

OAI221xp5_ASAP7_75t_L g601 ( 
.A1(n_474),
.A2(n_317),
.B1(n_320),
.B2(n_323),
.C(n_332),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_471),
.B(n_283),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_472),
.Y(n_603)
);

AO22x2_ASAP7_75t_L g604 ( 
.A1(n_488),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_488),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_484),
.B(n_418),
.Y(n_606)
);

NAND2x1p5_ASAP7_75t_L g607 ( 
.A(n_519),
.B(n_418),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_471),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_482),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_465),
.Y(n_610)
);

BUFx8_ASAP7_75t_L g611 ( 
.A(n_523),
.Y(n_611)
);

AO22x2_ASAP7_75t_L g612 ( 
.A1(n_512),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_496),
.B(n_333),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_511),
.B(n_335),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_479),
.B(n_418),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_SL g618 ( 
.A(n_553),
.B(n_617),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_553),
.B(n_519),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_532),
.B(n_413),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_567),
.B(n_413),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_SL g622 ( 
.A(n_573),
.B(n_413),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_534),
.B(n_485),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_557),
.B(n_485),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_537),
.B(n_485),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_606),
.B(n_495),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_564),
.B(n_495),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_572),
.B(n_582),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_543),
.B(n_495),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_547),
.B(n_535),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_544),
.B(n_498),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_548),
.B(n_498),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_549),
.B(n_498),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_533),
.B(n_583),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_545),
.B(n_481),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_546),
.B(n_481),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_538),
.B(n_491),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_595),
.B(n_491),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_576),
.B(n_516),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_578),
.B(n_574),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_597),
.B(n_516),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_561),
.B(n_516),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_SL g643 ( 
.A(n_580),
.B(n_523),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_550),
.B(n_516),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_554),
.B(n_523),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_SL g646 ( 
.A(n_613),
.B(n_523),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_555),
.B(n_15),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_563),
.B(n_28),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_566),
.B(n_29),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_559),
.B(n_16),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_577),
.B(n_30),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_577),
.B(n_17),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_568),
.B(n_31),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_560),
.B(n_17),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_614),
.B(n_18),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_569),
.B(n_32),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_591),
.B(n_33),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_539),
.B(n_35),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_581),
.B(n_19),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_589),
.B(n_19),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_607),
.B(n_38),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_542),
.B(n_40),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_565),
.B(n_45),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_599),
.B(n_46),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_610),
.B(n_47),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_552),
.B(n_49),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_571),
.B(n_20),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_SL g668 ( 
.A(n_609),
.B(n_21),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_586),
.B(n_50),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_590),
.B(n_53),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_593),
.B(n_21),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_596),
.B(n_54),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_587),
.B(n_22),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_603),
.B(n_55),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_SL g675 ( 
.A(n_615),
.B(n_22),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_616),
.B(n_56),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_556),
.B(n_57),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_608),
.B(n_58),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_611),
.B(n_62),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_592),
.B(n_63),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_600),
.B(n_65),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_551),
.B(n_23),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_536),
.B(n_541),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_570),
.B(n_66),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_630),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_634),
.B(n_541),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_636),
.A2(n_602),
.B(n_540),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_637),
.A2(n_602),
.B(n_562),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_625),
.A2(n_602),
.B(n_562),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_618),
.B(n_585),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_628),
.B(n_601),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_673),
.B(n_584),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_647),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_668),
.B(n_575),
.C(n_579),
.Y(n_694)
);

AO22x2_ASAP7_75t_L g695 ( 
.A1(n_652),
.A2(n_651),
.B1(n_683),
.B2(n_640),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_635),
.A2(n_605),
.B(n_604),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_651),
.Y(n_697)
);

OAI21x1_ASAP7_75t_SL g698 ( 
.A1(n_650),
.A2(n_594),
.B(n_605),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_584),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_620),
.B(n_24),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_622),
.Y(n_701)
);

NOR4xp25_ASAP7_75t_L g702 ( 
.A(n_654),
.B(n_588),
.C(n_575),
.D(n_579),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_623),
.A2(n_604),
.B(n_598),
.Y(n_703)
);

OAI22x1_ASAP7_75t_L g704 ( 
.A1(n_621),
.A2(n_588),
.B1(n_598),
.B2(n_594),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_619),
.A2(n_670),
.B(n_664),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_672),
.Y(n_706)
);

OA21x2_ASAP7_75t_L g707 ( 
.A1(n_644),
.A2(n_612),
.B(n_558),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_681),
.B(n_558),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_672),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_681),
.A2(n_612),
.B(n_27),
.C(n_26),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_655),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_624),
.B(n_68),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_627),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_675),
.A2(n_75),
.B1(n_77),
.B2(n_82),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_659),
.Y(n_715)
);

OAI21x1_ASAP7_75t_SL g716 ( 
.A1(n_667),
.A2(n_84),
.B(n_85),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_660),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_645),
.A2(n_86),
.B(n_87),
.Y(n_718)
);

OAI21x1_ASAP7_75t_L g719 ( 
.A1(n_629),
.A2(n_93),
.B(n_94),
.Y(n_719)
);

O2A1O1Ixp5_ASAP7_75t_SL g720 ( 
.A1(n_626),
.A2(n_96),
.B(n_98),
.C(n_100),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_646),
.A2(n_638),
.B(n_657),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_661),
.A2(n_101),
.B(n_102),
.C(n_103),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_666),
.B(n_106),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_680),
.A2(n_108),
.B(n_110),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_671),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_658),
.A2(n_116),
.B(n_118),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_633),
.A2(n_123),
.B(n_125),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_631),
.Y(n_728)
);

AOI21xp33_ASAP7_75t_L g729 ( 
.A1(n_632),
.A2(n_128),
.B(n_130),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_SL g730 ( 
.A(n_679),
.B(n_132),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_677),
.B(n_133),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_665),
.Y(n_732)
);

OAI22x1_ASAP7_75t_L g733 ( 
.A1(n_684),
.A2(n_134),
.B1(n_135),
.B2(n_139),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_641),
.Y(n_734)
);

OAI21x1_ASAP7_75t_L g735 ( 
.A1(n_642),
.A2(n_140),
.B(n_142),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_648),
.A2(n_143),
.B1(n_145),
.B2(n_149),
.Y(n_736)
);

AOI21x1_ASAP7_75t_L g737 ( 
.A1(n_639),
.A2(n_150),
.B(n_151),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_662),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_649),
.A2(n_653),
.B(n_656),
.C(n_678),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_L g740 ( 
.A1(n_669),
.A2(n_152),
.B(n_154),
.C(n_155),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_676),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_741)
);

OAI21xp5_ASAP7_75t_L g742 ( 
.A1(n_663),
.A2(n_160),
.B(n_162),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_643),
.B(n_164),
.Y(n_743)
);

AOI21x1_ASAP7_75t_L g744 ( 
.A1(n_721),
.A2(n_674),
.B(n_168),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_706),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_694),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_715),
.B(n_171),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_706),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_685),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_697),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_734),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_686),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_692),
.B(n_177),
.Y(n_753)
);

AO21x2_ASAP7_75t_L g754 ( 
.A1(n_696),
.A2(n_178),
.B(n_179),
.Y(n_754)
);

AND3x1_ASAP7_75t_L g755 ( 
.A(n_702),
.B(n_180),
.C(n_181),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_699),
.B(n_237),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_728),
.Y(n_757)
);

CKINVDCx9p33_ASAP7_75t_R g758 ( 
.A(n_711),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_SL g759 ( 
.A1(n_700),
.A2(n_185),
.B1(n_188),
.B2(n_191),
.Y(n_759)
);

INVxp67_ASAP7_75t_SL g760 ( 
.A(n_693),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_709),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_737),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_717),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_SL g764 ( 
.A(n_709),
.B(n_192),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_695),
.B(n_193),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_719),
.A2(n_735),
.B(n_705),
.Y(n_766)
);

INVx6_ASAP7_75t_L g767 ( 
.A(n_709),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_732),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_695),
.B(n_707),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_732),
.B(n_196),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_738),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_708),
.B(n_199),
.C(n_200),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_703),
.B(n_704),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_687),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_SL g775 ( 
.A1(n_710),
.A2(n_201),
.B(n_202),
.C(n_203),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_689),
.A2(n_205),
.B(n_206),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_740),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_691),
.B(n_233),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_720),
.A2(n_207),
.B(n_208),
.Y(n_779)
);

AO21x2_ASAP7_75t_L g780 ( 
.A1(n_718),
.A2(n_698),
.B(n_716),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_731),
.B(n_210),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_712),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_743),
.Y(n_783)
);

CKINVDCx12_ASAP7_75t_R g784 ( 
.A(n_690),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_732),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_727),
.A2(n_212),
.B(n_216),
.Y(n_786)
);

OAI21x1_ASAP7_75t_SL g787 ( 
.A1(n_739),
.A2(n_218),
.B(n_219),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_723),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_688),
.A2(n_225),
.B(n_226),
.Y(n_789)
);

NOR2x1_ASAP7_75t_R g790 ( 
.A(n_701),
.B(n_227),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_707),
.Y(n_791)
);

AO21x2_ASAP7_75t_L g792 ( 
.A1(n_724),
.A2(n_228),
.B(n_229),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_733),
.Y(n_793)
);

OA21x2_ASAP7_75t_L g794 ( 
.A1(n_742),
.A2(n_230),
.B(n_231),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_726),
.B(n_725),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_714),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_749),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_791),
.Y(n_798)
);

OA21x2_ASAP7_75t_L g799 ( 
.A1(n_774),
.A2(n_714),
.B(n_725),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_784),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_749),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_763),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_766),
.A2(n_722),
.B(n_736),
.Y(n_803)
);

NAND2x1_ASAP7_75t_L g804 ( 
.A(n_787),
.B(n_741),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_791),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_781),
.B(n_730),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_745),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_769),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_751),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_751),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_796),
.A2(n_713),
.B1(n_729),
.B2(n_232),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_773),
.B(n_796),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_771),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_769),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_771),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_784),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_757),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_757),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_785),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_760),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_748),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_748),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_765),
.B(n_793),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_768),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_768),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_750),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_785),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_762),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_778),
.A2(n_793),
.B1(n_765),
.B2(n_772),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_762),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_754),
.Y(n_832)
);

BUFx8_ASAP7_75t_SL g833 ( 
.A(n_761),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_766),
.A2(n_776),
.B(n_789),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_776),
.A2(n_789),
.B(n_744),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_745),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_795),
.A2(n_782),
.B(n_783),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_782),
.B(n_756),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_768),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_745),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_SL g841 ( 
.A1(n_792),
.A2(n_794),
.B1(n_787),
.B2(n_770),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_753),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_758),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_754),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_783),
.B(n_770),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_754),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_753),
.B(n_756),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_747),
.B(n_770),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_780),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_780),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_744),
.A2(n_786),
.B(n_779),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_785),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_777),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_755),
.B(n_785),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_822),
.B(n_761),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_845),
.B(n_785),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_824),
.B(n_759),
.Y(n_857)
);

BUFx10_ASAP7_75t_L g858 ( 
.A(n_800),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_822),
.B(n_780),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_816),
.B(n_790),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_827),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_824),
.B(n_746),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_847),
.B(n_788),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_833),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_845),
.B(n_752),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_829),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_843),
.B(n_767),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_843),
.B(n_767),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_R g869 ( 
.A(n_854),
.B(n_794),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_838),
.B(n_767),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_829),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_848),
.B(n_764),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_828),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_831),
.Y(n_874)
);

XNOR2xp5_ASAP7_75t_L g875 ( 
.A(n_830),
.B(n_794),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_845),
.B(n_792),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_802),
.Y(n_877)
);

NAND2xp33_ASAP7_75t_R g878 ( 
.A(n_854),
.B(n_794),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_842),
.B(n_792),
.Y(n_879)
);

CKINVDCx11_ASAP7_75t_R g880 ( 
.A(n_819),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_R g881 ( 
.A(n_852),
.B(n_764),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_797),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_R g883 ( 
.A(n_852),
.B(n_836),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_831),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_812),
.B(n_775),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_819),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_845),
.B(n_852),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_812),
.B(n_820),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_R g889 ( 
.A(n_799),
.B(n_836),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_837),
.B(n_841),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_819),
.B(n_810),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_807),
.B(n_836),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_R g893 ( 
.A(n_799),
.B(n_807),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_797),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_825),
.B(n_826),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_819),
.B(n_810),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_807),
.B(n_840),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_R g898 ( 
.A(n_840),
.B(n_819),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_798),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_840),
.B(n_839),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_R g901 ( 
.A(n_799),
.B(n_821),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_798),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_866),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_879),
.B(n_814),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_860),
.B(n_801),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_871),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_874),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_884),
.B(n_808),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_899),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_876),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_902),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_877),
.B(n_808),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_888),
.B(n_817),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_900),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_859),
.B(n_814),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_887),
.B(n_805),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_875),
.B(n_850),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_882),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_894),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_875),
.B(n_849),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_873),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_892),
.B(n_850),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_900),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_861),
.B(n_817),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_885),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_870),
.B(n_818),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_891),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_897),
.Y(n_928)
);

INVxp67_ASAP7_75t_SL g929 ( 
.A(n_889),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_891),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_890),
.B(n_849),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_896),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_892),
.B(n_818),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_856),
.B(n_846),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_883),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_896),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_907),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_903),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_928),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_929),
.B(n_832),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_925),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_928),
.A2(n_863),
.B1(n_865),
.B2(n_868),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_921),
.B(n_862),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_922),
.B(n_832),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_903),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_930),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_930),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_922),
.B(n_844),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_904),
.B(n_846),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_931),
.A2(n_834),
.B(n_851),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_914),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_934),
.B(n_844),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_907),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_909),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_905),
.B(n_858),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_906),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_917),
.A2(n_872),
.B1(n_857),
.B2(n_806),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_906),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_951),
.B(n_910),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_939),
.B(n_910),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_943),
.B(n_941),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_944),
.B(n_917),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_951),
.B(n_934),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_944),
.B(n_920),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_939),
.B(n_931),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_951),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_937),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_948),
.B(n_920),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_952),
.B(n_914),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_937),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_953),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_914),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_953),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_940),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_965),
.A2(n_942),
.B1(n_957),
.B2(n_878),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_967),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_963),
.B(n_948),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_SL g978 ( 
.A(n_960),
.B(n_867),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_961),
.A2(n_869),
.B1(n_955),
.B2(n_947),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_970),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_963),
.Y(n_981)
);

NOR2x1_ASAP7_75t_L g982 ( 
.A(n_976),
.B(n_864),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_980),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_974),
.B(n_962),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_981),
.B(n_964),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_979),
.B(n_968),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_978),
.A2(n_947),
.B1(n_946),
.B2(n_806),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_977),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_982),
.A2(n_975),
.B1(n_977),
.B2(n_935),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_985),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_984),
.B(n_972),
.Y(n_992)
);

OAI32xp33_ASAP7_75t_L g993 ( 
.A1(n_988),
.A2(n_971),
.A3(n_959),
.B1(n_973),
.B2(n_949),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_990),
.A2(n_987),
.B1(n_986),
.B2(n_935),
.Y(n_994)
);

NOR2x1_ASAP7_75t_R g995 ( 
.A(n_991),
.B(n_864),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_989),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_996),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_995),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_994),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_994),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_998),
.B(n_993),
.C(n_992),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_999),
.B(n_924),
.Y(n_1002)
);

NAND4xp25_ASAP7_75t_L g1003 ( 
.A(n_1000),
.B(n_946),
.C(n_855),
.D(n_913),
.Y(n_1003)
);

NOR4xp25_ASAP7_75t_L g1004 ( 
.A(n_997),
.B(n_966),
.C(n_811),
.D(n_973),
.Y(n_1004)
);

NAND4xp25_ASAP7_75t_L g1005 ( 
.A(n_998),
.B(n_946),
.C(n_940),
.D(n_926),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_972),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_1000),
.B(n_959),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_1001),
.A2(n_1007),
.B1(n_1005),
.B2(n_1003),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_1002),
.B(n_966),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_1004),
.A2(n_804),
.B(n_927),
.C(n_932),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_1006),
.B(n_804),
.C(n_936),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_1001),
.A2(n_947),
.B1(n_936),
.B2(n_932),
.Y(n_1012)
);

NAND5xp2_ASAP7_75t_SL g1013 ( 
.A(n_1001),
.B(n_969),
.C(n_912),
.D(n_947),
.E(n_915),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_1001),
.B(n_947),
.C(n_912),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1008),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_1014),
.A2(n_930),
.B1(n_856),
.B2(n_880),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_1012),
.B(n_933),
.C(n_954),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

CKINVDCx12_ASAP7_75t_R g1019 ( 
.A(n_1013),
.Y(n_1019)
);

NAND4xp75_ASAP7_75t_L g1020 ( 
.A(n_1010),
.B(n_954),
.C(n_909),
.D(n_911),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_1018),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_1016),
.B(n_1011),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_SL g1023 ( 
.A(n_1019),
.B(n_898),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_1017),
.B(n_930),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_1020),
.B(n_881),
.C(n_949),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_1015),
.B(n_930),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_SL g1027 ( 
.A(n_1015),
.B(n_958),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1021),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1026),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_1027),
.Y(n_1030)
);

OAI221xp5_ASAP7_75t_R g1031 ( 
.A1(n_1023),
.A2(n_901),
.B1(n_893),
.B2(n_930),
.C(n_886),
.Y(n_1031)
);

XNOR2xp5_ASAP7_75t_L g1032 ( 
.A(n_1022),
.B(n_916),
.Y(n_1032)
);

INVxp67_ASAP7_75t_SL g1033 ( 
.A(n_1024),
.Y(n_1033)
);

AO22x2_ASAP7_75t_L g1034 ( 
.A1(n_1025),
.A2(n_956),
.B1(n_945),
.B2(n_938),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_1023),
.B(n_958),
.C(n_956),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1030),
.B(n_945),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1028),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1033),
.A2(n_895),
.B1(n_923),
.B2(n_916),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_SL g1039 ( 
.A(n_1029),
.B(n_1035),
.C(n_1031),
.Y(n_1039)
);

XNOR2xp5_ASAP7_75t_L g1040 ( 
.A(n_1032),
.B(n_916),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_1037),
.Y(n_1041)
);

NOR2xp67_ASAP7_75t_L g1042 ( 
.A(n_1039),
.B(n_1034),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1036),
.Y(n_1043)
);

XNOR2xp5_ASAP7_75t_L g1044 ( 
.A(n_1040),
.B(n_1034),
.Y(n_1044)
);

AOI31xp33_ASAP7_75t_L g1045 ( 
.A1(n_1043),
.A2(n_1038),
.A3(n_923),
.B(n_911),
.Y(n_1045)
);

AOI31xp33_ASAP7_75t_L g1046 ( 
.A1(n_1044),
.A2(n_938),
.A3(n_809),
.B(n_915),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_1046),
.A2(n_1041),
.B(n_1042),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_1045),
.A2(n_809),
.B(n_919),
.C(n_813),
.Y(n_1048)
);

OAI22x1_ASAP7_75t_L g1049 ( 
.A1(n_1047),
.A2(n_919),
.B1(n_918),
.B2(n_908),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1048),
.A2(n_918),
.B1(n_908),
.B2(n_823),
.Y(n_1050)
);

OAI222xp33_ASAP7_75t_L g1051 ( 
.A1(n_1049),
.A2(n_823),
.B1(n_815),
.B2(n_813),
.C1(n_904),
.C2(n_853),
.Y(n_1051)
);

INVxp67_ASAP7_75t_SL g1052 ( 
.A(n_1050),
.Y(n_1052)
);

OAI221xp5_ASAP7_75t_R g1053 ( 
.A1(n_1052),
.A2(n_950),
.B1(n_803),
.B2(n_851),
.C(n_835),
.Y(n_1053)
);

AOI211xp5_ASAP7_75t_L g1054 ( 
.A1(n_1053),
.A2(n_1051),
.B(n_950),
.C(n_815),
.Y(n_1054)
);


endmodule