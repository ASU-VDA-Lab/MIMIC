module real_jpeg_18835_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_0),
.B(n_17),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_2),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_6),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_6),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_6),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_6),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_45),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_6),
.B(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_7),
.Y(n_128)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_7),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_8),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_8),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_8),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_8),
.B(n_275),
.Y(n_274)
);

AND2x4_ASAP7_75t_SL g278 ( 
.A(n_8),
.B(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

AND2x4_ASAP7_75t_SL g25 ( 
.A(n_10),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_30),
.Y(n_29)
);

NAND2x1p5_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

NAND2x1_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_10),
.B(n_60),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_12),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_12),
.B(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_72),
.B(n_216),
.C(n_322),
.D(n_339),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_174),
.C(n_197),
.Y(n_18)
);

AND2x4_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_151),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_20),
.B(n_151),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.C(n_112),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_21),
.B(n_87),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_61),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_22),
.B(n_62),
.C(n_73),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_47),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_23),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_23)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_32),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_64),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_25),
.B(n_90),
.C(n_96),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_25),
.A2(n_64),
.B1(n_140),
.B2(n_228),
.Y(n_308)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_41),
.B(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_33),
.C(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_29),
.A2(n_41),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_29),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_32),
.B(n_33),
.C(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_33),
.A2(n_38),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_33),
.A2(n_38),
.B1(n_68),
.B2(n_69),
.Y(n_335)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_38),
.B(n_80),
.C(n_103),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g339 ( 
.A(n_38),
.B(n_69),
.C(n_206),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_39),
.B(n_47),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_40),
.Y(n_271)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_41),
.B(n_76),
.C(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_41),
.A2(n_76),
.B1(n_118),
.B2(n_133),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_44),
.B(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_44),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_44),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_44),
.A2(n_206),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_49),
.A2(n_50),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_49),
.A2(n_50),
.B1(n_96),
.B2(n_97),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_53),
.C(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_50),
.B(n_66),
.C(n_159),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_50),
.A2(n_97),
.B(n_274),
.C(n_277),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_57),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_57),
.A2(n_111),
.B1(n_240),
.B2(n_241),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_91),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_58),
.B(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_73),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_63),
.B(n_66),
.C(n_69),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_66),
.A2(n_72),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_66),
.B(n_97),
.C(n_127),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_66),
.A2(n_72),
.B1(n_172),
.B2(n_173),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_74),
.C(n_84),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_68),
.A2(n_69),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_68),
.A2(n_69),
.B1(n_143),
.B2(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_135),
.C(n_143),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_69),
.B(n_84),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_69),
.B(n_80),
.C(n_234),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_69),
.B(n_122),
.C(n_132),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_71),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_74),
.A2(n_75),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_82),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_82),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_120),
.B(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_82),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_82),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_82),
.B(n_121),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_84),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_136),
.C(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_88),
.B(n_99),
.C(n_110),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_89),
.A2(n_90),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_90),
.B(n_182),
.C(n_185),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_90),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_90),
.A2(n_230),
.B(n_231),
.Y(n_286)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_96),
.B(n_127),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_96),
.A2(n_120),
.B(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_111),
.B(n_239),
.C(n_240),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_112),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_134),
.C(n_147),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_113),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_130),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_119),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_121),
.A2(n_122),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_127),
.Y(n_129)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_126),
.A2(n_127),
.B1(n_210),
.B2(n_211),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_127),
.B(n_132),
.C(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_127),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_130),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_134),
.A2(n_147),
.B1(n_148),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_135),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_136),
.A2(n_140),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_140),
.Y(n_228)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_143),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_154),
.C(n_165),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_165),
.Y(n_153)
);

XNOR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_163),
.C(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_175),
.A2(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_196),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_176),
.B(n_196),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_195),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_195),
.C(n_215),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_189),
.B1(n_190),
.B2(n_194),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_193),
.C(n_194),
.Y(n_213)
);

OAI211xp5_ASAP7_75t_L g322 ( 
.A1(n_197),
.A2(n_323),
.B(n_326),
.C(n_327),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_214),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_198),
.B(n_214),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_213),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_212),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_200),
.B(n_212),
.C(n_213),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_208),
.B2(n_209),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_330)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_256),
.B(n_321),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_254),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_219),
.B(n_254),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_250),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_220),
.B(n_251),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_222),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_238),
.C(n_245),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.C(n_233),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_225),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_234),
.A2(n_235),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_246),
.B1(n_247),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

OR2x6_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI31xp67_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_315),
.A3(n_316),
.B(n_320),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_299),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_287),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_287),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_280),
.C(n_283),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_265),
.C(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_283),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_286),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_285),
.B(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_290),
.C(n_295),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_313),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_311),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_309),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_319),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_337),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_338),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_336),
.B2(n_337),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule