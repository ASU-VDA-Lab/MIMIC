module fake_jpeg_8507_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_27),
.B1(n_21),
.B2(n_31),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_47),
.B1(n_24),
.B2(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_27),
.B1(n_21),
.B2(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_50),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_30),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_21),
.B1(n_30),
.B2(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_62),
.B1(n_65),
.B2(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_28),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_43),
.B1(n_28),
.B2(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_89),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_79),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_24),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_0),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_84),
.B(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_44),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_17),
.B(n_41),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_33),
.C(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_40),
.B1(n_37),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_53),
.B1(n_48),
.B2(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_40),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_0),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_98),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_90),
.B1(n_32),
.B2(n_84),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_72),
.B(n_67),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_97),
.C(n_84),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_53),
.B1(n_48),
.B2(n_40),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_59),
.CI(n_54),
.CON(n_97),
.SN(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_44),
.B1(n_29),
.B2(n_18),
.Y(n_100)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_50),
.B1(n_57),
.B2(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_116),
.B1(n_79),
.B2(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_25),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_112),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_15),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_44),
.Y(n_110)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_114),
.B1(n_69),
.B2(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_57),
.B1(n_25),
.B2(n_20),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_130),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_133),
.B1(n_134),
.B2(n_112),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_84),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_106),
.C(n_109),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_77),
.B1(n_75),
.B2(n_70),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_75),
.B1(n_70),
.B2(n_80),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_105),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_101),
.B1(n_91),
.B2(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_136),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_108),
.B(n_32),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_74),
.B1(n_68),
.B2(n_90),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_91),
.A2(n_74),
.B1(n_90),
.B2(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_81),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_70),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_97),
.B(n_103),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_150),
.B(n_157),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_153),
.C(n_165),
.Y(n_177)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_149),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_97),
.B(n_111),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_124),
.B1(n_140),
.B2(n_137),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_158),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_97),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_138),
.B1(n_134),
.B2(n_119),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_104),
.B(n_107),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_1),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_1),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_104),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_120),
.B(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_133),
.A2(n_104),
.B(n_49),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_83),
.B(n_49),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_151),
.B1(n_129),
.B2(n_124),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_144),
.B1(n_170),
.B2(n_149),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_182),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_190),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_181),
.C(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_126),
.C(n_125),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_136),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_136),
.B1(n_88),
.B2(n_115),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_189),
.B1(n_154),
.B2(n_166),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_155),
.B1(n_171),
.B2(n_163),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_193),
.B(n_196),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_144),
.A2(n_88),
.B1(n_25),
.B2(n_20),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_168),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_162),
.B(n_25),
.Y(n_212)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_194),
.B1(n_175),
.B2(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_206),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_166),
.B1(n_161),
.B2(n_147),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_211),
.B(n_173),
.C(n_186),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_159),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_213),
.C(n_214),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_221),
.B1(n_184),
.B2(n_173),
.Y(n_230)
);

FAx1_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_172),
.CI(n_161),
.CON(n_211),
.SN(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_55),
.C(n_115),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_55),
.C(n_162),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_55),
.C(n_58),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_186),
.C(n_188),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_20),
.B1(n_19),
.B2(n_57),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_58),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_196),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_183),
.B(n_9),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_15),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_234),
.C(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_191),
.B1(n_9),
.B2(n_10),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_191),
.C(n_3),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_15),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_238),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_14),
.C(n_13),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_13),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_241),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_249),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_213),
.C(n_199),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_252),
.C(n_226),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_204),
.B1(n_200),
.B2(n_207),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_247),
.B1(n_253),
.B2(n_221),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_224),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_199),
.C(n_215),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_231),
.B1(n_222),
.B2(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_255),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_252),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_214),
.C(n_210),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_235),
.C(n_211),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_263),
.B(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_211),
.C(n_218),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_227),
.B(n_203),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_278),
.C(n_6),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_248),
.B1(n_243),
.B2(n_245),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_271),
.B1(n_273),
.B2(n_6),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_7),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_251),
.B1(n_237),
.B2(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_227),
.B1(n_254),
.B2(n_12),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_11),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_5),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_12),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_262),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_278),
.B(n_5),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_283),
.B(n_285),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_286),
.B(n_276),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_6),
.B(n_7),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_R g289 ( 
.A(n_279),
.B(n_270),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_7),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_292),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_274),
.B(n_268),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_294),
.B(n_291),
.Y(n_296)
);

AO21x1_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_7),
.B(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_8),
.B(n_287),
.C(n_295),
.D(n_280),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_8),
.Y(n_300)
);


endmodule