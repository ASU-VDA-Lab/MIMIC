module fake_jpeg_606_n_144 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_0),
.CON(n_33),
.SN(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_50),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_59),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_27),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_26),
.B1(n_23),
.B2(n_14),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_73),
.B1(n_75),
.B2(n_81),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_20),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_58),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_20),
.B1(n_25),
.B2(n_12),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_25),
.B1(n_12),
.B2(n_15),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_8),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_56),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_82),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_5),
.B1(n_7),
.B2(n_11),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_47),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_7),
.B1(n_53),
.B2(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_89),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_93),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_64),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_73),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_57),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_72),
.B(n_82),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_71),
.C(n_78),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_90),
.C(n_100),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_88),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_78),
.C(n_70),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_90),
.C(n_98),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_90),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_119),
.C(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_118),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

AO221x1_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_69),
.B1(n_74),
.B2(n_92),
.C(n_68),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_93),
.C(n_92),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_111),
.A3(n_110),
.B1(n_113),
.B2(n_108),
.C(n_109),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_128),
.C(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_117),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_69),
.C(n_96),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_108),
.C(n_74),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_134),
.B(n_128),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_77),
.C(n_114),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_127),
.B(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_137),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_114),
.B1(n_126),
.B2(n_124),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_126),
.C(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_85),
.A3(n_102),
.B1(n_69),
.B2(n_57),
.C1(n_54),
.C2(n_61),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_138),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_54),
.Y(n_144)
);


endmodule