module fake_jpeg_4490_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

CKINVDCx9p33_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_15),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_43),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_25),
.B(n_22),
.Y(n_35)
);

NAND2x1_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_19),
.B1(n_23),
.B2(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_14),
.B1(n_10),
.B2(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_18),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_26),
.B1(n_14),
.B2(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_28),
.B1(n_0),
.B2(n_4),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_22),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_52),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_24),
.B1(n_33),
.B2(n_17),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_28),
.B(n_42),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_52),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_46),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_49),
.B1(n_47),
.B2(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_57),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_53),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

AO221x1_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_28),
.B1(n_47),
.B2(n_6),
.C(n_7),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_47),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_63),
.C(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_64),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_67),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_67),
.C(n_6),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_76),
.Y(n_78)
);


endmodule